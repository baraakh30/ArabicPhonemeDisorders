`  �   ��?7�㾦8��f����x�s:Ҽ.->Q1?q�q�j���?0A�=P{$���c�-Ӕ��P�<0"Q?rK�?��I?�&Y?�6�3c2�z������y?1�>�F�>S۾`��>7�,?��O��Y��� �>G��?���?��l?P�F��Wѿ㶗������붾�>x�>�s>�s��닽=��'<�󊽁1T;�< >�>���>�΅>��J>�~2>� X>�5����"�k*���䔿T�:�����T��A�;�lr�@¾�x!��˰��;	���*�ؽTM�L�?�c��Hp��AW*�p��A?ᑤ>�2�>S��<�S�<�&��iû���u�o�p��Y���"�͹ ��sؾ[����-���z��e��y�v�?l��{�k�3?�5��r�<Ի?�*�=�=ʹ�>�\=�5>�Ď>�+�>���=�`,>��=c�{>�և=:��g���m:�׏Q�~9�;p�C?l]��~����3��d߾W���p�>�?ŦS>��'�������x� ��>2G�o�b���˽�� ��c�>ǽ�>��==JɻR����w�V�u�=担>�>J"m�#���)/�|��=�{�>�U���>��
>�� ?�0}?i ?)�i>�&�>���<Ӓ�>�[�>sk��so�< =>�J?5?�A0?�C�>d�j<�I[��D��=��=E�`��&>��=n���"f��޽�����S=>��=��={��}#Ƽ����x�����>Q�0?'��>z�?RШ���3�>y�����*>>w>��>Q�
?kE$?��?�?9>�Z����׾��%��=�>}�>�C>�4�l�3!����>+G>j�?H�=?����w���v>�cB>P!�>cL	?��?V�>_~>�����ɿ�v���d%��=���>8F�>'/��I%>Q.�>�u��F[���>���>:��>(v>�H">�O><s�<�T�>թ>�<��C���X��?=���~�_�iЁ�{���9k=��)>�!5>h<͖�=� 9;U���8��t�v�nt?VZ�>��ͽ�J��ob����F�ž�j?2D>=��>ʠ?\I�<��,��a�C�q����A?F�i?h��>��}���R���|>����+�>�4�> [p=䙔��#�;�+����� ׻>R��>�W�>!�:��0I�p���|]���8>��i=՟���?��O?v�־X���^'�)5�"���}˨��3{��룾�T���@�s�9���~���|����R>S��>���?8�}�r�<}�ƾE��8=q�Z���t�=v&>:��=ꪽ�>aK�I�!��"��������k� ?`��="��>^|%?��9?+�t?=Y?�0:?1{����N?�� ?/V�=��9?�DE?$L]?E�Y?�E}>cW/>���<�Y�� $��.��2<|��>��M>?m>�A�=�>��D> ��=����)^�Km�����3]�<#7>ť>ǋ?�A$?nC��������U. ���?=,�=v�S>�ļ�:e�Q�<L�s>�p?�M4?��>n�O=s޾� ������>�=oC?�*?4�>��<$��=��߾��]��E�=�L>Yhռ{~��5}�-S��r�ڽ	4�>T�>f��=��o>φ�?��?��>�����(*��&o�_�G��e7�H�Խ���K�d�fb>�2��d~Ѿ�⑿"���)m�6��=��E�Xr����B=R&�>�Ņ>mٖ���>��<�'6��t�=-�8>�٣��ہ>��?�#?�Ś>� �=���6�B�k?s�Ҿ�ca�љ������)��l�=���>��o��>�3�>yz,�Y���CN��=Ė�?��?x��?�X�=] Q�婓>D[�>��>�M>�J���q]�O%=��W>-��=�J���M��>>���X�la�>2mx���¾���~�I�/"���$6��6޽�˾���e;���?侌n��oRy��m4�_��jP��ł���(��w���{�d����6վ!�Ծ%��?���?��$>�`�<��E:�k���Po�7馾���b��o箾d޾�6�t�F��,���=��.���O�K`h>��#�U���{p�w�#�/P�����=�3?��sBپ���a��y��=�n��N�b���5'���>/�o}X?R|P?+�ܾ����6��W��l�>|�>�$�>G�a��հ���>�B4?��?�!�M?����t�<��=���?���?��??��P�"/A���ű��M?�:?t�>�}��W; ;�M?V(9??��>���6��L�a��>�~[?\�N��Yb>��>\s�>���@c����%��ؓ�$���8>�4�|��a�f���=�]/�=�"�>ǩv>Ox^�8ޮ���?4���s���AJ��^4����>�Q?A�7�6�<�H�>�eս���w%���,����!�K?� �?��F?@�k?Z�/�P�L�k� >Йi�l�"?�3�>Q�`>B���O�>�.
?=u\�e�D�-U^�SQ,?�0@#� @�y?ŮO���п�����H 뾺+>X��=�`>����>�Wz��J|:#�>X;w>	��>��z>F�O>Qa>�p<>�]>x�����Z���T��zYR�*�	��"�w�]��<�����[����%z�@����/�@�ýL�X���������r��������=$	?�$d>�l�>&Nֻ�U߻iD��f
�� �����V���A���L� �����=��搾��ϾK� �ijؾ ��>{��zt>��>�;�;>��>�E�{�>�!?=��~��!�=�yz=dX�=��=�R�>q�x>�u>l��=�����l����8��\�R�.�4Z@?�_������4�ݾ����nh�>M�?b�M>/(�Ɣ���z�N]�>��C�&`�{�̽Ç���> N�>�W�=֨�����t��M�˗�=/��>r�>�c���=���/��£=���>����d>X 7>7�?���?�K?�*>L(�>A�>>��>�8�<�
�=��>h�o>V.?�;?Pz/?7�>��v=�D�H�=�!>C���B���>����1�/>9��<
��@l=X,v=Ys�;���<1�=_����b�,�=ڪ�>�`8?���>�#�>�:�{M?��I��C��!>�2T��[�>���>�?bL�>��>�#>	W���ža��A�>��8>�[�gYr��8��x��>���>"�J?�q4? _ż��Y���<BD�=m�>�R?�%?��>ߌ.>����Q����˿1n*��s-��, =�ZӼ���=VDܽ��=���q
��"�>D�>.�?\��>�]>�ʊ>��=v�>���>R��=�ټ�O
>��;=!2$�.��=UZ�= �ཁ��=�)?�Hu����j�!�O�<�ȓ�9���J�N��<9�?Q�?�F��=���=m�[�hĲ���>?4�>�R�>�z�>�On=���_�T�8{E�I����>A�_?��?؇=�`%�=r��j$߼���> ��>��=��j�k��~-��8�;h��>W,?�Μ>?�#��1[�P�o�v!��ȭ>,S�=���	2�?[2?�����$�Y4�>TM��ؾ�l��}Ⱦaj���Ҿ��!�U]W�Ӄʾ:�̊����=(3�>���?1	���J �F��� 	����j�m���ڣ:��L����=�R�<Kw<ӧ-��(.�H�P5��/�� !?	�>Yp?�,?�D?��?��>ZJ?��:�Ou?X�>�)�>��)?�S?-PR?�?�z�=�4�=�;ӽ��?���w��.ڽ��=C$q�>�.>|pA>���=�fi=��<���=�_ʽGB˽S�=�R=��;;9S�=�Q�=�,�=k�=tt	?��#?�޵�Ƀ�=R������;=�?�=i>,���	~D�C�7=��a>�{?�[1?k��>mR�<�ݾ���n��a��=\�?��*?���>Q�V="�>���3+2�9�&>�aI>;�'r�Tվ� ��4k��>�U�>'	>�ug>���?��!?�3�>��(��+������3�*�n=��i\μ���>DF,>�վ��;�j~��D�[]h�T�>\`��q�#3�=���>D��=;P�D�>U��</��=I��E�>�7�>N�!>���>U�?�@�=�į�O�������r?����7�"pM���2����>tYo>p7+?&�LPB?E��>�|���g��[�z���?�:�?'��?DG�?�-�w�n�s@>�&?l��=]�>�%='H����y���>�=,(��Ƽ���p���[>�\<������澥��k�׽����"����̒��G:��������0ƾ�j�����5�OB���:��%ٽ���鐾�Ǿ�����?��?m�Q>ù�	/�	�=����~���G�������	��th2���v�?{ž�#侒G�dp>���0��6~>�(
��H{���z����rz����=� ?Jb��������p�����;�4��}S��ʔ��H���6����[?gKO?e�f(-����7��1?�w�>�3�>cž��y����>��>�B;?H�=ă{����|�=g��?�]�?X0??��D���?���R��x?<;?�v�>�;��}Ͼy7��V?��8?�f�>���0���Y�6}�>��^?�O���j>��>��>;ؽ�]����:�Ǒ�+�r��lE>�Y����	�3fd��A�k��=\��>�m>{�b��֩��?�Ŀ� ��B��=M�J���x�?d�:?�e����O�0?�?�>����y�c蠿��"�f?z�?\�m?=�K?�.�2�*�T�=�{(>V��>Y�b>;�=�����?�5�>����.B���Y3�ص6?���?�?:5v?ѡh�ĺͿ��������ҏ���30>
��>a�=>���!<>���=�7<��=�>�ܵ>Vݤ>��W>x�'>�k>���=kς��'�x����
��m��+���	�\"���˾(Oa����>��3l����}�d�Ͻ���;���#1��W��SE���N(>B	?:��>�>:�8>�{>��i���������'��*�"��c����;v;�)g�{���[D�
i��@�Ž����P�>��<�;�=�+�>J!��=�מ>�Q�=R�=�;>w�)>7�M>H�">�O>�x>	�8>���=¬{>&9�=�������o:���Q��5�;��C?D�]�Y�����3��p߾ʏ�� ��>�?A�S>J�'����y�%��>�:F�}�b��˽ӵ!��2�>n��>��=�2Ȼǌ�M�w��X��=�}�>��
>6_l� ���C�,��=lf�>|�ʾX`�=�mO>�?y�t?@�,?�0�=�j�>qnS>
��>�$f=ܬ>O�>�ŀ>}�?�`;?d�3?���>Ĕ�=�ob��f�<&�=ȃB�P9�
��ɞ��N���s=�K:�HV}=Ȏ5=�!��&�a=�N�<*K��q�;Uk�<���>P�9?ȝ�>�_�>�E$�q~=�ܹF��c�eC$>�,�:��>+P�>��
?�/?5V�>�I6>����)̾��@�>�]F>��\��x�;~�J�>��c>J?Z�3?��W�	�o��;=f�= �>��?V�(?Z=�>�">���G��'̿��?��a��
�>錚>g��;�n��ӭ�>F��>q�Y�zo>�ҝ>�R�>I��>�HU>�i�=�;O�,��>���>�I�=��Ƚo��==�A���<��T黈3üa��sW=�Vo��A����<B4�=����N򽘾j�$�����=0?���>ǧ�==���yҾ�r����륾&1?��`>��(>�n?E��U��r}����i���ؾ�>~l?4�M>�Ab����=�/">%>'��>tm)>+RP=T�}���>dә��Խ�Y�>���>b�>�Ƈ��Q�`:_��^!�L�Z>�)�;V���T�?'�F?fG�g��=v6�f�F������,��#��g,���}�<��ޟ>�b:�$6�e䯾r�-���>���?UC`�'1�=̑�,_���R���*�)-=���=6��>K�=���۾Y�9�����$j��W^>��?�/>��?�`??�V? ��?� ?�f,?�ȼ��K?<v��v x>��?��D?��X?X'?�ω>�+ʽ墲��%��v����/��tټn���ӭ=7m>G@>����=rb>���=V�@>��< )
>5�e>���=���=3�>���=,x?�#?�$����x���#�=&��_W<�P>�<O>��s�`�둗��=B>2�>��)?���>9�=R�Ͼ���`��]�=8�?��1?��>*��<�P�=E'�i�ys�=k�B>��Q����jh羛���;$��o�>�ی>���=rΗ>Ȋ?ڗi?̑�>�֞��1���E��$�$��][>j������`���P<u���iQ/��yw�hig��L'���<)�,|�=��=H�=Mv�>#�)>ͳ>m��}{����ܽ'Z;ې>2�>} ?._�>�H(>���,�žcB����q?�yD��N?�����G�/����d+>'y?^Cﾽ�7?)� >�܎��౿M�}����>�3�?=�?�ܙ?��9=\�v�oWf>�S�>���<銩<|�>�S`���>�،>�ڽ�����~�Z�xӺ�>B�$������=����߽�ا�I�C�}u�����G��@ൾV���C�C�p�+�2����$�����/T=d)�qC�����g�޾�`�ڑ�?)m�?u��>e�*=��,���.��*�7�<qmҾs���_z������k�π��־W6۾A�.��E��]J�5y�><5����x���\�e�<��E�� �;>�|?��ƾE������<�v7>���Hu,��.��!��Xѽ� r?QY?�jоt
A��W�.4��S?6G4?��? Y���\��	 ?!+?r	+?F�\��J��+�>�f>C��?�K�?q�??��O��}A�F!�"��&?
�?�.�>Ȋ�v5;t���
?-�9?�c�>T��S��g�*�>*v[?�aN���b>��>^4�>^�𽂃��v&�����ր��:>�����մg�?�=�9��=��>N�x>TX]��ٮ�b�>�<���`��4��P�6y���>�N??��T����>씨>��=A��6�� ͙�=o��8[?�l�?�"?ξS?R(�w
D�7��'�=���>�>X�/>S����>��9?d����z��"�?aR�?��?�.�?BpS������k����e�;
�$l�=m6�=�n>���8�=�Y�=�u��l䝼^�)>�:�>De>��@>��4>��%>�>�v���I�9O��&�r�2r�F3B�"�뾌�F�//)�<j���:������þQ����!���#��D�-i1����</Vþ�Z�=Q��>xbZ>�O�=�MA>�V/�Ѽ����m�JM�V�¾C$(��%� !�������"-��O�G�a7��>���Z�|��>����>@'�>���=:;��^��>�2�=H�">��s>6�8>k��>
_>0 �=��>24ý�q>��y>�)�=sń�s‿�E:���P����;ˉC?9\�;����3�(�߾�4��$�>��?�S>4'��|���Zx��^�>?�?��a�2˽��,�>�v�>�ָ=�4��P ���v�tB���=K`�>�>,����U�����!l�=���>'Pھj��=�ɛ>�P&?�9e?��.?��=�8�>��1>z�K>�>y^L>�;t>���>}?{+?O*?g��>2;>X.i�y(ػ�/�=6���.0�����e|ۼ�n<���<TΌ��U=���=vyL��=Fh;�L1��f<]�U=�
�>��7?޺�>e��>�t$�Z7�:�L�y����(>�$S��7�>��>hs	?Wd ?K��>t�%>����ž뾩��>�n<>LjY��9u�}D2�:Q�>�Uq>OsM?��0?-���iz���=5J�=�>�>��?Ҹ%?p�>	�'>�&D�����Ͽ+���} ��{��8�ɼaW��E3�i�'�� �;4v4�rj	�
���6L>�Cy>l��>�JU>�r>�.>-��>5�J>A�=0��=�mt<��(<d[@���J=���"�^��&�X�N�T���������z���Z�T��1}!��:����>j^�>
mm�������r۾^Eо
?ڳ�>��>��>�T_��$�!�V�eOF�t}��:z�>��^?�ҳ>q�G��X�=�	�=pG�=w��>V��>d�=O��B0���V�� ��=�&�>��?Z��>I�~��c��9y��*��Ȗ>��=z�����?��\?����w�-� �F�F���	�~�=U�?p^��߱��p!���9�[@��3���x�tR�=j�>6�?�z|����=)N�������샿�ǰ��#X=�Yu=6/�>��C>' +�Y"���W�c�վۘZ��;1�>5�U>�\>OB?��)?y��?�9/?���>���� ?���I�s>�X@?�\?�6d?��O?ⴋ�u`$�5t��aUR���>��eε��_�=iS,=D>�Ei>}b,=4/=t�������J=�T�	=Q�=���=qz�=S>��=�?��"?�)ܽ�>�s��
��!�<>AWP>�z`��-g�عq;�[>-�?k	0?��>�Zg=l�ھ�l�r! �ZY�=v�?��2?��>�9�;H�=�"�Q�����=|7U>��_�É���U��a!���>P�>=��=�u�����?S#;?���[uA=[��������T���#=w���{-�>���>!ш=�w��b޾�������KC}�i�7�g�����=��I>�oI>N�>�㔼#6a=��I�,D�4�H���M>	�>��>	�>��>:�C>~dɼ��*�ξ.�	y\?-�/�y��<�����d[	�P$�>ץ>VAھ�f?�������'B��Irv�:�U>u��?��?1w�?�a�=I����>�7�>�G�=��+>H�ν��]��=T��>�%4�y~Ҿ9��$<����=�s>�~��k���Ի��ߣ�N�����#���I�^b�g����b��a���[���&�Q�����I��� ���6b���>��U����W��z�2���+�A]M?'�d?�+�������G�����z��G��=��ݾ���9�����/=�>$�F
ݾ����%��/��.�=���%9z>�_�Y����_p�M�.�q$d�'zO>@�,?~�Ҿ1ࣾwy�Fc+=�j%>�<�"��$���P-��d��}W?�;4?�������O�+��Ѡ=͸?���>�T>�*��2WսmϘ>ؕ2?�#?ڷ��(J��.C����s<�Z�?zR�?A�??I�O���A���y���1?6�?���>�����̾z��#?��9?�ͼ>8� g���;���>ޛ[?`;N��Zb>���>�G�>'�ಓ��(&��7��0=����9>d�J���Jh��$>��ԧ=� �>v�x>�]�C����?�Ŀ� ��B��=M�J���x�?d�:?�e����O�0?�?�>����y�c蠿��"�f?z�?\�m?=�K?�.�2�*�T�=�{(>V��>Y�b>;�=�����?�5�>����.B���Y3�ص6?���?�?:5v?ѡh�ĺͿ��������ҏ���30>
��>a�=>���!<>���=�7<��=�>�ܵ>Vݤ>��W>x�'>�k>���=kς��'�x����
��m��+���	�\"���˾(Oa����>��3l����}�d�Ͻ���;���#1��W��SE���N(>B	?:��>�>:�8>�{>��i���������'��*�"��c����;v;�)g�{���[D�
i��@�Ž����P�>��<�;�=�+�>J!��=�מ>�Q�=R�=�;>w�)>7�M>H�">�O>�x>	�8>���=¬{>&9�=�������o:���Q��5�;��C?D�]�Y�����3��p߾ʏ�� ��>�?A�S>J�'����y�%��>�:F�}�b��˽ӵ!��2�>n��>��=�2Ȼǌ�M�w��X��=�}�>��
>6_l� ���C�,��=lf�>|�ʾX`�=�mO>�?y�t?@�,?�0�=�j�>qnS>
��>�$f=ܬ>O�>�ŀ>}�?�`;?d�3?���>Ĕ�=�ob��f�<&�=ȃB�P9�
��ɞ��N���s=�K:�HV}=Ȏ5=�!��&�a=�N�<*K��q�;Uk�<���>P�9?ȝ�>�_�>�E$�q~=�ܹF��c�eC$>�,�:��>+P�>��
?�/?5V�>�I6>����)̾��@�>�]F>��\��x�;~�J�>��c>J?Z�3?��W�	�o��;=f�= �>��?V�(?Z=�>�">���G��'̿��?��a��
�>錚>g��;�n��ӭ�>F��>q�Y�zo>�ҝ>�R�>I��>�HU>�i�=�;O�,��>���>�I�=��Ƚo��==�A���<��T黈3üa��sW=�Vo��A����<B4�=����N򽘾j�$�����=0?���>ǧ�==���yҾ�r����륾&1?��`>��(>�n?E��U��r}����i���ؾ�>~l?4�M>�Ab����=�/">%>'��>tm)>+RP=T�}���>dә��Խ�Y�>���>b�>�Ƈ��Q�`:_��^!�L�Z>�)�;V���T�?'�F?fG�g��=v6�f�F������,��#��g,���}�<��ޟ>�b:�$6�e䯾r�-���>���?UC`�'1�=̑�,_���R���*�)-=���=6��>K�=���۾Y�9�����$j��W^>��?�/>��?�`??�V? ��?� ?�f,?�ȼ��K?<v��v x>��?��D?��X?X'?�ω>�+ʽ墲��%��v����/��tټn���ӭ=7m>G@>����=rb>���=V�@>��< )
>5�e>���=���=3�>���=,x?�#?�$����x���#�=&��_W<�P>�<O>��s�`�둗��=B>2�>��)?���>9�=R�Ͼ���`��]�=8�?��1?��>*��<�P�=E'�i�ys�=k�B>��Q����jh羛���;$��o�>�ی>���=rΗ>Ȋ?ڗi?̑�>�֞��1���E��$�$��][>j������`���P<u���iQ/��yw�hig��L'���<)�,|�=��=H�=Mv�>#�)>ͳ>m��}{����ܽ'Z;ې>2�>} ?._�>�H(>���,�žcB����q?�yD��N?�����G�/����d+>'y?^Cﾽ�7?)� >�܎��౿M�}����>�3�?=�?�ܙ?��9=\�v�oWf>�S�>���<銩<|�>�S`���>�،>�ڽ�����~�Z�xӺ�>B�$������=����߽�ا�I�C�}u�����G��@ൾV���C�C�p�+�2����$�����/T=d)�qC�����g�޾�`�ڑ�?)m�?u��>e�*=��,���.��*�7�<qmҾs���_z������k�π��־W6۾A�.��E��]J�5y�><5����x���\�e�<��E�� �;>�|?��ƾE������<�v7>���Hu,��.��!��Xѽ� r?QY?�jоt
A��W�.4��S?6G4?��? Y���\��	 ?!+?r	+?F�\��J��+�>�f>C��?�K�?q�??��O��}A�F!�"��&?
�?�.�>Ȋ�v5;t���
?-�9?�c�>T��S��g�*�>*v[?�aN���b>��>^4�>^�𽂃��v&�����ր��:>�����մg�?�=�9��=��>N�x>TX]��ٮ���C> ߴ�K�&�Q`q�u5,�jh߾0ȼI�?B ��^_>��T=Fb��'�A��9��@��譼R�a?A1�?Y�Q?�_?|� �ՠh���,�l�>�m*?k�8?bum>�Nݾ�_B?6p�>FW¾jB_�$���BD'?U��?�?�lo?�^G�m�տ�A�����Pԥ��!>��K=�=��7��/�=l�{��G=�婼d�>���>1|y>>Y�&>�GZ>��{>�>���>(��w������B�?��%�� .�'�ǾT'�ĸI��(�`�޾����aÍ�R򰽜h*��*�K���e=�u��)��>�6�>���>KT�>e�>�OO>p>������a�����2�!��l׾�����6����x���������о�|���
�j�'?Զs<�߼��>E��_�h><�>�β=�=��>x��=e�V>��>8{|>���>���>�6d>sÞ>A>8��������.�wҽ��>��9?��ھ��E�W��U�z6���g?�b3?V8�>ģ��p����r�9�>Q�!����<�4"=a�9�g�=xe�>-A�=�̀>yVe��������=9}�>��i>c-�=x\���3)�ǅb�=C[=[�>�ľ� >��d>��?�Nq?��+?���9��>�L>��x>��>}8�=��.>�eb>\v?�J?T�6?c�?�=�=���t��A���9�,����V"��15�:��<���Kżŧ=�%�=_���1=��<�
=0�=Ȼ<�M�>)�-?�m�>�G�>�]�׷1��F�/@i��$>�a��G�>w��>���>(��>H
�>IsT>;�o<f���5��v��>�~o>�a��x�w%�;*�y>#�m>�0G?_M=?�.׽0b�!��=�^==�Y�>`�>v�'?e�>�~>򥒽���/�ܿf�/��C	����;����-��mC��%��[�X��T��	��[ǈ=xn>◐>Y�>{�\><�:>4�>ߓ?��>���G�>�g��;d�-����i�=YY��ׯ!�W��]d<����@�潡�m�y��cc��?R��=c���?��1?�(->P��ɳ��}��	�q%0>< ?�>�Y�>�5`>@��A_�R�R��p6�IA?�{p?��V?�g �C�,>�&�=��={�>0��=c�8���r>^����=��=Z>Ó5?�$>�GG��8\�� j�����S�R>�(\��%t�R��?�F7?M,�h뎾م,�=6r�o��v�
�r�A�����7��I��1����}d�x{��]�>_�>�d�?߼;��=��Ⱦ
 }��Q��xɾ��=v%�="��>���>kK	�!���t�E��c�,c=za�>sK?��O>���<�F�>��_?Ɗ?ӻ?�N?��>b�(?@��9�/?�A/?it?J��>:8�>�5�5.���z>��˾W�0�����G�ս!�";X6��H��=��>�3�<w��=q��i\�:�W��eu<\��=��=Ȝ�=-�(<3)>�u�<�?:� ?���"�H�Mt(�K����>�?>S^��<֨������B>�� ?�.Z?�0?*�=�^%�ʸ��*/�H��>�?�j)?,�-?���=�]�;R�޾�T�}E<�ǧ�>/�=�p��ai�a��.�������<H���y>ٲ�?�:]?�h�>���=���Bj��1f��*P�>=4>&&�>l�>S��=����XU�A�x�S_�������Cu��=s8=��=��>ٕ�=3�>�Z����@���H����=w@_<wn
?mE�>c�>��>L��<�پq���P?����.e��iE��^��f7�>S-�>�~�=p+)�;dx?�� �iX�������^��n$?���?Q��?zB?���a!<�͐>ۡ�=t�X>%�P��载]:5�*��W�^>nǻ;h�Ѿ�4�ǁ�=t�,?��$?�^0�$'���m4��^��ǿ1�O��=�����ܪ��.��f¾�����a������~��?=K�	��Ö+�T���@������� ������J�?B��?i�>�==U*�3Q����[_���5���ѽ(����RX������!��(��)>���7��!�CI��S��>�yY��Q��X�|�>�(�2)^�{�>>'/?-�ž�(���g��2V=�^$>���<lv�֊����b��3�U?�:?�W�!m���ӽ�>�8?���>!V >�r���)�ө�>9�4?l�+?���2��{֋��:��{/�?Ƒ�?��??�O�݀A�L��m��*?�x?��>����S�̾j���?�9?���>l�^�����>$�[?�nN��ob>���>?>�>�C�δ����%������z�9>������EKh��>�L��=�ՠ>�"x>r]�1M���t�=<<���"8�Z.���W۾G~���⵽�?�	��g�>e�1>c�r=&�9������P�K=��Z?���?�n?�q?�9�g�p�����-��=��?�5?�ƥ>p2�/a�>/�>�]����3�o4��m�?Z��?�b�?�Qc?_m*�-�οY╿�8��K���4�>�R�=���=^�*��	�=ͫP��>�=/7�=b�i>�̽>Y�z>�p>��>}�]>��+=�%��SV���������7E���-��[8�F��� o�5Ϥ���0�U���Ѿ�ݽZ��Z�!��;���;>�@�M�!ֈ�H/�=/\�>81k>Q޸>�ϔ>ѱ�=�Ӭ��׾�������?<�� ��� �����c������j���'߾����W�Ҿ���>��(���h=Ɯ�>𣓽D�>X�>4�=���>v�>�.�<�';>ݞ�=_s�=�4�=��h>E#;�>�.>�
E�$(��R�������4�S�w=)0?eu;��þ �>������U2�>:�?G�n>,�e獿҇���>u(G��ˬ�K�7�'Y��~<>6�>���=�@�;0�>~b����=�9<>�#�>S�S>��?=	�U��;��ף>R�>gk���=�c�=EC&?�p?K�2?)~C=F-�>F�X>	�>2O�=�Q`>E�>�;�>l�?�i,?�?���>���=l�|�1�>�`�=��-�?���{-׽3���-e���<j��M+=hLe=H������A�<KX�b=��=Bn�>��9?���>CX�>�3�j�;���I��h���>��3� �>��>�Z?���>Ο�>L�+>�!���ƾ��辬)�>%]>>bB]���s������(�>Dx>^�L?�M1?6J��Z���J<Ƀ�=&��>��?�)?X��>�(>s���[S�d�Կ;� �g�%� �D�����ɉ<F.B� eJ��y;�I����=U{p>�0�>#�u>�/B>&>�!>k��>*?>���=��=�<�:�����<m�"6=Et-��m;�Lj�i ���뼋���E����3i�ܢ3��5������S?��/?R�=ʛ��>��KE>��\��i��>���>�/!?��?�=��7�{b�QR9��y�=<`>V?�;?Uo��km�=�Ț��N���"A>�$!>�}>��r=����ܻ�"�>{?B�	?`t�=(�:�N�T�et��I��,J�>��T=�}N�}��?L�F?v���F6�����{<>����7כ���;��w���Tž�{���*��ɾ�#��5"�Z��=un�>�ɬ?��I���>[9�)̔��V���Ms�N[Q=m�W=��"?b|=��N���1V,������W�D�+=?�>�_�=���>U"?UKP?,a�?VGW?o�)?��=*�4?m�g>{?/�?[}w?�\?*?cx��)@;>���<�]�d��@T��xS���kU�Ό5>M�=>,�=���n>9r�=x/&�Mη=�X=]�<.��=xN�<�a]>���>�K�>�?N�	?�����s=0����Akg>-@��I�D>�-L��/��T&���n>M�?8�Q?�X ?�>��%�.�񾙧�{�4>k�?�>�>��:?�f->8nνacԾ���Ama���=?P[<�0����7����n�����Ayn>�"���>Cz?GoX?�,?�&L��9!��>�����m�>�}���?C�?���<1-��ژW�%�w�;�����,��T
��"�u��=��=�> >�>�na>�">��	��
���7�������X[=��>���>���>�a?>���<���ô'��9e?�c�;�t��c���`�z�=Yc�>��>3�+�+�?�󏾣'��Q��ܭ;�S�?3��?�<�?J�I?բ��
����b>�>5�><ѣ�S�W�5	+=�½�ϧ�>4���t�5ɾݾL>��>1��>#EK��Lؾ$gS�ڵY���ѿd�W��������EM[��辸G��{����m�A,��tn�
򸽥�'�`���\.�x"��������&EȾ�yv?�k�?�oh>�=0x�ě@�E���/�=�a���)�����J��"��T�(����Ҿ�� �0�쾡.ѽ))�>C*Y��%����|�\�(�(?���$>>r/?;ƾ�ô�
�� �g=��$>�0�<�pﾑ��������
��eW?��9?����"�����x>�?Ș�>v�&>�%���z뽘�>*
4?�h-?D����n���i��Ri�?��?�??�#P�*�A�~�����?��?b��>d����̾�{�?Q�9?٤�>��5Z��0����>L�[?k'N��Ub>E��>n�>G�M�����&�ja������0d9>���3#�Fh�@.>����=�Π>Yjx>�6]�<쮾���=�;G�:�Ґ�C� ��پc�^���>�O��0d=������7�G���<?�� *�=�w?��?��?�	f?:����qV�����!�>s�	?H�>��?�о)� ?ʜ�>6�5��/'���p�� �>�y�?�	�?��x?�D�i���%��I��BC����'>�W�=��=�X��\�=�N�<��L=+�r��M�>�)�>�`�>��T>2
�=�>�ZR>����a�!�n2��5��UI;�d��`_0�9���+��־	�������}������s������Z3�G�����<�����>�TX>��>cL�>���>�:>5�"y��C�
��$s��?��Ⱦ �#�	�o�%�;�r��_�_2ؾ�.����q)?S���|#�;,Y�>.�֢�:E��=������>4��>�"&=�k�>f�=��=.F�=P��=GmR>*?z>�~�={����)��eX8��L�\/�;��C?�[��n��mk4�\>ᾟި��Q�>��?��S>	�&�����y���>0�@�I`�*�ý�����>���>ޗ�=����x^��%q����ʼ=��>>����7���Jb��=E�>?5Ͼ�9�=ƒ>��/?��v?%�:?j�s=���>+5>徦>�>���>�1>���>O�?�m-?*.$?���>�.�=��s��	=>&J={r�~���������"�kY�;���;�A=�z%=��=�r8<¨=�=s�לI= 3�=� �>�%F?U��>�z�>�A=���%�'�.��L�A->�\a�D��>�� ?(�?vv?<?�>���=���h|��@ ��C�>9�>s�T�q�j���o����>y��>Hf<?�-'?�:��L��_:��9>l�>O��>(� ?��>>�3>`="��mӿ�$�@�!��fP�g߈;n�<���M�(�7�-�Y�����<�\>J�>��p>�E>��>�<3>�R�>�HG>�ф=�=�:�;Z�;�E� �M=�
�+DG<V�P�ꆯ��$Ƽҟ������I���>�k:��8ټ�d?:-?��9>�7���L��=o��0A�>!�>��*?�,?��P>	;��� �r�a��L����>L?�-?���f��>�~��6�f�K>��>\g,>S2��ʅ������>$ͷ>m2?��=���?_u�f	u��d���'�>�6>M����ɗ?J,a?���7�p�,���E�|�侷I?�*�i����� ����&7�ﲡ�" �����'`�>�B�>�?�����q=u�����^q������Q4>�	L>�N�>�滻5�꾷;t��E�z��w��=�'|>�9�>8�>��>���>��<?C�?�L? rf?gx���@?�r>7�?R��>�g?:� ?��.?d,ӽw[u='_�0
�=�����䠾�)�u�	>�>�>=K�>:�����޼@��=|�?=��9���l��6l�=�]�=�#>|>t��=" ?�)?��M�xPl�P.�G�.��7^=�bX>��R>�e�OӾ8D9�m:>RE�>��6?��>CZ=e ;u0)�,S
�73>@��>י)?�?Ģo>Õ��9U��s�ս�=��|>1������0��X�z1����;�o>�>�C�>ٳd?��K?XV?2����H�wB�m����>���=[�>�2	?�h�=֟��/*-�y�y�����k#H��������h���j�=B��=\��>�k!>�>V=w��>��K����
>5y�>{u�>1�?�,> M���X�RM*��:]?���|�����6��wO���&X>/��>O�+��?k���J�����������>���?w��?�Q{?��7�sZ���i�>�k�>(n�>��3����b>xǒ��L�>P�@�t�þ0��'��;���>�?�5S����.��j���,ӿVO�w��_�¾}�a�r�Ͼ8��+̺�ԛ���Љ��i�o����W������x�|!_�ks��X���Q��"�?�C�?OȞ>���<#=F���C�s���x=p�������Ⱦ�ا����z"�b�-��
��,��о�aѾg��>��Y�U5���|��(����p5?>-!/?�cƾBᴾ���
\g=�7%>�'�<|<�B���������WW?��9?^N����� ���`>L�?ub�>��%>�����{�>�34?��-?��t��o.��!E��n�?P��?b�??�O�ϋA�L�8���6?j�?W��>㢊���̾S��� ?G�9?z��>��)b���8���>��[?�)N��Db>���>:P�>�'𽣣��j&�=@�����3�9>k
����J?h�{'>��x�=	��>�xx>��\�����t�=<<���"8�Z.���W۾G~���⵽�?�	��g�>e�1>c�r=&�9������P�K=��Z?���?�n?�q?�9�g�p�����-��=��?�5?�ƥ>p2�/a�>/�>�]����3�o4��m�?Z��?�b�?�Qc?_m*�-�οY╿�8��K���4�>�R�=���=^�*��	�=ͫP��>�=/7�=b�i>�̽>Y�z>�p>��>}�]>��+=�%��SV���������7E���-��[8�F��� o�5Ϥ���0�U���Ѿ�ݽZ��Z�!��;���;>�@�M�!ֈ�H/�=/\�>81k>Q޸>�ϔ>ѱ�=�Ӭ��׾�������?<�� ��� �����c������j���'߾����W�Ҿ���>��(���h=Ɯ�>𣓽D�>X�>4�=���>v�>�.�<�';>ݞ�=_s�=�4�=��h>E#;�>�.>�
E�$(��R�������4�S�w=)0?eu;��þ �>������U2�>:�?G�n>,�e獿҇���>u(G��ˬ�K�7�'Y��~<>6�>���=�@�;0�>~b����=�9<>�#�>S�S>��?=	�U��;��ף>R�>gk���=�c�=EC&?�p?K�2?)~C=F-�>F�X>	�>2O�=�Q`>E�>�;�>l�?�i,?�?���>���=l�|�1�>�`�=��-�?���{-׽3���-e���<j��M+=hLe=H������A�<KX�b=��=Bn�>��9?���>CX�>�3�j�;���I��h���>��3� �>��>�Z?���>Ο�>L�+>�!���ƾ��辬)�>%]>>bB]���s������(�>Dx>^�L?�M1?6J��Z���J<Ƀ�=&��>��?�)?X��>�(>s���[S�d�Կ;� �g�%� �D�����ɉ<F.B� eJ��y;�I����=U{p>�0�>#�u>�/B>&>�!>k��>*?>���=��=�<�:�����<m�"6=Et-��m;�Lj�i ���뼋���E����3i�ܢ3��5������S?��/?R�=ʛ��>��KE>��\��i��>���>�/!?��?�=��7�{b�QR9��y�=<`>V?�;?Uo��km�=�Ț��N���"A>�$!>�}>��r=����ܻ�"�>{?B�	?`t�=(�:�N�T�et��I��,J�>��T=�}N�}��?L�F?v���F6�����{<>����7כ���;��w���Tž�{���*��ɾ�#��5"�Z��=un�>�ɬ?��I���>[9�)̔��V���Ms�N[Q=m�W=��"?b|=��N���1V,������W�D�+=?�>�_�=���>U"?UKP?,a�?VGW?o�)?��=*�4?m�g>{?/�?[}w?�\?*?cx��)@;>���<�]�d��@T��xS���kU�Ό5>M�=>,�=���n>9r�=x/&�Mη=�X=]�<.��=xN�<�a]>���>�K�>�?N�	?�����s=0����Akg>-@��I�D>�-L��/��T&���n>M�?8�Q?�X ?�>��%�.�񾙧�{�4>k�?�>�>��:?�f->8nνacԾ���Ama���=?P[<�0����7����n�����Ayn>�"���>Cz?GoX?�,?�&L��9!��>�����m�>�}���?C�?���<1-��ژW�%�w�;�����,��T
��"�u��=��=�> >�>�na>�">��	��
���7�������X[=��>���>���>�a?>���<���ô'��9e?�c�;�t��c���`�z�=Yc�>��>3�+�+�?�󏾣'��Q��ܭ;�S�?3��?�<�?J�I?բ��
����b>�>5�><ѣ�S�W�5	+=�½�ϧ�>4���t�5ɾݾL>��>1��>#EK��Lؾ$gS�ڵY���ѿd�W��������EM[��辸G��{����m�A,��tn�
򸽥�'�`���\.�x"��������&EȾ�yv?�k�?�oh>�=0x�ě@�E���/�=�a���)�����J��"��T�(����Ҿ�� �0�쾡.ѽ))�>C*Y��%����|�\�(�(?���$>>r/?;ƾ�ô�
�� �g=��$>�0�<�pﾑ��������
��eW?��9?����"�����x>�?Ș�>v�&>�%���z뽘�>*
4?�h-?D����n���i��Ri�?��?�??�#P�*�A�~�����?��?b��>d����̾�{�?Q�9?٤�>��5Z��0����>L�[?k'N��Ub>E��>n�>G�M�����&�ja������0d9>���3#�Fh�@.>����=�Π>Yjx>�6]�<쮾���=�;G�:�Ґ�C� ��پc�^���>�O��0d=������7�G���<?�� *�=�w?��?��?�	f?:����qV�����!�>s�	?H�>��?�о)� ?ʜ�>6�5��/'���p�� �>�y�?�	�?��x?�D�i���%��I��BC����'>�W�=��=�X��\�=�N�<��L=+�r��M�>�)�>�`�>��T>2
�=�>�ZR>����a�!�n2��5��UI;�d��`_0�9���+��־	�������}������s������Z3�G�����<�����>�TX>��>cL�>���>�:>5�"y��C�
��$s��?��Ⱦ �#�	�o�%�;�r��_�_2ؾ�.����q)?S���|#�;,Y�>.�֢�:E��=������>4��>�"&=�k�>f�=��=.F�=P��=GmR>*?z>�~�={����)��eX8��L�\/�;��C?�[��n��mk4�\>ᾟި��Q�>��?��S>	�&�����y���>0�@�I`�*�ý�����>���>ޗ�=����x^��%q����ʼ=��>>����7���Jb��=E�>?5Ͼ�9�=ƒ>��/?��v?%�:?j�s=���>+5>徦>�>���>�1>���>O�?�m-?*.$?���>�.�=��s��	=>&J={r�~���������"�kY�;���;�A=�z%=��=�r8<¨=�=s�לI= 3�=� �>�%F?U��>�z�>�A=���%�'�.��L�A->�\a�D��>�� ?(�?vv?<?�>���=���h|��@ ��C�>9�>s�T�q�j���o����>y��>Hf<?�-'?�:��L��_:��9>l�>O��>(� ?��>>�3>`="��mӿ�$�@�!��fP�g߈;n�<���M�(�7�-�Y�����<�\>J�>��p>�E>��>�<3>�R�>�HG>�ф=�=�:�;Z�;�E� �M=�
�+DG<V�P�ꆯ��$Ƽҟ������I���>�k:��8ټ�d?:-?��9>�7���L��=o��0A�>!�>��*?�,?��P>	;��� �r�a��L����>L?�-?���f��>�~��6�f�K>��>\g,>S2��ʅ������>$ͷ>m2?��=���?_u�f	u��d���'�>�6>M����ɗ?J,a?���7�p�,���E�|�侷I?�*�i����� ����&7�ﲡ�" �����'`�>�B�>�?�����q=u�����^q������Q4>�	L>�N�>�滻5�꾷;t��E�z��w��=�'|>�9�>8�>��>���>��<?C�?�L? rf?gx���@?�r>7�?R��>�g?:� ?��.?d,ӽw[u='_�0
�=�����䠾�)�u�	>�>�>=K�>:�����޼@��=|�?=��9���l��6l�=�]�=�#>|>t��=" ?�)?��M�xPl�P.�G�.��7^=�bX>��R>�e�OӾ8D9�m:>RE�>��6?��>CZ=e ;u0)�,S
�73>@��>י)?�?Ģo>Õ��9U��s�ս�=��|>1������0��X�z1����;�o>�>�C�>ٳd?��K?XV?2����H�wB�m����>���=[�>�2	?�h�=֟��/*-�y�y�����k#H��������h���j�=B��=\��>�k!>�>V=w��>��K����
>5y�>{u�>1�?�,> M���X�RM*��:]?���|�����6��wO���&X>/��>O�+��?k���J�����������>���?w��?�Q{?��7�sZ���i�>�k�>(n�>��3����b>xǒ��L�>P�@�t�þ0��'��;���>�?�5S����.��j���,ӿVO�w��_�¾}�a�r�Ͼ8��+̺�ԛ���Љ��i�o����W������x�|!_�ks��X���Q��"�?�C�?OȞ>���<#=F���C�s���x=p�������Ⱦ�ا����z"�b�-��
��,��о�aѾg��>��Y�U5���|��(����p5?>-!/?�cƾBᴾ���
\g=�7%>�'�<|<�B���������WW?��9?^N����� ���`>L�?ub�>��%>�����{�>�34?��-?��t��o.��!E��n�?P��?b�??�O�ϋA�L�8���6?j�?W��>㢊���̾S��� ?G�9?z��>��)b���8���>��[?�)N��Db>���>:P�>�'𽣣��j&�=@�����3�9>k
����J?h�{'>��x�=	��>�xx>��\����v��>�p��fM�gkG�3��`F(����<][?g��>D�i>��>��'�q��ɞ���V�NH?��?�QR?<M4?�R��Q�����:�=Hv�>��>!�=���.r�>o@�>Z��ւq�a�{�?e;�?;��?FCT?�o�%tο-����й�I��Ѽ�=q��=��B>���(��=/ׄ=�/�;:?Z��%>�W�>�P�>h*�>�v>ڊY>}�@>�����O$�b�������>�G���j�kz��&e��>�I¾�kǾ���нr�}�����xν�D������6�>���>~r�>�S�=�>�>� ����t	�2�Ѿ ~4�4c�o��e̾m���G��?��j�����7�}>y�=���=W��>�=�->���>��;~]�>6�n>� �=���>{0�>��V>��>�8>АE>�2�>�g0>|���r�����m¾��C���W?'�����ΆѾ`5,��J�%$��2��>0{>Q�B�B=���0��T��>�c�.]�\(*����=�t?��>N>����>�H��o!@����=���>��M>�K�=C��W���:h">ѓ�>���Y8	�v��>�?y6�?-�b?�F>���>��>~+>W吼�F�>\d	>��>l9+?N�?	%?� ?�׏=���2؅=��]>D����H�kp��KY�y�<�����ѭ�#�x=�D����$>��f<ʈ�>��ƽ�+��Q�=�0�>�kA?"L?E�>��,��i,�U�z��J�k��`m:�H�%?�
?c\ ?�{"?/��>W3>�=�����(�Zd�>h�<�|�qfs�o�>O�>2��>�`�?��>��=�5]�+��r;��l>n�A?A=?��?@�$>���P �9)��(�����A�h�ƽ��u#Ͼ/n��@M>��&�h}���kV�*#5>:�=�/X>�k�>�>!�`>\3�>�Ag>���=���=�=Է�:�W۽[� ���ܽD1�=?iH�Ntͼ��=�����;���b�S��оѽ�¼�?&?���م�B�z�k����=��"��> �>G��>q�>B�=�e��$Z�΂F���^�U�>g?���>!YQ�!)�=l����<�,�>:/�>�>(>�-��K��㘾6���@ѿ>]�?N؜>Y6���+O�12l�2�����>S�<D�нy�?"[?u� ����y�&���[����������� �v�����
`-�t.Ǿ]�������=�-?��?�$=	갾��w��e���¨���"�+�$�"D	��?.�?I�z�H�ξ��Y��V�}��FI��D)=
uO=��.>s��>��>�r?ϵ&?�?v�f>PA/?���>S��>��>i�5?�`?6�L?���>;v?��>vI�=��+4��Aֽ'+���U�=`�>�j�>�����~r=��{=�'>� 9��$��R�?ॼ�-��<���>$�%>s?�#?�{Ͻ�1:���ڼ�����<�~>�N>��G�ھd�&��9�*[>>o?��0?`��>Ѯ�=y�۾�i�F� �d�=�??=�0?�f�>��<�t�=M���u��T�=��O>ҏ^��+��J�[��w�t�>�T�>t��=��>Kz|?�
R?�%?������9����vxL�l�g�� ��XZy>��>�'>�=ȾO�M�%�E�K�T�?�-��6��h����/>��.>�wx=��(>Qrd>�C>�����}��OF�<1Q�=Z� ���>��?2Q*?�:�>�MR> �g�`�I?Η��2�<ܟ�Ѿ�7�Ʒ>ѻ;>R��n?~C���}�@奿�=���>{�?��?�d? "B��1���]>P�W>!
>W:<�6?��!��:��s2>�O�=�Wz��N��r̉;�z\>�=x>��ǽU�ʾ���W`K�\}��	L��n��&���3��(�¾ő��Z6��g����HἛM�^�оǩ>�e�=���&�XSi���������r�?�m}?�m>YE*�\�� ��R(Ծ=��i���B��e��+j� ʾ,���߾gA��	]���+�J����?�+���J��C����yȾT�C��p[=0k?J;��"X���2�!n>�|ս��X��m��0��Ѳ���.�Lx?'�?M̾�����6=��"=��>��>@�8>��= D=��>���>��S?Z�?>9���������=�*�?�y�?�sa?���A M������`���?>\T�>\2?p�j�����f#���}�>��?G�>�dK�����-�]�/?�?�r���A@>f� ?6�?ԓǾۣ�P�r:�������a>��-=�UӾ�+���þc
_�DB�>~�,>.�[����v��>�p��fM�gkG�3��`F(����<][?g��>D�i>��>��'�q��ɞ���V�NH?��?�QR?<M4?�R��Q�����:�=Hv�>��>!�=���.r�>o@�>Z��ւq�a�{�?e;�?;��?FCT?�o�%tο-����й�I��Ѽ�=q��=��B>���(��=/ׄ=�/�;:?Z��%>�W�>�P�>h*�>�v>ڊY>}�@>�����O$�b�������>�G���j�kz��&e��>�I¾�kǾ���нr�}�����xν�D������6�>���>~r�>�S�=�>�>� ����t	�2�Ѿ ~4�4c�o��e̾m���G��?��j�����7�}>y�=���=W��>�=�->���>��;~]�>6�n>� �=���>{0�>��V>��>�8>АE>�2�>�g0>|���r�����m¾��C���W?'�����ΆѾ`5,��J�%$��2��>0{>Q�B�B=���0��T��>�c�.]�\(*����=�t?��>N>����>�H��o!@����=���>��M>�K�=C��W���:h">ѓ�>���Y8	�v��>�?y6�?-�b?�F>���>��>~+>W吼�F�>\d	>��>l9+?N�?	%?� ?�׏=���2؅=��]>D����H�kp��KY�y�<�����ѭ�#�x=�D����$>��f<ʈ�>��ƽ�+��Q�=�0�>�kA?"L?E�>��,��i,�U�z��J�k��`m:�H�%?�
?c\ ?�{"?/��>W3>�=�����(�Zd�>h�<�|�qfs�o�>O�>2��>�`�?��>��=�5]�+��r;��l>n�A?A=?��?@�$>���P �9)��(�����A�h�ƽ��u#Ͼ/n��@M>��&�h}���kV�*#5>:�=�/X>�k�>�>!�`>\3�>�Ag>���=���=�=Է�:�W۽[� ���ܽD1�=?iH�Ntͼ��=�����;���b�S��оѽ�¼�?&?���م�B�z�k����=��"��> �>G��>q�>B�=�e��$Z�΂F���^�U�>g?���>!YQ�!)�=l����<�,�>:/�>�>(>�-��K��㘾6���@ѿ>]�?N؜>Y6���+O�12l�2�����>S�<D�нy�?"[?u� ����y�&���[����������� �v�����
`-�t.Ǿ]�������=�-?��?�$=	갾��w��e���¨���"�+�$�"D	��?.�?I�z�H�ξ��Y��V�}��FI��D)=
uO=��.>s��>��>�r?ϵ&?�?v�f>PA/?���>S��>��>i�5?�`?6�L?���>;v?��>vI�=��+4��Aֽ'+���U�=`�>�j�>�����~r=��{=�'>� 9��$��R�?ॼ�-��<���>$�%>s?�#?�{Ͻ�1:���ڼ�����<�~>�N>��G�ھd�&��9�*[>>o?��0?`��>Ѯ�=y�۾�i�F� �d�=�??=�0?�f�>��<�t�=M���u��T�=��O>ҏ^��+��J�[��w�t�>�T�>t��=��>Kz|?�
R?�%?������9����vxL�l�g�� ��XZy>��>�'>�=ȾO�M�%�E�K�T�?�-��6��h����/>��.>�wx=��(>Qrd>�C>�����}��OF�<1Q�=Z� ���>��?2Q*?�:�>�MR> �g�`�I?Η��2�<ܟ�Ѿ�7�Ʒ>ѻ;>R��n?~C���}�@奿�=���>{�?��?�d? "B��1���]>P�W>!
>W:<�6?��!��:��s2>�O�=�Wz��N��r̉;�z\>�=x>��ǽU�ʾ���W`K�\}��	L��n��&���3��(�¾ő��Z6��g����HἛM�^�оǩ>�e�=���&�XSi���������r�?�m}?�m>YE*�\�� ��R(Ծ=��i���B��e��+j� ʾ,���߾gA��	]���+�J����?�+���J��C����yȾT�C��p[=0k?J;��"X���2�!n>�|ս��X��m��0��Ѳ���.�Lx?'�?M̾�����6=��"=��>��>@�8>��= D=��>���>��S?Z�?>9���������=�*�?�y�?�sa?���A M������`���?>\T�>\2?p�j�����f#���}�>��?G�>�dK�����-�]�/?�?�r���A@>f� ?6�?ԓǾۣ�P�r:�������a>��-=�UӾ�+���þc
_�DB�>~�,>.�[����ϙ�>��羍�>��{.�����{�Ʉۼ^��>Ulھ�.>_\�>Kw�=��.��͎�CY���D=�_%?Me�?�X?2N5?g��45��J�w=�����ܣ>�2�>�q=�8_�mz�>{��>�jݾ�S��\��1?�o�?~��?�7C?��j��Rտ�a��G�ľ/�ž�_>u��=�vK>�Ȩ�)��=ԇG=<}�<�	���;�
�>r��>��>5>.#>v�*>`��>��Lٖ�e��UB��T����V���1��#��E���Lv�������[=y-����}??��yc�t����v!>z�(?t�?v��>�ި��C�=z�\����b���i��6�Q�+����ů�8d�I�ľ-*������Zu��q�%����?l��>�" >l��>hzr; >F>�ժ<��~>��>�Lo>��>���>$��>�F�=�9(>|2~�Z��>�9�<^~���k��3
��쨾-�.��n\?�Qf��վ�_
��,�$���Q�=�=�>V�=��:�e����6c��>(F��xI�+�'�ٴ�=��>M��>x>e>J7h>�+ܽ�x���>-�EX>��>��'>M׳�㿾_� �%�0>f�>���é�V>��?	�?[OC?63�<���>�ƌ>\d�>J�>��>�pj>uo?� :?��e?r݀?0��>�]�=н����<���=�\���+����=�Z=����Q�����g>J��<9w�
Yּ��q< ����V��9輖��>��Y?�G�>�ϼ>w�Ž�F�}Y���&�ܽK�¼y��>��%?vC?��'?�c�>4�;>����q��3�� �>�_�>|eP��z���ē�9�>	�Ƚ� ?S/Q?s�*�qT!��e#�t(=e!�>X�?O%?ID?,m>s�b>��	�#Jܿ&?3�~C�N���������<�n���y�;�Z�����w���2��ټ=�ǖ>�q�>�J>��=�(0>y��>�� >�g2=D0{=2.��Ǽ����a�>k^=�<�{̽­�=W�=-��_hK�K�wV3��H��9��z�> z%?(1��Ǎ��'�^����K��Ƣ�>��>W �>9�>
.�=D��V�L��{J������I�>�r`?�&?4�V�%|�=.�����u$�>o�>�_�=����1������|\0>��>8�>�_>�a���gJ�O	l��`�B8�>�=����T�?�j?;���Ⱦ=���Q���>�	5��P��d��:첾D�����8�ơ�~��u�⾩�Y��40?L �?Lbܾ�~��ؿ߾�ʀ������0��D>�������>�v�>|�v���Ͼ��$�� ��aV1��� #�G�5<��=||�>T9?180?2z2?M�]?�����7?X�>D4�>b\�>5?i��>y?6a�>ё�>�`>�<������g�;=«нO� >�@L>n��>'O��覯=�x<>?�;h��-y��*s>��#�t!�;��E>^�ڼ\�>�s
?/X5?`�<�=���q5�,L9����Ì=�ȵ>��V�B�=ͻ�>��?��?s�?�?�=���L�����]��t?�N>?^L*?zͶ;�%�>]��� ��?>�/>Yb=R3��#�z^=ŷ��c+�>�}�>�-�=�b]>=h?��??x�?u���TN�3eY��n�"q�]�>n�>�2�>�>���-���\���J�i.�(ʽ�J~�#�=J�>�&>8
A>Rª<1���6(=^!ܽ$���C�/=e>�<�[�>W�>�?Z��>��Z=�&վ�� ��H?�����q�.l���Zؾ�iw�A�C>4&>�9㽴H�>`t2��z�Ҵ���h4��	�>l�?���?eg?cLQ���ܽ�b>;>��>��e��2�@*�F\w�sS5>��=��n�弑�E{����m>��m>ᶰ�`9���Ѿ�S��􋽿[N��D��T�о��־��ƾ�U���:���s��2��2��n۾iz���Z��O��H�����C���� X����?o�?���>BL>}6���-"��"���c��(��x��_j	�]3��LG��m���4��R%���8�\�V?䝈����Kٔ�&���f=F�9�Q'%?9$��VE%���A��p�=�]ҽ'?Ⱦ�'�?9��OU��45D��-Z? �?�̾���#�����3 ?���><c�N=�<[f���1>G��>47?��?��ӕ�`񜿧r��Ԧ?c!�?�T?�j}�B��N��zQ�>��>��>�!!������iP�>)��>R�=��=��ާ���>��u�>��?~����|>�?��>�o����Yr��7���+ b�lf�>I�=eo�����>r��܂����>��>�ˁ���ϙ�>��羍�>��{.�����{�Ʉۼ^��>Ulھ�.>_\�>Kw�=��.��͎�CY���D=�_%?Me�?�X?2N5?g��45��J�w=�����ܣ>�2�>�q=�8_�mz�>{��>�jݾ�S��\��1?�o�?~��?�7C?��j��Rտ�a��G�ľ/�ž�_>u��=�vK>�Ȩ�)��=ԇG=<}�<�	���;�
�>r��>��>5>.#>v�*>`��>��Lٖ�e��UB��T����V���1��#��E���Lv�������[=y-����}??��yc�t����v!>z�(?t�?v��>�ި��C�=z�\����b���i��6�Q�+����ů�8d�I�ľ-*������Zu��q�%����?l��>�" >l��>hzr; >F>�ժ<��~>��>�Lo>��>���>$��>�F�=�9(>|2~�Z��>�9�<^~���k��3
��쨾-�.��n\?�Qf��վ�_
��,�$���Q�=�=�>V�=��:�e����6c��>(F��xI�+�'�ٴ�=��>M��>x>e>J7h>�+ܽ�x���>-�EX>��>��'>M׳�㿾_� �%�0>f�>���é�V>��?	�?[OC?63�<���>�ƌ>\d�>J�>��>�pj>uo?� :?��e?r݀?0��>�]�=н����<���=�\���+����=�Z=����Q�����g>J��<9w�
Yּ��q< ����V��9輖��>��Y?�G�>�ϼ>w�Ž�F�}Y���&�ܽK�¼y��>��%?vC?��'?�c�>4�;>����q��3�� �>�_�>|eP��z���ē�9�>	�Ƚ� ?S/Q?s�*�qT!��e#�t(=e!�>X�?O%?ID?,m>s�b>��	�#Jܿ&?3�~C�N���������<�n���y�;�Z�����w���2��ټ=�ǖ>�q�>�J>��=�(0>y��>�� >�g2=D0{=2.��Ǽ����a�>k^=�<�{̽­�=W�=-��_hK�K�wV3��H��9��z�> z%?(1��Ǎ��'�^����K��Ƣ�>��>W �>9�>
.�=D��V�L��{J������I�>�r`?�&?4�V�%|�=.�����u$�>o�>�_�=����1������|\0>��>8�>�_>�a���gJ�O	l��`�B8�>�=����T�?�j?;���Ⱦ=���Q���>�	5��P��d��:첾D�����8�ơ�~��u�⾩�Y��40?L �?Lbܾ�~��ؿ߾�ʀ������0��D>�������>�v�>|�v���Ͼ��$�� ��aV1��� #�G�5<��=||�>T9?180?2z2?M�]?�����7?X�>D4�>b\�>5?i��>y?6a�>ё�>�`>�<������g�;=«нO� >�@L>n��>'O��覯=�x<>?�;h��-y��*s>��#�t!�;��E>^�ڼ\�>�s
?/X5?`�<�=���q5�,L9����Ì=�ȵ>��V�B�=ͻ�>��?��?s�?�?�=���L�����]��t?�N>?^L*?zͶ;�%�>]��� ��?>�/>Yb=R3��#�z^=ŷ��c+�>�}�>�-�=�b]>=h?��??x�?u���TN�3eY��n�"q�]�>n�>�2�>�>���-���\���J�i.�(ʽ�J~�#�=J�>�&>8
A>Rª<1���6(=^!ܽ$���C�/=e>�<�[�>W�>�?Z��>��Z=�&վ�� ��H?�����q�.l���Zؾ�iw�A�C>4&>�9㽴H�>`t2��z�Ҵ���h4��	�>l�?���?eg?cLQ���ܽ�b>;>��>��e��2�@*�F\w�sS5>��=��n�弑�E{����m>��m>ᶰ�`9���Ѿ�S��􋽿[N��D��T�о��־��ƾ�U���:���s��2��2��n۾iz���Z��O��H�����C���� X����?o�?���>BL>}6���-"��"���c��(��x��_j	�]3��LG��m���4��R%���8�\�V?䝈����Kٔ�&���f=F�9�Q'%?9$��VE%���A��p�=�]ҽ'?Ⱦ�'�?9��OU��45D��-Z? �?�̾���#�����3 ?���><c�N=�<[f���1>G��>47?��?��ӕ�`񜿧r��Ԧ?c!�?�T?�j}�B��N��zQ�>��>��>�!!������iP�>)��>R�=��=��ާ���>��u�>��?~����|>�?��>�o����Yr��7���+ b�lf�>I�=eo�����>r��܂����>��>�ˁ���˭>��򾯏K�C,���������=Ě�>�1���n�>if�>v�>� �x��W�y�7M��2�1?ܐ�?�a?�K?h#<�����ذ>�\���lJ>q �>~�=bɒ�X�O>�O>%�ﾅTK�.l;E]?i�?�[�?FSj?{hO��Ͽ򟿄�Ҿ}@޾�b�<@{=���>?<�<�1�=�w6>~,��E��\�=���>#`>U�x>(Y�>D�>KfJ>>Z��G�����;ٖ�M9��4�Ei�W�!��-�.��O1���M������m�����:=�볽!������ɾ�u>�?��>#I>-ª>��W>�����龊7ݽ쳾=���h��\��r=.��|�@$C�kQ���uC���������m�>N1=��u>��?�8�=\$�>0�>� ����v>��>�i>��n>���>��,>��>�XE>׭>�v?>���y���Ō�¥��ö����Z�a?�z�3�
���|��I��PB�Ə���>��=<�\����C����>�k��u���V=j����<`"�>���>R��-=��Q;?����T<�_<�@5��={�=
�"rI���n>�>�ҷ���(=�,�>5�??�C�?uc?�>yR=?��>���>@��=�8�>`�V=(�>%�!?Q?�C`?#3?�n�<Lξx��;i��<��9��=�"�=��;����;�J����ڢ�;>'R�=o�%�K�Z�'�ν���<�}�>��j?�$�>׍/?��<��!�T�[������9�>�{���D�>��M?v1?�O�>�u?I?�?;a߾� �L4�>I��=;*V���^�j��&h�>�x>��?I�P?�yP�j5�zҽ,�#=�˿<O��>wP?.S4?�C�>6t8�� �|�ɿp%�`@�z4\�F���\*=��켟O��=q����
�%��={ߞ>C�Y>:v�>%k�>�>�Q�>���>7i�>zW�=��j>\��= fD�s�ν>����H̽��ܽ����	�7m�:�"�����K���)�$d���	����?�V?�3ļ�jּ��C�ܡξn���7��>��>X�>�`�>���=J�T`T�0�9���̽��
?Ar??8 ?}�?�p=if��u���h�>�ʳ>YGY>62|�r�&���j�D�=[�>�?{�>[3�K~c��f����W�>?>-�U�@��?�"e?�JH�nJ��H�;9O)��D	��H��6jL��C¾��⾐���f7E���߾����|�9Z0=z	?M��?!v��
c"��� �#ٝ��c���ᾨo>��;�C`�>Pt�=����'G�=��f���[+��%V}��U���ּ��>��>$?�>��>?e	8?�4?/U=���>פ�=�d>�?D>Bv?�� ?��?��>K��>xNx>R��=;���e��O&�=,��� ��=�8
>�>��=3C<v#>���=�����3�i�<�s�<�B&<E�U>�#>rC0>r?�N*?���`==Ȼļ���V5��	�=�J->��=�l��@��=Aڍ>���>�/?��>f5=����V�#^�[�g=q? G?��?� m=#x>�×����b(u=���>MI=8�E�~s��/��5�j��>�a�>k�}>�7�>/�v?�16?�@?�,����[�1�����v��V���SL>q�G<oˉ>���=vs��b{R�d_��vQ����	���`��2�>-B`>2�>M��>�L�>V>�<���=0��[# >����>�EA?�e=�d*?RM�>k]O>��|��X��}$H?��������(���/̾0Rʼ(�>�2>o`ٽ �?��ykw�f̡���=�	��>.M�?�z�?�>e?��5�U����Q>r_>��>3�ѻ�T2��:��<@����(>R@�=�:v�v�� �p���g>$l^>�ܽ�*��QgϾG������8J�+f�= o����P�*�Ⱦ@a���_�=́Ծb���F���}�� %V�pBo�L.e9�袾��"�
���I��
��?�kW?VՀ�IY���"�B� �I����=�2����d�a���8���ƾ
�����ܾ��1��9E�tg
���>:�]��䚿����M��8���`=��?�ܾ��Ǿ�Y��<���҄`�����琿���=e��|f\?{�?ŉ��$I��w���	8gt�>��>l|=�d/�k�㽝0>mz�>Js'?�t�=O����>���!����?���?Y�J?�i8��?�0�(����?��>T��>���>�����j¾\�n�Đ�>��>�MY>-��6n��� L��O�>��e?�r�K�q>W?F�>}���O[Ͼ_5=�龌��#�>��=~+L�5򮽡fM�.��'%u>���>�� �C���P�=�|��g[�����9�!�GG�a9�=�c�>h���=��=� ?Os�V^2��#h��b��9�Ƽ0�o?"��?��F?Q%r?�R�4J���V�PO�=ӱ�>��>IC|=��	��8�=r6?(���蚿_%���>�Y�?�A @�ng?	`}�eй�z���]�x�����>��>�u�>p�2�J�=�=A�B=�k_<Y>!��>��?>��m>�P)>T[=>-`�>s���g�����餿j�S�j�7���#��@�f��]M�h�Ҿd�	�SG �
�½���r72���ؽ�V<�o=μѾ�yO>X��>Z�? ?�e�=h{j�������˾0�h�Ac$�K��UB��5�E�H�,����$C�ߒ˾(������m���H�>��O=`�6����>�Y��MF�<��i>�=�<���=��=Py>Jy�����=�{j=5��=GM�=_�� v>���=bR����~�.�7��_N�WjK;��E?VU�5T��¶6��l�F������>G�?ֲY>@$�*���!2y�E��>{�B�~�U��ȽC�8����>(п>��=#(�O��Br�y�ｷ�=�,�>�J>i￼b���CW����=��>�tԾj��=�){>>(?r�u?*�4?�w�=ܚ�>8Kd>�>�l�=S/N>�/U>rl�>��?M�8?˻.?#��>���=F�[�2R=Hd1=�A��X����J���"���j<^�%��	E=,�j=�6,<��V=�(=��ټ��%; ~�<���>�d#?��>X��>�B�64:��I�N
�=��,�奆=���>���>��?�0�>/�>��=#�(N5����d$�>��=�j���z���pf>��M>��\?C=?%��=����r3=�	7>���>�G�>��?�R�>�9�>=������lӿc$���!��킽�N�Kш;�<�"�M�b8@�-�������<��\>Q�>�p>�E>��>�:3>YR�>,IG>Gф=t�=02�;��;��E�A�M=���<G<Y�P��G��g*Ƽա����0�I���>��<� =ټ�H?q?o��e�Vq������B�J!�>A�~>?H��>��7>J���YmK�[�5�)=��&"�>m}?ۊ?�5ҽgm�=y�ѽ����3�>ӣ>^\�=$�Q�E��K̞�8�]���>͇?�.�>����B��W�(Ҿ�K�>��jr�Vw?��O?��.���I�F�O�R�a�ξV���T��a�=�����d�J�>�	��H��f�׾�}���=�>u�?+sc�"b�C����}�N����A{�<"��>}#?���>}��=� .��5�g���GľN6n>��4?�N/�iF?)�!?͋?�t9?_�C?��?� b�^a?#�þ\��>�C�>��.?�V?π-?.>���;X-_��M�������:a��⪽��#�h��=�G>�)>�7�=�%�=�>A�=�:<�Z�=-J>�>�F->�ƃ=ʠ���⌽4�?�4?�ӳ��*<���;D
E�ZJe=na4>��7>	s��c��(�	�&�C>���>rk ?�V�>���=�5׾?�6�)�>��?�,?���>�]T=�B�={=��O�N�@�c=��J>gw���,��(�羗٭�:�����{>��>>���=8z�=��f?�E3?�8�>"Z���	5���Q���˾܂羧ő>l��>he?I�U>͵���YQ���~�mS���pҾ���>�X�L|=�u�>pr>E��>�>+�1>_U<l���w������S?�MG7>5s=b� ?2+q>2�'>�Va�!���/}?�v�fr��|t����z�=��?�����h�>2@�>b?>�;��)���d���?��?'�?��?i|��AP����>�>R>i��>k�>1?��4����=�j�=;�8>����KE�1�:>5uK>�p>�p���D��(�(�(Ţ�@����!@��
����Ԃ�Q�����þA�%�M��<�:n(��o��I��u��3�_,#��$U��:徃��Q��?�Ղ?,�R=�Q�^#����X��@C^��d|�r0���!�����<Mv�y�����ȧ�`+>��W�ml�᷐>�y8�����B�s�HG-��6=�=�>��!?G���)�������=I�(>�7�<��������ט���,�X?�@:?�۾����2���==�?���>�E>����NY��R�>�+?��0?�Oü?։�g���]L����?���?��c?M!�P���Ӿ>\?�ɖ>!Gj> v?��ǾwŅ�c�>���?��B?u��>����󅿥�$���<?+�Q?K<�O_�>ٛ	?κ�>M����ž7
�>VԾ9���I=��	���.��J��S2���D=��>�RG>����n]�ED�>�t��pM�����-!�"`ܾ�cR=��?�\!��s?�{ջ>�-:�w����_�V��>A�L?{e�?���>���?{~3�5�s�z侺nʽ�X�>|+?�B�>�"H=7�>5�?c��@��\�,��h�>��?>�?��d?L]�Y�ۿYؘ�����j���M>ƞ >\{->C������`�%S�;���_�=��>b�~>��T>0�?>ŗ$>>g���u{�ي���X���h>�lq�/N��R�:E�� V�H��Gȫ��˵����X�.��L���t9��h���|��Ǝ�!��>^�?G0?�ȧ>��Z>&>=4�������p���*��+!�D��� �¾+��񃤾��X��4�e�� $��ky��8�>�*�<�it=F�?
����	>�E�>����+��<g�>˗�=�a>G�>5iP>�&>�:>�N�=�>m�O��$��ڔe�֠���<�G�>a�w?�O�=����D�����_H��?��3?�D�>�����2���,L�*��>'�������c�<�q���Ξ<��>P��>��<�ω������ü�z�>r�z>W��>PK���v&�6��Y��=�>�Ǿ��~=��	>�.#?r�i?Ĭ8?��=�W�>.9�>s
R>�A�=�A>H�>�<>d� ?4VV?	�3?̬�>���=Ii��7�=�=4}J�PQ���f���F��~���<A���w3�=��=���<?_;y��<{�%�㡘�#t	=���>�
3?���>R��>�e޽oB��x@��4���=7{��*H�>I��>]_?N�>u�>��>I�}�ߪ��U��P@�>��=��p�vX��j	����>`6u>�3Y?6�"?���H�7��<���=��d>`�?F�D?`��>��6>J^������G���Z�l��>�����<��H�+�5�u%����=�iB�2�S@�=���=t|!>>�=��>�+�=���=��>�s2>���=��<H(09��ͼ�Ո�6w�=�\=<��>Z=���^�ޮ8���:��G��ϊ�g缌a�����P+?'��>hl>R����؃�<�*�* C��X�>6��=�5�>�4?#C>Ö���9�K�q�u����:? !h?gV�>z���N)>�C*>��>v>Y�&>���x��������&����`=��=��?���>`�n�9��Rz��ǩ���+>�aI<oN���i�?*�^?�)
��4���s,8�f��]1����I�!�����D��D^2�����.
��=��H�H=,6�>:��?D틾c�=0�ľl�����������jG>J�=���>�I>F_n�U�i�2���Ͼ�jI��l6<l$�>�P���)1?7?�� ?�kA?z&]?���>Ė�S�?�����>)�?9�b?=�?A5?�U������PD��I=9�E��A��@Ͻ�|��D�=0�8>-	�>'�k=!̱��V�="��=F�	>�z>,#u>cR>̥�=�t[=�=h�C>,Q�>S�>Z����S
=X���`N�iy�>X��>�ϣ>J�=�ύ�:���[��?�?�2�>ơ�9�.���ھ������>2u
?�8?���>94�=�._�wG#��I��n�:;N�=�N>�˧�����$�ܤ���v�<��?>i�b>�9f>�T?��5?t~�>{�=��(��rr��!�i]9>�{�=/ۆ>�K	?[9u>7�$��R3�I5����c��(��j ?����A�/=}��>m�Z=a0�>
*�<~I>�����%�����<f�x��6�=4�~>r��>�_6>��S=,Xw�\���1_?\:5�ک^���(�I�8����U��>���>%KżCv�>$�>�zG�C����- ��?�&�?���?P09?J��H��e$>}�	=L�=7�V>��4�/q��~�����>М>󦫾����*O=o?&[l>
Q��ڸ� dI�fz��ȿ8�2����;ܟ�)��e����:�z�!��뾿	��(�����ba<���׾�&�|���-s������V۾U�?��S?d�k=lO�=`���m �)p����A�C3���И��
��ߩ¾���������ľ��þ����a��#쾨��>KT��Y��W�f�xN3� �[�W��;B��>d� ��]����xj9>�P�=I��=j��<Ҏ�L���h[8�-hs?��+?� �Z�����+<>�<�>�->dOJ>�ݴ��^��΋>�2?�a??����U���:��.�C���?.�?z�;?Zr=�V2�B���� �m�>8��>�,�>�	N�z �����P�?xg??C��>�	�;ɇ�}�!�i�>>�x?�\�=�=>}�>Tݥ>�]��zF�������F��x{�k�)>�+�<tc8�,�;�~C����=�j�>9'm>�aF�T�߾d��>l$��aQ��kq�"���e���0���?�0Ͼ�<�RW>$t�=؂�q��>d�����=��(?�ε?�"?��\?������Q�H���Q=�>Y�>-��=�v`�z+?%J�>��׾ p���9��.�>���?���?�?T�^̶�{���D�d�҂�����=6
�=�/>�r ���+>�h=l���!�8=]	3>�	�>�~>�t>�'>bzF>l�=�?��������<͔�OlJ���0�Hr,�m/�v��?3m�(v��C̾tξ�җ���~�{ⷽ_�l��
��f5��i���g6V>���>l�>��>��>�x-=i�ɾ���͚��"�v7�fCھ�\��w����򘾕"���{��� �5k+��v����>�7)=�~)>��?"��>��wT���b�<����M��>���>��;>a"�>wʃ=��=->u��
;{>�V�=?���i���WY9���N�w�;��B?�,_����{ 4�t߾�)��Ֆ�>v�?��Q>��'�"����x�Ay�>�B��dc��tν���r��>��>�Ӽ=қ���
�c\u��v��-�=Gԅ>�#>�3Q��X�����.J�=��I?ݫ���0>%�0=�2�>v ?�?��>���>���=�c�>R��=�ۍ�|��>�Q>d�:?��=?��B?��G?��>
�]�"�>�W�=�b@���,����&��==�\��ʇ<wl&>��.>\E�<g���	��;m	+=�I��";����@�>ED?�>�>�I�>z-i��@?�I�H�D#@�ku>w9e��I�>}o�>�?fp�>�E�>�� ��{�fy��J[��"��>JS>��G�� ��AA��R0>6�X>��[?q�Q?<e�=��E��0%>��=���>��>�-?ۡ?+�"=�3>"��mӿ�$�;�!��xP� �;��<���M��n�7N�-�)���s��<�\>8�>��p>�E>��>r<3>�R�>�HG>�ф=��=A8�;p�;i�E��M=�jDG<'�P�^����$Ƽ������N�I���>�@:��8ټ��"?^מ>��l>UV<*����C�L��s,?�"?:�?N?M?��>�*���#?�q�G����)�>|G�>v	L?a��>��/=XX�=y{c>e�M>X`T=�ԡ���)��G����Y�=�I?H[j>dA���&��[���;�> 什[3�o��?��?�����ҾI:�� 0�s�%��>�����#[���˾�0��#�
�#��M������q?D�?��R�)�:����L���t����=�ڿ>?�=R�?��>wBi�;��)A��`��$p>��?�����^?W<9�3�>5-�?�E�?Nea?|�*��.(>S:�=��=QA<?#8R?�sU?���?
>�= .��k�ܾ�-��+����^�A:>KH���[$�?�<'��=d(���-7>�V�<�=xl=��=p��<B�t<���=I�=��n=	@�<�	?E?�Gj<k��=N��;��h�ï�=>0D> ��=���9ɽ�+�?"z>�j?ۮ?W�>�"�<S.��%�þ�i(�	��>��?�>?NM�> ,> ��=�F#�1܁�%��<������͠��x�3�:�p����>h\G>�?=P�E>�K?��W?�4?��3���+�����iᾷM1=1/��L�>Ճ�=���=]��T1��V���j�8��O�<]?���>M��=r�!>ݵ?W��>Ĥ�='�;��T����뾩3����zR�>��Z>�?�>D�l����?� �,?�[/��e���2��⾯����O�]��>Ue޼�u,?�J��ꆎ�����j#��ȉ>ɡ�? �?*;o?�窾 #M���>�b><G�>�}��d8�7l����̯�>7wX=k]��g7��[�p�%�>5z�>����}�ľ-OH�+����7��3&1���Ͻ��Q���o���V���T=�ڟ3�<z`�V
���k�ǰ�d\;��si�����4$��p��S���y+?��S?)<���;a��cJ���׬�=[ᾧ�R��
j�G	�<����F����=���d4�?����/ �#�Z>�LR�e�]��_�����-��=��?rؾ�],���.�\����>4h����#��������=J�#?�<N?���w�0�����`�N�>W��>L6k>¦}�ӡ���/B>�kC?i�#?��=;
��}��z�=���?��?R B?3`Q�/�>�������?�e
?���>�w��(�ɾ��ڽ$	?��8?�>z?�o���:���z�>{�[?ЄQ��Sj>���>�"�>���
O��_��۔�"ɇ��v@>���#"���\�M`7��=?�>�kr>�\�(-���<	?Q�E��zV�EF_�1�($���2>��)?6�A�6[q���?r1>�K)�@���q���F<H?K?[�?��2?A!5?�c��Vоa,�r�t<��>�v�>K�+>����4c�=�?� .��>�����>��?�{�?�� ?�(�y���;p����]s侙��=���=|�B>v#���g>�h�=^������Fl?>�}�>�>(�><�:>��=��k<�~�p��Ą��⮤��=��� �)f��#2�>Ӭ�=�I�0�&��{������GKh��k$��T��#�N�� �����Նd����> ��>G�?MU?���>�@�=�¾��i��:��x�	�����aLᾹu���ھ��W��u�n����6�ޓV�6�>�#<㊉>�?2�L>�>��>]$�>�6e<cv�>HF�>��>Cs�>� q>���>{�Q> ��==�c=��|(��M�L�-�}�B��\"�;j1?>잽�<q��\C�:p
����ؔQ>q-?akb>����ӑ�f���]�>�t�Uh�������<<3�>�Ʒ>tZ=*�)�r�G����Y)����;��>�l >�`l����p�
�ҥ�=`�>�A��^��<���>�?fJg?k�a?:�<AF�=Zv>��>&�>���>�o�>7	�>|?�D0?<?��a>"y(>'v��]�q>R�g>ПQ��W�N���f�����e�>\��0i���l�=vv]>��=�@=��ƽ��=��<(!�>O:?4��>~��>�x��+��P3�,ʙ<��>��5�
��>2b�>�>y��>��>�BI>�+>��3�:v�l#?�9���Jq���[�� ̾V/~�ڝ?\��?��S?��># %>R�>��i>ļ*>�R�>*M?.�?*"?=��_��]��Oӕ��sN��o���>��>�2&<��K�jú>m=�~{��V���=�f�AG>�}>��=��R��"��cѶ>��>$L�=��J>��>�Y�=���u�˼jh��������B=d�8>v�>��l=p�u�\3f���=�-�<��(;ʿ7?��W>^�Q={�=�W���)�����#?F��>�a�>c�?P!h>7-ʾ�
�l�1�1{2=3�>L�!?ի�>�X��s4X>�p��`	�8G�>S?��+=K���zn���߾�He�cx=#��>[kr>�r>�\?k��Rq������>2#Z=�z =*�^?��?3�ǵ����^�S����EO�>W����f������������L��u���O)>1�?U�?��n��r�<\p��j���9���������>�[��b�?&�w>���о�����󾍾���2�J:D?�'`�*� ?�c7?�?��?$�s?�O*?쌚�o?9�=�9p>$>�>�@L?X1@?mn?{�2>��">�ik�uj�=Q���|@���W���Pؽ^�>S�L>'󶼝h�=d��=�z
>.:%=�-�=m���ì��e'>al�=~�>"#=�5?�?��s�@�gԽ�3�ƅ�=�k>��c>,��@��|K�=��>*%�>s�?��>F��=ߝҾ�@ؾ�������=��?�]-?��>1��=�$!<Ѩ��9�Z�¸�=�K�=�9���x�2�Ͼ񵖾N��`?>�7Z>;;�=b�>J�S?��x?��>`_�����N��}2�H��= -�>I��>�{>�Bi>��h��b���e��n����V�P��>�e�^�(=�>8>�#��2�>.��=ҧ;?*%�� ���R���7��u��-�=�+�>���>���=��=�;�?��q�`?A�>�D<�7����\��^�>��?�G��R�V>|�>��N���(��)�J>���?s#�?��?r�c>=aY����>�F�=RW�>��=�>�@)���J�ݮ=�@>_៾���q��NZ`>�>�沾��@~��Q@������(�Ѷ���|��=���`���۾/�v��f��P#�k������
��t�)���H���S�^�I�%[���5��0w?P�g?7s[>��G>����%�����C����x5�sƾ�ݾF��N���v۾��ٚ�w�
�=�����>�mI�th��"W����`Gk�z�=�� ?6��e ��ɽ���=��	�;�����Β�J�=��N?ܓl?�%'��������f���>�?l��>g侨.��G?ž>?�/?��=�q����v��N��9�?�a�?�,@?��P��?��,���A]?��?�G�>od��E�;�m콾�
?��8?1j�>'��H{������>TY?34R��	f>��>�
�>����@��\'��i��]c����0>x������l�c��>��z�=�]�>3�q>��_�u���4u�>"XѾ�E:�iQ3��-���;�AC=c6?�XE���`��>�7����%1���L��.h�M/M?��?͗�>�c?}O9�+��t�w�����>�>F?�U>t1E�WOu>��E?ے���膿�B#���?�*�?��?~�e?_�R�0ֿ�Q��X��h���'$�AU>�>`�$��U�=� �;Q��<h� >�b�>��>�v�>�sc>i{�=g�=��s=-���� ����������m�����!�{Y�I��p�7�u�پ��b��B��ｻQ�����<@�����31�:;���>�?xu�>�]?���>Z��=dS5�z;���˾�_�[�"��	��;ξkD��WXI��>��o�ā�f�]�o����K?K�����,>�1?]�*<�}�T�>���=A�߼�qp>��=w�<��>�Փ>�L�=�>��ѻԧ~>#%�=ө���!���J:�H<T��D�;��D?��[�KЛ�k�2���پ�ɨ�%�>?r?jpX>g�&�F0���_x��c�>4�E��^c�T�Ƚ�F����>`�>.��=<y��G��,Jy����^q�=���>[>�$����b��=b�>fX˾�3�=��>& )?8u�?�9;?�o�<�:�>�n�>��>��=��V>�E�>�Ě>��?�p1?�?j��>�H�=�o�o��<�XG=��Z�b�̽,�4�ۤ��O�X�*=���<U��=���<Ef0����=��"=������ȼ+�K��\�>N�*?0�?��m>܌>Ư=��N}�2R����=K\����>�a�>�.�>pW�>6n>8W >U�G���B�V���?�$�<ƈ�O����E��^�=t��>D�?�@?��"�6�1�l�>~��>@`1>5}�>��C?��&?��=;i(=���4ʵ���}��$����5�il��x.�;ɋ�HgY=	.�>P|����=|/�>_Q�>-�/>lI��-O=�`�pE����>p+>v��<�7�>{԰=�kx��m���}�=�(����<�C*�������˽L��Q���c��ǉ�<���<5��= 7?ٶ�>��;/¾&� �?3��,���J?�I�>a �=|$�>%�"?���� V�f�:�N�=��>6?|[�>��r����>��OΜ=,��>@�>3>��~�]���ݽv��c>���>�� ?'煽z"`�s;4���ȾW)�>Ļ�=y�<��?'��?2f˾,ߐ���a%8�T���������qz�PT����4��j ��G
�f���hž�fR�*��>��?��@�b>������������N��Ѯ>\ ���>[�>o �;|[8�t(���(�;�ž�y<U�C?{����>�¹>��0?�'0?
J�?S?o��eH?�>V��ɺ>�4?��8?6�'?��0>V��:�:����>��<��C�Y��:�<#��=r �=j1�=��h�h	����=WR�=���oX�=�R>6��=�7�=ϕ�=Z���:�=��?Z?��ϼP�8�˚\>�7�Y>5mN>�ڟ= >��`���uZ>.�?+�>-'g>�W>\�m��W�����d>� ?��V?~��>ZJ=�.>%�3��z���ex��ź=ˊN�t�|�O��1����Vr�|�->�L7>��=`��>�Ki?9>u?��?&����qH�Q���7<�NZ�>$8���?��a>>���{媾�@Z��>��Mo��e,��?d�&��"���>�~�:T��>�����D�=P�8>r�i�v�L��+>�o,����>;yZ>⼝>�IY>'
����=�w�L�s?_�c��.�~�C�t�vz�����>��> �����>y��>#kt�)�̿<4���[?3�?,��?���?[ľ2�y�$"�>H�>|�z>�7�=t�ý�諾����l�>��==��ܾ���酽�t[>b�0���#�����9���*�3�����@��1�����6B~���r�Ⱦ������Iz+��`� �<��0���?��7��慨=CȾ#Zh���?�=�?�|�>EwF>�پ?���"=��c>Iiܾn����������T�������$i�?)(�5���0�ﾜ��>8~9��_���gl�j ��f��eC�=11,?j�ݾ𾾷�'��ջ@9>=1&���_$���&���սܒO?�I?�G�E:����@��=�b�>��>|s>�U�� V˽�>�9!?b�%?����c���J��#�T=&�?_T�?m4D?��"��r7���)O�����>�1?�>u���"��3�l�T�?�7?���>G"����O��%�>vpN?ll�TS�>���>�>���y j�����2��� ڇ��j>�(�;6��J�G�����[R�=/Q>�!{>]+�A¼��P�>X3���N�<�H�@���\�֗�<��?w��2�>b�i>�>��(�D������u��L?�o�?�/S?ܥ8?�D��)��1��Q�=O�>�F�>z~�=�]�MM�>�/�>���qr� ��U�?"$�?~��?�Y?�m�A�Ϳ�Q��%լ��e��=��=��=��@>_�潛�=�"�<���T�B;J�>Mϯ>'�>[��>��J>R�I>H�L>��T�'��ޡ��ڑ��E?�/���r�pg~��h	��������\о'Bоz�罦]�K��4.M������:��,�>v��>�[<d>�c�=��>��=J�վ�2־ж�k�'�J���~	��^�i��C��3վ�.��E���z�� �9y?��+��H�=%�?�`��R(=W+?��E>4F�>���>�b�>��6>hw�>���>$�r>
�>੽�3>UӬ�p��z��di>�yS��$^����[?L���=�޼Y�+�=�E��n�|>><�>/f������L���M�>_�t�Dۼ�i�����=]d4>x�?�2>zt���"!=n���W����^�<��>���<�30>,�㾏þݞ=>�/?�����ޅ��|><�? O{?�p$?�> �?ZHO>�n[>FC�>��>C��:3?�Q<?��'?c�V?fZ�>9�n=k�����껕bH���7=���Ƚ׽ɿU�g��'uӼ�|�=(��=V=.�I=p�=�J��摽l��k�>��T?�� ?�?)���W����j:��v>f	�>��&?|��>`��>�b,?��>c��>)QM>�Z�^� �ɭ�>W�r>q�1�X&w�o��=�%�=��=]�f?$�Y?�g=L=���.�����9<��>�?}I�>\��>36#����w`ӿ<$���!��y�����I&�;�<��NM��|�8#�-��<��s��<_�\>�&�>�cp>c�D>�u>cF3>�K�>ڎF>i��=: �=m"�;{;N�G��9L=����1J<�'P��f��%�ż����W���ZJ���=��z�Y�׼[�?Q�?f�8<�v������&�c#�>��?T�?��>��)=������W��m+�� ׽[L?��q?t��>B�/�TbO<��f��W�v�>q��>�>6腽J�j	���;c�>z?xI>�V�h�N��Ac���~Y�>�pۼ!n����?��S?a]5�����%���`��� �9+�C����z��G�˾ 52���Y������6�f���yf>
��>�C�?�fP���>�b� ����N��Z�7��@7��>�}�>��M>ɯ����SPV�z�Ѿ��R�>9�@G3=�q4>r'�>*%?E{+?	dl?)V"?W�>=����>�)= �>��? #"?`b�><�>��>���>!�<>�b��L�'/�!�7<tD���>8�=7e>5O�=��.>r(>��=�U)��P���yn=�=ٲ=�8�=ԱB>"��=��
?�p$?�ʽ5"�~���$�ڕ�<�{�=�tS>me7�ޙ[�>ø;��\>>v?��,?p~�>FT�=��־;��.����ǲ=�?D�/?�.�>��<���=�羉�y�{^�=�>T>�p|��C������}��� �>SD�>76�=�?>�̑?��J?�)?|���+!���~�0@��b�e���
���>���>�X�9���X�{�b�O�b�,�?�7��[�$�'��@����<o:v>1܍>�_�=
��>[�+>[���|�P�V+(>S!�>.�?EX+?�'?�<�>��>�=i�:�	�ÒI?�ɟ����
Y���:Ͼ�r!�%Z>�M>>O����G?���
�}�ƾ���=���>.`�?���?��d?|C�NV�0[>i�U><>`<٢:�o�uЃ��4>��=��z�������;��X>�2x>'ʽ�1ʾ	X�b�;��ȿr�{��>4��0 �.�ܾL#J�æ�����Љ_��e��i�����$D���dc�cm����������7�j���?&�=?��=��6>��E��
ȾZ�۾JM�=����B.��@w�@2ѽ
�ҾB򖾀�Ҽ`�^����?��ȾZI�>'�+� >���-��r�C�߲����{>��??��5�FP��/�����i�y�)>������%���~p�X
?��>�lI�qZ۽���;i�b�⨫>n�?~>D�7��$��-��>:&?�Z&?�ž��j��c��hĽR[�?»�?M@?T*N��D�3��S�&�W��>�8?��>MI���Jξ�x���?��1?8��>�%�I1����ܑ�>˾a?$�_��g>���>��>+�G/��uC��
D��ߘ�\!>�%�W�&�5U��y:�J-�=n�>x��>nP�+Ű��P�>X3���N�<�H�@���\�֗�<��?w��2�>b�i>�>��(�D������u��L?�o�?�/S?ܥ8?�D��)��1��Q�=O�>�F�>z~�=�]�MM�>�/�>���qr� ��U�?"$�?~��?�Y?�m�A�Ϳ�Q��%լ��e��=��=��=��@>_�潛�=�"�<���T�B;J�>Mϯ>'�>[��>��J>R�I>H�L>��T�'��ޡ��ڑ��E?�/���r�pg~��h	��������\о'Bоz�罦]�K��4.M������:��,�>v��>�[<d>�c�=��>��=J�վ�2־ж�k�'�J���~	��^�i��C��3վ�.��E���z�� �9y?��+��H�=%�?�`��R(=W+?��E>4F�>���>�b�>��6>hw�>���>$�r>
�>੽�3>UӬ�p��z��di>�yS��$^����[?L���=�޼Y�+�=�E��n�|>><�>/f������L���M�>_�t�Dۼ�i�����=]d4>x�?�2>zt���"!=n���W����^�<��>���<�30>,�㾏þݞ=>�/?�����ޅ��|><�? O{?�p$?�> �?ZHO>�n[>FC�>��>C��:3?�Q<?��'?c�V?fZ�>9�n=k�����껕bH���7=���Ƚ׽ɿU�g��'uӼ�|�=(��=V=.�I=p�=�J��摽l��k�>��T?�� ?�?)���W����j:��v>f	�>��&?|��>`��>�b,?��>c��>)QM>�Z�^� �ɭ�>W�r>q�1�X&w�o��=�%�=��=]�f?$�Y?�g=L=���.�����9<��>�?}I�>\��>36#����w`ӿ<$���!��y�����I&�;�<��NM��|�8#�-��<��s��<_�\>�&�>�cp>c�D>�u>cF3>�K�>ڎF>i��=: �=m"�;{;N�G��9L=����1J<�'P��f��%�ż����W���ZJ���=��z�Y�׼[�?Q�?f�8<�v������&�c#�>��?T�?��>��)=������W��m+�� ׽[L?��q?t��>B�/�TbO<��f��W�v�>q��>�>6腽J�j	���;c�>z?xI>�V�h�N��Ac���~Y�>�pۼ!n����?��S?a]5�����%���`��� �9+�C����z��G�˾ 52���Y������6�f���yf>
��>�C�?�fP���>�b� ����N��Z�7��@7��>�}�>��M>ɯ����SPV�z�Ѿ��R�>9�@G3=�q4>r'�>*%?E{+?	dl?)V"?W�>=����>�)= �>��? #"?`b�><�>��>���>!�<>�b��L�'/�!�7<tD���>8�=7e>5O�=��.>r(>��=�U)��P���yn=�=ٲ=�8�=ԱB>"��=��
?�p$?�ʽ5"�~���$�ڕ�<�{�=�tS>me7�ޙ[�>ø;��\>>v?��,?p~�>FT�=��־;��.����ǲ=�?D�/?�.�>��<���=�羉�y�{^�=�>T>�p|��C������}��� �>SD�>76�=�?>�̑?��J?�)?|���+!���~�0@��b�e���
���>���>�X�9���X�{�b�O�b�,�?�7��[�$�'��@����<o:v>1܍>�_�=
��>[�+>[���|�P�V+(>S!�>.�?EX+?�'?�<�>��>�=i�:�	�ÒI?�ɟ����
Y���:Ͼ�r!�%Z>�M>>O����G?���
�}�ƾ���=���>.`�?���?��d?|C�NV�0[>i�U><>`<٢:�o�uЃ��4>��=��z�������;��X>�2x>'ʽ�1ʾ	X�b�;��ȿr�{��>4��0 �.�ܾL#J�æ�����Љ_��e��i�����$D���dc�cm����������7�j���?&�=?��=��6>��E��
ȾZ�۾JM�=����B.��@w�@2ѽ
�ҾB򖾀�Ҽ`�^����?��ȾZI�>'�+� >���-��r�C�߲����{>��??��5�FP��/�����i�y�)>������%���~p�X
?��>�lI�qZ۽���;i�b�⨫>n�?~>D�7��$��-��>:&?�Z&?�ž��j��c��hĽR[�?»�?M@?T*N��D�3��S�&�W��>�8?��>MI���Jξ�x���?��1?8��>�%�I1����ܑ�>˾a?$�_��g>���>��>+�G/��uC��
D��ߘ�\!>�%�W�&�5U��y:�J-�=n�>x��>nP�+Ű���>�dؾ?.P��G�Zv��u<��4�=R�?g���=�)>�>�#$�┿4�������8?�T�?�EK?n\(?�� ����� ��~>��>~ɨ>j>���BA|>��>�!��BR����L�?Q �?���?y�f?��q���տfc��<^��5GоH'>+2�==+Z>޿g�pĮ=c!.=;[��b�q'�=:@d>�E�>�t�>�E>�>��!>"چ�n*����;Ӕ��:��;�t�u?_�P��~�����)���㾛m���ꪽRv��+���������r
�������_=���>�_>�Ӥ>�~c>��e>p��:��ʾ��a�vژ��ͷ��X��IC���ྎ)f�3j�0}4�i�����h���Z?n��=�z|;+�>l�e�R�b>ws>���>H`�=��@>���>l:>�L>:�>�|a>C��<k�T>L��=(Q����!�T�z�]��A��x?�=�HM�u��=��.�
>���=݊��˿�ʉ��Td��4�>���<'����F�X#<�O�=l�>�DB缏o��������^�>µ>�x|���=g���n;�� p>{�,?
y�)����"վ%�>O��?��?�#>#�"?���<�yٽ���>J�?��U>�v�>��O?��i?�pF?<�?��>_����r���]_=��-��>=�̽��J=��üH�������$C<lw���)ּ�쪻N/���v;�`=�4�>II=?qH�>���>ĕR�9I�
�6�@|���=}Da���>U"�>�L�>�L�>���>s>�=���ӾR�ľ���>��>ɴQ�{y��M�=��>2�>'yT?�jF?k��`۔�Ј>C�/>]�>��?��0?cR�>�.j>3콂��h�ҿ�Y"�D|!�V���(s�3M;�v;��X=�г:��"�ui��<)�\>J��>�3l>X�I>J!>{.>*��>AA>.�=��=�Ua;�S��c@���=#��4G<!���x�n��@��7���&TP��=��^��Oʼ��?B�5?�ځ=3h���K޽��z.žJ`�>"?�]H?��6?��W>R���SoE���"��{��R��>F%t?��&?�D��->s~�<	5�h�/>�Ι>���=�����Kj=��*��]��˼�>���>�X>_�R� r<���j������>�����r��/�?�n?��W�ľ�-8�P�#�R�#���=YWx=��������D��i}2� g�*2������e��?��>��?C�w���;>�!��e��?m>�����Y��Z��=��a>+U=�J���P��#6#�`Y ��Rr���4����>l�=F?%�+?c��>�c?���>W ?�sg���?�˅>�=�>C�>s�?�8?U�?h՜>V�S>��>8H+�;\��ɚ���ѻL�ֽF�Y=�+L>-�!>Ts
=�c�=6x�=N��=�^��2&�=������<�37>�~�>(��>��R>�4?�)?��k�<⑼3[=��3��c#=dg>�vT>ㆽ�W��'=Ϋd>�K?�4?m�>�r;0�̾)�㾶���@�=h??g*?��>��0=���=�1׾��/�H>�P>4⎽����T�꾋���Z�� �>�܏> �=>�7>@ԅ?��3?uM?K*=���^��X^� MA��𡾿�x�x˚>��=o�>���*��;-�!�m��fx�j�/�F���ݿ2�J�g=ie=5���_�~>��U<j�\>��8>�()��s��,�=�Q|n>�
�>�J�>
.;?�:q>K��kZ�:־|�I?蛡�km�G����nоL
�S�>��<>+���?�����}�-��WF=�Ȍ�>���?C��?B>d?P�C��(���\>IV>��>��/<�>����|����3>D�=�}y�y����;� ]>xGy>=�ɽz�ʾ�2侗�H�?�˿�`���	>)��"D�dg���~��|^�Z�����G� �s�ɾ�׹�Ur��(-��v���õ��dྗ�����?jl�?��q>�c�>��k*�`p���=�]+���H=d<?��a�%����ѣM�,,X�DtI�?�H�N|�c�z>���3���b_���(��!���K�>Q�-?��۾�塾�!�x8k��{=k=�����9��饘�_��TG?%�?=������~�9ݣ>*�:?��>\�>H0���p��ht>&I`?��J?���Cb�J��w=7ÿ?5�?)0=?�wP�,%C���	����*?�_?���>`N��\�;:���*?��8?=��>����e������y�>�PY?e�O���X>���>�җ>[��g���Kq�1k������bB>T04�&
��/Y��.�R��=@��>�T>@-V�η��'x�>d�澈QM��I�k��l�6[�<
r?@��z>[�m>l�>-�%�^ދ�m������\>J?���?϶S?��7?�Y��� �%W��8ֈ=	*�>�(�>���=���C�>�.�>j����p�� ��U?ۆ�?���?Y�Y?@�n�:Ϳ.q��J޹��vؾ�>crs=��x>�,���=�/��i�����ي�=t��>�֛>��>�>�<>H(I>4����1&�?!��l����R�	�6��A��pQ�����^���� ���fE׾�λ�y�����w�N��JK�<�;�C-��Ξ>���>S��>�S�>T�)>?8u>\���ga�� ������q%�C@Ӿ��Z5��U×��A�������+�k)*�l]n��?�웽��J>j?��-q�=��?�9&=��|>B��>���>G#�>���>1+c>d�=W(>���=��{>^\�=�*��Y���f:�JQ���;X�C?n]��0����3��+߾�x��l?�>�?K�S>r|'�ַ����x�K��>$sG�r�b��H˽�w�
i�>���>��=�Uٻi��x��JｬZ�=ێ�>�=>f�g�h������f-�=��>gǾ=n�=��F>�*?�{?ҿ9?��h�>t*/>���>=!�>�n�>s<5>���>AA?��;?+�<?�u�>H��=�TK��^/�j�x<����H�������p����7�g�U��=<���<CpC=�tI=���=H�)<Z�����<2d�>L�:?i �>�MB>�k����u6"�⺑��W�>��_>P?�-?�8?ί?G7�>��=��V�w|�������>Gρ=8�q�H���ܻ<���>�h+>�9�>��?��=세:�mr>̓4=��?�OI?RUi?��?���=�����|�ʿ�f���R�+Y7�?��y=�ѻ��U=�<��/^�m�b�*�V=RWx�;�>l�>1Zq>Fq3=$n�=��>�1=3]�<c��=��=oT>v�Z<��=�*h�*����(P�Yg=��=����z���Tt��(�?=��=8خ�̈́?;�?����v���܅��1��D��G�>���>V�>��>�I�=j4�u�\�R�K��xd����>-b?Md?�gS��R>K����=<. �>H�>|�8>�y�<h�}���k<� �>L?� �>�m��JP��ii�m��8�>����懾+��?�u�?+�&���\q����R���>�y�=/�˾�4���E��m2�9!����A����g�h�0?#q�?����>	!��2���5x���^�k�=���>�N?��=r��_'��:^2��)��ׇ�oM�`�>K��>��>K}U?hc�>��n?×C?�A�>�x��N�,? t���m�=�y�>�B?!h�>�?S	�>��>GY">u4����ɽ���j�=8h<���<��= ��=�P=B� ��ȼl�J˽C���0�<� x�(� =K8�<��=�>ړ?-(8?���/w3>��4>=V�=�L9> �&>B�ý@�`�k�S<3n/> *?�X!?{T�>$�m>����,�a
��
�^>II?��?�E?ν0�
��<9��HV���raH��˾|���?�l���`+�7�k>I�q>�<��l>�y?��;?U�>���F]>�J�6����vH���->��>K!>��߾)3D���g��\�U4�k��==���W}=�ɍ=�m�=[��>�r4>=��=V'k<&�;>Q�^ZV>�fI>��>��?�73?ʏ�>���=�����=	���I?����/������Ͼi��-b>��<>w�8@?Y���'~�i����<�^�>5O�?��?vc?��D��-�A�_>��W>�>oK)<(�>��~�+���ȿ3>�>�=��y�/@��}7�;4[>=|x>UE̽k#ʾǼ��F�'��ER��o������o���yپ���y�~�e㯾u�x��$׾���#��#�3��̃��=:��Me��Џ�ܢ���{�?��?�J^>=Z:>:D-�C�I�
���l�=�	�� ������h�h�Ƈ˾+�߾C�ܾƵ8��l<��6��'����>�R��Nc��!�F�3�Y�ɛ�8u����f?N0*��B>�B���.�����e��*ꚿ�)���pK��~z?��5?�>���ܾ����53>r(?]=?&;�>Y{�,�=�Z>�U$?�A]?�w>�l��R��]c��<�?�q�?Z�R?��z��7���.�����~�=E�>���>@-�󻋼���310>j�>��J>�C\�i��~~Y�i�/?cu�?������>� ?��>�%f�:���;
>��M<Kp����边�J����=�l��}z��E�>'�~>6�徇�����>�dؾ?.P��G�Zv��u<��4�=R�?g���=�)>�>�#$�┿4�������8?�T�?�EK?n\(?�� ����� ��~>��>~ɨ>j>���BA|>��>�!��BR����L�?Q �?���?y�f?��q���տfc��<^��5GоH'>+2�==+Z>޿g�pĮ=c!.=;[��b�q'�=:@d>�E�>�t�>�E>�>��!>"چ�n*����;Ӕ��:��;�t�u?_�P��~�����)���㾛m���ꪽRv��+���������r
�������_=���>�_>�Ӥ>�~c>��e>p��:��ʾ��a�vژ��ͷ��X��IC���ྎ)f�3j�0}4�i�����h���Z?n��=�z|;+�>l�e�R�b>ws>���>H`�=��@>���>l:>�L>:�>�|a>C��<k�T>L��=(Q����!�T�z�]��A��x?�=�HM�u��=��.�
>���=݊��˿�ʉ��Td��4�>���<'����F�X#<�O�=l�>�DB缏o��������^�>µ>�x|���=g���n;�� p>{�,?
y�)����"վ%�>O��?��?�#>#�"?���<�yٽ���>J�?��U>�v�>��O?��i?�pF?<�?��>_����r���]_=��-��>=�̽��J=��üH�������$C<lw���)ּ�쪻N/���v;�`=�4�>II=?qH�>���>ĕR�9I�
�6�@|���=}Da���>U"�>�L�>�L�>���>s>�=���ӾR�ľ���>��>ɴQ�{y��M�=��>2�>'yT?�jF?k��`۔�Ј>C�/>]�>��?��0?cR�>�.j>3콂��h�ҿ�Y"�D|!�V���(s�3M;�v;��X=�г:��"�ui��<)�\>J��>�3l>X�I>J!>{.>*��>AA>.�=��=�Ua;�S��c@���=#��4G<!���x�n��@��7���&TP��=��^��Oʼ��?B�5?�ځ=3h���K޽��z.žJ`�>"?�]H?��6?��W>R���SoE���"��{��R��>F%t?��&?�D��->s~�<	5�h�/>�Ι>���=�����Kj=��*��]��˼�>���>�X>_�R� r<���j������>�����r��/�?�n?��W�ľ�-8�P�#�R�#���=YWx=��������D��i}2� g�*2������e��?��>��?C�w���;>�!��e��?m>�����Y��Z��=��a>+U=�J���P��#6#�`Y ��Rr���4����>l�=F?%�+?c��>�c?���>W ?�sg���?�˅>�=�>C�>s�?�8?U�?h՜>V�S>��>8H+�;\��ɚ���ѻL�ֽF�Y=�+L>-�!>Ts
=�c�=6x�=N��=�^��2&�=������<�37>�~�>(��>��R>�4?�)?��k�<⑼3[=��3��c#=dg>�vT>ㆽ�W��'=Ϋd>�K?�4?m�>�r;0�̾)�㾶���@�=h??g*?��>��0=���=�1׾��/�H>�P>4⎽����T�꾋���Z�� �>�܏> �=>�7>@ԅ?��3?uM?K*=���^��X^� MA��𡾿�x�x˚>��=o�>���*��;-�!�m��fx�j�/�F���ݿ2�J�g=ie=5���_�~>��U<j�\>��8>�()��s��,�=�Q|n>�
�>�J�>
.;?�:q>K��kZ�:־|�I?蛡�km�G����nоL
�S�>��<>+���?�����}�-��WF=�Ȍ�>���?C��?B>d?P�C��(���\>IV>��>��/<�>����|����3>D�=�}y�y����;� ]>xGy>=�ɽz�ʾ�2侗�H�?�˿�`���	>)��"D�dg���~��|^�Z�����G� �s�ɾ�׹�Ur��(-��v���õ��dྗ�����?jl�?��q>�c�>��k*�`p���=�]+���H=d<?��a�%����ѣM�,,X�DtI�?�H�N|�c�z>���3���b_���(��!���K�>Q�-?��۾�塾�!�x8k��{=k=�����9��饘�_��TG?%�?=������~�9ݣ>*�:?��>\�>H0���p��ht>&I`?��J?���Cb�J��w=7ÿ?5�?)0=?�wP�,%C���	����*?�_?���>`N��\�;:���*?��8?=��>����e������y�>�PY?e�O���X>���>�җ>[��g���Kq�1k������bB>T04�&
��/Y��.�R��=@��>�T>@-V�η��U�<>�� ��1C�M+:�I��R�C���<C��>]���k��a>�%��B.9��g���Z��l���y?�ͮ?��0?�~<?ݵ�����W�.���=���>�
�>>� >x�8��7�>Kb�>����)fh����Mm�>���?�T�?��,?�h3�vԿ@��� ����ma����=M'r=��/>7�f�=����G�;*��=�>>p��>l�F>�l>� o>�@>�`>���]+ �\h��3ف�=fE�������q���B��#��Q϶��J�ٌ��GE���<�GI�����!c�XT_����>A:?d}0?�`>�hD>���}0�k�����؃4�At!�j7	��b���6�-O��E���
-�BH7�G�#�jB?��=L�	=С�>�N��5�a=�L�>o�n�BG">�q>�Ș>h s>��=�p>-��=w �=�{>۩>u��=�n{��'��=1��0��+�=�Q?_���7���6��<ӾS�X�-��>��?��@>8`-�f�����|����>�	�駊���;v=��x>���>�^=�I=�Qv<p2��Е���<��>f6>>#z�<�_g����Ʊ�6P�>`վ`P�=��s>=�(?v�v?��6?H��=OG�>{t_>1T�>�p�=�uL>�qN>u�>�:?�v9?�2?gN�>첾=��a��Y
=�XD=��;���L�M������68��<w�&�?J=F�t=/�;�b[=�I=���w�;Z	�<V?u/G?���>��>?׌�����?���</5g>To(���>��?��2?�?��>�z��׉��/�[���3��>�;>:td�ˈ���齍�>��s>�wg?��??��}�V񫾶�N��>ˤ?�?g?>��>�<�=�v��.l�i�ſ�T�dƾ띘���7�������`H�<
�B�~&}� ��;��Bʮ>���>jY�>5]�>��>Ε�=̘�>5C�>B��=X!4�����h����];���^���ܴ�����X�wǊ�3 W��כ�J���!�b�]=��O�?�k??Nn�=r"���8��� ������=�0?�Q?�C?&<�=�Ҿ|.���u���
����>/�?�i?)�����=�ۊ��oԼu�=	!">w�=�JJ>I#=��<��>�09?xW5?�q>
a��f��>�����I�?y�=B�(3�?Άp?:� �$q�V����k��9
� ���?�=�hۙ�K ���:#�@*�縷��P�����Wz�����>"�?�����ۂ�����T"���~t�AQ��z�C>��
=�l�>J�>{�D��1���0�����85h>~W	?v6�>�H>~?��?�ې>~�?�(>?12	?�w��@�
?�₽)��>̪?�H?Y�D?�w�>t*�=j=�:
�l�X��3t�d�����L>b�R>x5=�N����@>��r<����!��?�<��>����:�n��<��m�9j�=���=:��=�F?�/?ְ4�Q6�|���\챼Q`�>��=�j>���=28оԽdq0>�;?Up.?��>$������F	�����K>�z�>�k?�?�3�;+��<~���̾m��b�> ��¾���fW/�d6��}@X>|�e>M�j=���>IG{?b�9?t�[?t�1�&Ke���O�J���]+>� �>�x�>+�3?��> �����V�ٌ��:��4m4�Q=�>L�7�Wה��a8>��>	J�>�SF>0Ȍ>( 	�_A��*J��w���������>p�>�
?�A�>��g<���}� �=�:?>}վ��i��S���ؾ�8>���>��>�־�C?[�>xۂ�iY���I,��zC?��?sj�?��"?�/���=���=�+>��n>%���3`�l<>�"=T5�>�g�>�ꢾ������s<Ƨ�>���>�ˡ<���]�
��ؽv����tQ��L���˾�I����о�r���o΁�Z`�r�:�a��~����̴׽�<�ꝅ��u��Q���i��?3��?�N�=h'_���'�#��uTܾG��=鈜��Y�������C�����6�ܾnB��32���&0 ����#C�>Z�\��+��6|�!�*�j����^>V8?��̾�������D�S=��>p!��⾜���o���ѽ�W?t�;?�d�!����(�>�?0��>l[%>�������}l�>�7?j,?�W7��ύ�����W�U�?r�?�B?]� �j<�6��v꽫�?I�?˺�>�i��hϾ���&�?*�??�n�>�J��L���>s����>~�K?�T��vV>�T�>,ԓ>���"���er��3�����F%E>f�5;�\�[�r��<�@��=K��>׏�>ˉ>�����Q�>�ۛ���a�kOn���)���:�6O<�� ?^����<f��>�>�G�#�������Sj<:"J?�ë?�F|?�f?�
��fQ��W��F�n>�T?�?G�G>�h�'�=�i!?�b�ǘ��/R쾒2/?���?u� @��n?^2n��ؿS@���	���F��l�Q�/D�=ƴ�>v� ��Ѣ��6���<���<�])>BR�>��>s�=>�[>,x�=H��=4����,"��Ԣ�e薿�>/�Q%������K�ٯ��gP�I �P���➾A���Ҭz��a���\p�(��3㔽^�X���=>{�u>]��>3X?rBs>;z>��z�(�ܾ<^羊���H��x-�Y͹�EZ����R�� ��������@�.6#�D�E?����˼��>��R��̨�>��#>+�f>�0	>���;d�=��=�)Z=!\�=8�s>�q�'b�>�}껛����r�l� ��Lc=�����a?,9��⧾�U;�U�.Nv�?�?�U?��>��,�d0����,�:��>�<껒������z��BP=I
?�:�%�l����Ѷ��R?�>ew�>Ȏ>�����\D�4;���Q>���>N�־��=�y>z�(?6�v?�>6?��=}d�>oa>[ӏ>���=M>:?Q>���>��?�9?l1?b��>���=\�`�=!�:=��>�0*W��6��)q߼a�$��e�<	{3�~oD=��w=ݟ
<�_=��B=��Ǽ��;+>�<P�?r�H?r[�>�#p>L���� ��*4�AU�TF>��a�M��>C��>��?�B�>�A�>ko:����]d�<"־N�>�"m>�S�=l�����`�>EVW> �?4pI?�/S���	t>�=f�>��.?E�S?tl�>z&E=s��:��&�ѿb���(�h�y��Κ���W<��=�p�<�Y�>��h��5u=�-�=��@>��=r�
��\=YdE>7��>1$?��J>jL3=���b�e��9~���o��=��-�]'y�ak��\X=�ݱ�Ӈ���K�_ ��0p���༕�|=E�?:�X?k�2>:�Ƚ]��MP_��`�ae�>�r�>��:?�I?۸<~w6��K����]���*?�+�?��>8��nE0�_�0=��>���<Tw$>l�$>���m��J�}=��=��?�{.?�Uk>_�m���y�Z���/�W�>�<%�ϙ�?FC?��'�.��:uX�y�w�*� ;>��9����ݾ��C
(�փ��-���8��q>�}�>\�?ht���L�=��;ec��طB����֌="�'>��\>Ӡ�=�%:�SMҾ���ZѼ�)i<��>��?�Y>?o
>ބV?[م??�?�?N�>�d{�o�	?�����>j=?e�G?b�?� �>�u`���?>aB�=��꽷�}�9��=O&�=���;Q��<��$>w>�d�<>:=4�
�i�̽-/��Xp�;S�Y=�J�=�=@=�;�=�1>�?gn#?v����8 �R����+���2�>��;>�zq=����Rb�� g2;ڭ>Y�?3�?�>�ċ:]���ݾ��(�SUp>ʕ�>y�F?E�N?r�����-�9����Ӹ=��>ch
���� U����ӫ$�J@�>9�>�%��=b�>Ht?�6?r�0?X���F<���q	h�i�0X�>]��>1@f>��9>���fy��݊�p>���q3��Up>_&��Q=����g]��Ky>aj�>��=i��\�H�G�o���=*�B>�f�>K��>t��>a�f�+=�ƾ*l���D?#���wY0��� �f�;���=[4 ��۝<�}�X�>N���눿�d���_5��M�>�l�?R�?��b?*��@����S>&={t=��f>D8��4����i>b]�>�m>�d���B���K�=`�>��>s��I�;]󾬠�gݱ�jUS�m���4龕jҾ�wѾ�=�����m���&�+.ƾ:\(�o�d�����AH۽�LS�p-���Gɾ$r����?�ߌ?FYa>7o>=@�C����$�4ϒ���W���M�O�ڮ��|���ƾ�+��8,�K�3��`5����/�>y-k�6Ґ��5w���/���S���/>5*?��þwp���-!��'��X+>Ej�=�����み����p�/��a?�
2?4Ѿ"B�RL��l=���>�5�>F2>�n��"C���j>^N/?<t-?�=]��(��oч�Y��<U�?H[�?'(H?GIi�1�E�iK
��Eg��a?��?~��>K��� �˾��[��>��:?�R�>����r�:����>F�c?��e�'�>W*�>`�>�[?�/¾��=�㏾�X�Ғ4>'7M��읽`]F��b��<ݳ<��>\j�>A<�ٖ����B>��ʾ�UI�,�]���'�R��ϊ�;C��>�f��ǻ1>�ԍ>B�z�V8%�?<��؂|�~�����H?�?#�d?�cf?�8��b;��~b���.=-?sj�>�p�>���$>$l?�����Dw�dB��24?�]�?��?��U?�I�n������8�����;��>Z>�1>�V���d>�NK<e�G<�=Ϻ>�X�>��N>?��=ٙ0>�)+>���>�yx�F� ��ߣ�������6���Ҿ�������d Ҿ��d������ɭ�N��%�����
��R���I�	��<�������=���>�?�1?C>��>��P�k%Y������<B��AJ��E	��"�ץy��y��%��; �T�T��z�;���gA?IH=S�)>ۍ�>�}����;�^c=��g>[dv>Xi�><��>�)>ȫ:��p>�4�=�Wu>w�	>�Q�>�(>ү|�kʍ���#��T�=a1F?�+�x����B�M���X=���>��?k>w?��ߔ��q�m��>�<�sY�v%����ĭ>���>4��=C��<d6��+�h�|��K��
ɴ>��x>;֥=�[��CT�>�*�!��>�o׾�1�=��r>��'?�
x?��5?���=��>�b>�l�>�0�=��G>N>AW�>��?��:?�1?^��>c��=kC_��=̵D=�;��,[������o�n���ɝ<�;?���3=��v=ϰ/<	�h=S=H)Լը�:���<r?e62?Z�>�>����k1��&V�>�\��T>�Q�f�	>�<�>5*#?�>��U>�$������9����}�>�'c>�x������� ��8�>�?g%1?6�?�L&;�;��R=Xd�=�S?��?�< ?E{>p�>��/��)��F�8�%�G �.�
�g>�7:C���ȼ���>����Y�<�zo>��>T�>�[�=D�j=�Pj>�\�>��>���=��%=�$%����)�!�)�z�Hᖾ\��&��B��=�=;<;���t 2<ԯ�ih4�: ������H?�$/?�Ë>a=�1�S?M��³��?��	?V��>�{J?)S�>���9I��kp�m{�
�?�9�?���>�Q���.=
�Y	=� �=r,>S��� _>�M<W�a��$�>���>�6Z?"��=����zv��	��e�����>�~l=�.?�7��?�c?��ԾI����ξE�]��3���t>���.㋾�U���s ��\&��PZ�;��s½�;>���>��?x���c�2��~����~�C��� ��>c�%�w(>�4�=�6��i���9��r$@�t�>��>��?6�>)�?k�?4?Y�w?��?�?N���2M5?�_�<��b>LV#?�wH?i�F?�J�>x�<K�=�v�&�0�y�c��1��}�>�#�>�(>[
>F&E>#�`�]a8<��#�~�=%��=®K�U�=�>�<NA ��_>N��=��<>+?�,?��k��v9��h=[L�]4�>K&>A�S>�Z�4�	���7��KS>?n09?z�>I��7Y��S�1�	��P>��>I�[?�8 ?*'�����<�f��iN��?{�#�>�J�c/�����2T�����ۋ>��>�'��Vi@>�n?��S?�?p~A�@ ?��w�����&��=�W��ް�>��>)�>�:<�$�N�Ś���x��"�T7=�A��㦼��=`)ɽq��>�<H>�"�<b~�CQ�N�7�'
����b�1Q�>�1�>�o�>��>Q��>�ϾRR���M?�뾏�l�9w���¾t��>6as>�<p/��,�"?���놿�莿�����B?���?0>�?C?�Ij��f���c>�en>(�>���{ �?�k=�o*<he�=,N(>�Ⱦ�������<��>��>I���v�񾐟� �k�O+ɿ�BX�����_��������ܾ��z���;���n ����6�����>����s����?���>���ɸ�ֳ
�O�?S�?N�>>����*2� Z8�e[����a}�vL=R3��c�ξh�������������ě"��=ɾ3u��3��>TPY�E���U�|���(�a�O=>rF.?�ž�!���t��/g=�%>��<s��[�������y�ÓW?�:?�2뾦R����MO>��?���>kR%>�����;�)ё>�33?Mh-?�x���&��j����ޔ��{�?���?�WD?d��'d=����Խ9>	?5?�z�>o�e�U�ɾ�7��*?RFA?� �>���́�[s)��x�>I?(?��q>2��>�6�>	Wؽ3>l�����*����M);�>�q�~��;��$��R�>6"�>��>�pr�Lﶾ�3>^��%>K�����43������q&�j�>�
��\������>iچ=t�)��岿P	��h7b�ְ4?�?�Dg?�d?C����*�����~f��/�9?V�?����Լ����>���>OR��&���i2��8?�-�?�?�Pu?F]���ܿ��������w�G{C>��=2�=4�M���H<�i�<�R$=yS�<2��=Z�>�X>c�@>1G>��S>��<>����������%ʄ��F���S��4Tz����Ȁ������uľ-�˽&PĽC�<��NB���� \��ɏ���0�< Gw>|Q�>ί?vބ=(�t>�b���+�P�޾����<7������$��mr�<E�p�	T�YT��c�w����߫\?#� ��S�=x��>k(���"�=]v�>m�,>���>&��>�F=���=�A�;E;�=@q}<��k>��<���>����0���Gs��HK�d5���(�`�U?p5[�[y��+S�i��]����>��<?�S�>���ր��@$=���>�:7<ʽ�!= ����=}��>a��=�ݰ���=�v���BS���E>U}�>AQ�=%|��|1��������p=]��>�{־8o�=��w>��(?��v?B26?�4�=��>qub>{�>Ғ�=L>LQ>瘈>��?��9?E�1?���>j��=�`�(T=�/8=�>���V� ���7�}G%����<�K2��G=��s=��<��^=��B=�N¼���;��<�{�>I6?��>ێ�>H�>��@���G��q�X� >=h���>׆�>��>���>���>�,K>����̪��'Ͼ�-�>G^`>+e�k�y�$�����f>�(�>�cI?�2?�����$|���	=���=�I�>�D ?�K(?;|�>��$>��ǽ��XHӿ��#���!�L����8��~>;α=�L���+��R,�K���j-�<�:\>~�>�p>0�C>?�>Zp3>L��>�JI>v3�=�/�=v�*;< =:��N�BwW=�t���9<ɁR�툋��üGE��U����UL��E����tἙ*?ѝ8?�'�=��>��N)F��&߾�F?v�~>�6Q?��?o��<iξ��E��e��i2��;?Hw?���>����=�s�jx=��=��>���=F�L>6��=�툾�!v>J�#?��:?95�>�W;��1���x��4������>n�W=,)���ۤ?��I?ܳ�g����{0�N�S�Me.��Ŕ<�������h�ć�ݝ'�?���h�a3�tM>��>�	�?g����I�=��>ߠ�\�X��#��.��9�1�<�z%>����ڪ[����<پ��g8�=���>T�>݄X�)��Y^N?��D?n�?��'?��'?;���:>x+�>���>�y?�?�<? 7�>{���2���}�/)�����큅���=?>�=�l	>��i=;>���3ۨ��1>p
o=���d�̽��0Z%���=6ca=}V�=S��=�|?�-?X�ž�������m=�c=��=�Ó>�����i޾+��=��>��	?,�8?#��>v�7��z����բ5�S3�>�?�2?��1?G��2������Pܾ2"=��$�>E�ϼX\E��3��C���;��6�>��>Uə=$�f>�x~?V�@?>F!?���j�+��*v��*��8S�5�����>D�>ϒ�=0־~�4�'�r��^���/��c�R�L��<�<�j>�>`~A>nM�=��>�Z=����5ҽ�u<���U�>'l�>_�?j�O>El�=���`|�$nJ?1&���1�{�J���9���Ē��A?�o�_>�¾ ć�����r��?�,�?�p�?��N?�4&��yz=@��=v//��M*>tx�9�]���/���'>�@�>��K>�U��[����Z>���>���>�iû5��w����c<�Gֿc�(��&��Se�������B�7����XڽnX�?��u�����%���}2���U��[վF�R�t�ˀ�?�g�?(��=
AP��I>�p0�B��_>Ѿҽ�{�j����θ�R/�|���D�h��= -�p
�J���yM>C�]Ǆ���q�i�&�e�����%=X�+?��{��ž�����g�=Iy>
"˼D���R������J!�)�o?�9?A�о;�$�T� �>Ӿ�>�(�>c
>3o���A��_]>%R)?`&?�Pսm,��@��/��k4�?��?�&l?�	ƽ aC�/,�����}�A?p:?�~�>\ҋ>���>V��X�Q?ֵ�?�O?X��ۏ��J��I�>r�?��g>�ef>�$�=����T��<��U=�z��5t<�ǽ�����CI�!P��dn=%E�>LY?`#�>h���OE�i�>�͠�
ZE�ϞS���C��_���8����&?K%���̉>���>�oV>��X�V)��XЄ�K7t���H?-��?P�M?n?nA,��(E�N����Hg>X.?`��>$:�<��쒥><��>��l�y
Ѿ��??���?���?$�j?�\i�g�׿�����2���H��<zU(>Lb>�F��ފ=> �z�k��8�^�=���>�bb>���>㥉>�_O>' >�����S$�WȮ�������X� �}u�Cl��D�֤�����Ⱦ����&����^N�Uo���0⫽��=�c.��m�N>��E>;�>8F�>󯽬�>IEf�	P�}�I�E`U��2�ņ��z��Ϧ�����4�a�D�4��j5��$Լ�s��"?z.w��!���>���=Kj�;߉>6!>�X>�@j>��j>�i1>6�Ӽ#��=p~�< ^>���=Ř>a��<�
��Zb��b�#�y��t����]??�J�ۖz��0����P������>|�?jDX>T)�r���}1t�>��>~��J�U=f����.�E>���>���=V��� x��q��|v�p��=�+�>�B>W���x��\
�'��=�D�>��྄i�=�a>�n(?q�q?D6?)��=Ƽ�>��C>���>p��=��H>��v>�d�>��
?t�'?s�5?�!�>�0�=F�^�|*�=�ń=|e��N�RY̽�������ش�(��[59=΃.=a�ީ=ѩ�=����n�X<(�=&c�>~�??\��>���>�2�*+J��QI�t�c��u�=��Qu�>�՞>�@�>\5�>�J�>zc�>�{x<�����ؾ���>�Z>>�e�
����L��wU>N;[>dQ?YGF?�7�<9sJ�p��=k3�=��>���>^�&?ͮ>��%>�ܽ���y���0�㾆P���Ek��=���<����@����4�����
B�ӊ���T>R1>�>{�>\�K=��=��>I�>M3>E�>�'=i��<':�<����tM�=_ $>�O�<G�<��;��b/��1�O^}<
b�5�ŽT��"}�>D?�t�@W�<���l6��G^��D?l��>C�.?��>���=V��]z�e�~��z`��/?��S?��>�R�ێ��2V2��d>P#g>y��>�>�j
>Ę�>���`k>�""?�e-?v�>�ѿ�ɣl��Ė�\$�T�-?d��V5���?5@?�U��K¾�<�֖3���������	R\�0��I���Y����8Fо�����>%?st�?�ߗ�z
j��AȾ#Y��>S���o�ļJ>2ё;ғ|>�x2>�6z��	�O��ͽ/h�=�J�=��>A����*=m��?��C?G=,?�W�>�Q>�-�0�>�J1>%1%?� ?f�?Պ>��>�s�qJ<������𧽗�Q��I�Ӯ�<!n'��ϻ=$��=o���O�<`��=��M=�[�=!B�"�9=#o�<s=���<�>�`>�O?��!?z�7�<wQ��Y=c����>7r�>�>ېs��$��c����=�0�>'Y5?[��>9"��'������0��+>�q?��1?��?�O����>C��!������ֿ>�/9�aL�������n���K��v>D�>�H�;1bV>��~?q�@?�0?1��Y5�j/k���,��颽���<��>Iц>|�G=�߾�8��m��T��^-������A�͊�<��>�1>_�8>�ʶ=�O+>�ٔ���ҽ�ｍ�H;h
���>���>�?�J>RU=�l��O�!?J����g~%���A=�m���A�}�\�� ~<	�?�H�����:Ҟ��F2���>!�?ŵ�?S4I?��ݾII�=X)t<�;�<��>Ř�>�/���3�� =���>�>�>�ݾ"ѽ�%�O>#C�>7d>}�K�jy��������ſY1@�
�ܽ�b���ɾ���/z��&ž��F��E��׾ō��!h��R��_��dJG�]��hN���Ň����?���?�f�=tf����m����SvY>ȃc��G�y�f�Q��m����FǾ�ξZ3�Х����?����>�	�����r�`��.�"��=;$>Y�?�]ž�Ry�Y?�6���Ձ>�4�>��ü[=x���������m?�R'?�R���GԾK$����}>V?���=�ʾg4�`d8<��M?�ci?-�W>So��hx��q-&�k4�?�4�?�rl?�ӄ��NV���3����;�R?aw)?�ӱ>h\��`�����^�9?|�?/H?$䕾F<���S>���=�v�?i�_��?�>��>���=)Fa��]ҽ��8>�l�+��=�θ=�`�g����设 {�>�u�>�Ȅ>���%>�~�>�
�!���菿�:F�[~>��ʽPW ?�P��A>~�=�U�>S_��ψ�tÕ�tC���)?�u�?���?��&?h���3��"_�>��>�&n>�.>P�t�����>�o> �2�p����)Ӿx0�>h0�?�0@_>?�������:���u���SuN���e:� ��Z��>ʮ�<u��=�U>0j+=T��=�t>%Y�>�V�>~�5>2{1>V:f>�?>�	�����\䩿�ꁿ+9���0�B����Z���,��/}�`,�mGT�ϛ��lx�� �6��o��n���D���<�����ǽ��?b�>��?~��>o�$�6=�ss��HW����� �r#������־�%��D(>�⮽sAž��C�J5�=�?�J>t�1���?�{�>�\(>9K�>	F���L�>���>L��>�E�>Ar�>Bz�>K3 =��=Fd:>�{>("�=_)������u:���Q���;a�C?1�]�@i����3�op߾����t
�>�?j�S>��'������x���>�G���b���˽, �>Z�>S��>���=>�Ȼ�@���w��_�=���>U#>?`l�����>����=���>:|���>�ބ>�=�>��?��!?|�'>�?��=��>��=u��=9�>^L>�#?��8?�?�9�>1�>]�-������c>��¾�=�«=	N�т�=K:��*+>>�F�J����=U�.��q��J�ս𢗽�b��w��>��??���>�V�>�X8���8�+;6�q46���= 3�;�X�>{�>��
?�
?���>�>k�ؽ;�Ծ��߾��>�*>�}Q�WOj�%l��C^>w�>��X?|2?��=|8l�W��AM�=1��>�d�>�2-?�k�>�?G>�����#�Կ�22���A{ �Po�g�*=�� ���н���TSU��v���`=�ti>���>��r>n2_>��I>�/X>g��>�R>�v>w�A=�`#��BU�����;�D���
�����D���
��{�������˼᥺�U>��[7��$�?O�?�f�H��:����vH�;�>���>!	?V�>y��3$���]��|K�%�2�M?�|[?ĉ�>6xv�N�L=��D<�^ü)[?<��>+%�=�kn��6I<������=��?��?^ʼ>��g���z�E`m�Y���$>�(=V)����?�Gb?
m.�@>�e��!sA��Eo��. �aG_�:`����8���~-����'�������0�ʽG��>V�?Ŭ¾p/=�h{�)���'F��h{�XC� ���=;%)>p=Ӽ>�Ѿ,��t= �L�ξ?�J�j�@>��>5�?��>�~5?�=?�FT>�lQ?O=(�	?�`�=�c)?4?.�7?��3?w�W?��=D� �Ŵw��u^���q〾Q��<C�X=S8>}O�=��o>��">T�<�ї�wq�<zߑ<�.M��L=�� 	=2��=v7>���=��?K�%?�̽��"��h$�r�=�O�=_�F>�E���U�G��;��b>�n?I�1?��>[�5=Bt߾)Z��z��*ٴ=x�?2�.?���>+<��=�t�{v�(��=�5S>_�|��R��$���!����ɒ�>+>.��=$J>VC�?{&?���>����	��aڐ��f��Bӻ�ހ����>�m�>2�>��n�����rv�;�Y���a����������u�=<�<��<0[�=���<yW0>����������>�u>�>�?���>��J?�	z>�'S<�g���V'H?9����%��������I?T<�*y��$> ;�I�M?Ӓ	����ѥ�c���=��=���?���?}�z? �<%JB�,V�>_	�>N�|>v�<��K��Ё&��M"��[�>{��=��w�ھ����&>�>Ch�����z0�����Կ�`\�;��o������ �B��Z���jE��þ6`��� ���l�����eɽ�B��w�W�m�z��庾�쾶-�?�?r�>�P�����	w��/��� �����TZ����Ӿ�w�jQ��߷Ծ;�>!���M��{6��@�9��=T#~�'M��$��&m��(彫��=�r?P�ȾR�+��c/���=�>E>���U#�*"u�?v��<]�=�q�?f�n?T4Ծ��\�Q,�/u*>�]?W�>�?�lK����c�>v@;?��5?"Ù�[Ύ�%tC�Ҵ����?E��?s�??�pP�IB�m�����T?�|?�F�>����̾�^�`^?[�9?+�>�e�<O��tG����>�\?ȒM��a>Ok�>KS�>�@�c0��t�&��<���p��5)9>N���H��M$j���<���=��>�z>+�[��O�����>�������w�����=�7>�!b�?�H?ޠN��%���D=
��>�'K��\��	%����=�TL?b�?�?��?�I�n�<���>�?��]�J<&M�>�O7>��o�L�=5-�>��#�q���[{c�?@�?�u@��@?ݰh� 뽿��������T��g�;$~a=�F$>%�޽Sv�=am=)��{�A�ޭ�=Gw�>�TF>v��<�@>�*>�>e���^� �����������f� �
�\������E����񳽐q3�����	����Dq6� &����`��_����䏟��)>h@�>L/>� ?X-�>\��=\Q��������
#���྾�����l+�#����4��/��]�j�
KԽZ�6��-?�=��=x��>�F(=VE�=|L�>�;�<�L=d�H>x�> �>��>+F�>`t>>���=y� >�f>!|`=���,-���><���Q��X;/�A?+G_��Л�q5�a���ɪ���>P�?L,A>et'��Z��@y�v]�>�7;��]���ʽ�f��ȇ>���>4�=�G���Z?�POv���߽ĺ=�Ņ>u>n�E�6Z��� ����=�	?1��r�>>]d�>Cj�=�3?N�@?k��>�o�>��d>	?K��=���>��>�t�>�?�w?���>�J�>D<�='t���b<�%>��6�NGM�����Z�p=㽽o�$>�Z-=��4��{�=�>	>߀�;�p�k5ʽS����>�p?��>w{�>]\���T:����>����@>�Bݽ��p>��> p.?f>�>�K�>4>f��n
��V�cf�>ga�=��D��Ap��-�<a\?��b>��J?*"?��=�z����> �y>;3E>諠>���>p>�>݋�>���=n��iqĿ"	�=1��>о&�|�����%� �Kø�z���hZ��$���g>l�>��6'8�3��fhR��"�>).6>��">͎=:�?>�n��2=�?�=7鋻%^���=���=�Sk=��4<����>�|�=�ǔ=�����>�?�&����9��<Y��eQ��\�>e��=�~>R�>��L>, M��a���>�v_��?v"�?���>�ľ�ע=[��Ã�,�?}�0?��>��[�u@�=ļ� }x����>��a?<9�>����>|��{�3���I�>��<>Lm���?kl?�ܓ��d���'�\��A�J��榸������о�:�ql��n4�žn�����>���>s��?2���~_�=�@�(���]a���"��h ?�m�>��>/Fa>uc;�s�Q�#[����[���9��|�R>�>��>K%�>���>�?�>}�"?E�7?G=N�?A	�>1��>,��>m�>�}!?3&2?�K�>��->��y=W<�j�]�
[J�nIv=��=G/>tp=�N�=��ƼC\0=��>��z>�H�<�c�_��=6������<,�$`>�! >�?6?,߼:!�=�$��q��=6��="0q>���;&q���<��>��>Z�0?t5�>�׈=�a޾�z�4lȾI�=K?�?���>�U�;ck_=�M���\�R��=\�>Z��`塾��ž���������I>Hʒ>;�,>�>�/�?=Y
?��5?W/�;a�m�lp��8��l��>{��>��\>;] ����>�8�>�Y�F�_���@�wx��9�R�1���#1>z%>�t�=x&�9k��3��>ɽ��s�d�V�̷H�)<�4��>b�?�-y?��->�� �7WܾS�$�^�A?~������K����g�՛��lE=:�>����՟>E3���Hh��iǿ�`�m�=7�?)�?��?�4���Mi����>���>=I>y�������oʇ=�Ƈ�5p>�I>8�W��k��<����R��>d��Ȃ����*��HԿ�A�2�<�nྦྷ2�)�w��m�Ѿ��ʾ�@�ݦ������#[���ӽ�K�V��l�����U?reW?��=���]t��b���޾2=꼰��Pþ����3��.��$�۾��̾4B���5�m}�
s���g>��6�+L�������&��ʿ�=l����6?dI�Wi߾��`��>��_�6>�z���:���e�񹴿�?�ݏ?ߢ�?���Bq���-����>�S2?�O�>�%?�ܛ�]�Q���=isF?H-/?f�1��Ė���R�d����?�+�?g�B?ЪF��U6���ؾQD���>��?O��>�㑾,����5`?��:?kŽ>��N|�q���K�>l�`?�'.�ZK>��>�}�>�i �6匾 K�]_��������=�1��V+�Ǣ_�������=9��>��>��D��C��(�?o'۾����4ƈ���� t��I��"B??�D���=�ߤ=
R>O�Z�*x�����<�	6?;E�?9��?�X?%ץ�^5����8>�ཱི��=B�=�]>5��dЋ<<�"? ��&����f���?*h�?j�@���?���]U�S��=Ω��=���>N#=,�>!��o�=;8=e�󽠍��OX�=��>�<>�j�>�<>��C>�/>�����#�h��+Ԉ�wl(���'�W�6�C�����0��]*�ږվ�̾F�'�� �N?!�o� �Y�ؼ�����R>��>u�>%��>Z��>�N�=�l��v�;h�kV��:z����������6����Z�ӼI���k��ՐB���A?j���Ȳ�V[�>cwu��xZ=3O�>������=�9��Ct�=�5?E�5>eф>��>X�e�L�2>%WA>��=l����(���v-�Wߦ�⫼��G?j3K���Ǿe�V��t˾�n��	I]>���>G�9>��;������z�	5�>�����|��
w��>RϮ>�#�>޴>����^�'�ʾ������=��x>���=Zk=⵾ �&�A�->� �>��ݾȑV>��d>7a�>�k?
�K?�J�=�!�>�Ï>��>���C[h>Y�>�%�>v??l?�?�~�>�� >|"��E�=��|�NŊ�mOཀ����4-?=�������9h:0�e���=e1�<�
,�)�<��=Y�=d�?&�L?�a�>���>߫����G�)�1��D�]H�<�T���*�>�+?y8?]�?t��>�l�=:��;��پ�4.�k��>k;>M�B�=;^���G����>�lk>M);?�F?V�}=<s;ɠ�<Uk�>���>b ?��>$�>��[>{�P���Z޿������q�j�P��?n�<U�
��6?�ε=jmV�m5��A�=>7/>�΄>���>���>S	$>��k>Zx�>�E7>��==13>�9�=X���Wǽ!�J<�_K�y=hF=�D�;��:�vڽ�UE���R�粺��빽���9�?��7?ۜ?�?<��H���<�>_�� ��>%0�=��b>e�>�$>�l�t�*�>�����?~mz?�>!���7�=	Q��I�>�^?�-?#E�>9y���[	>4ʤ����=) �>��h?i�]>WU�=fV�����h-���>�%G=^D�D��?#;?��о�H�-M���.�]h��sO�5t<�� �y����$��.�r9�����g�D��0�>��>��?خ��f�=�i�zՎ���~��?��\>�#�>�W�>�i�>�B���"�,J%�3�����ѽj �>j�'>[v3���>Z�'?H�?��K?��W?z��=~�?���>6��>��>�$?�z%?/@?��?q�0>I�<� �΃&��D�v�V=Z�����$>-�3>u�X><��=�c�<SJ=�h<�N����d.���=`�=78����=�s�=<a?�&?\T�/C@=Mr���%��<���=��*>[�V��p3�{	�=���>��(?}1?�w�>-t�=�.ݾ=[��̰���Y=0�>ۙT?�ս>��=#�>Q=ܾ�����J=.�>���Q����̾�Ⱦ��=�$n>�Ò>5xQ>�k_>�z�?���>N ?�S���a�5��&R��;�=�AL>�)?�>XS��V[�Z'���ra��sg����։-��:Η�=�7�=:���;��wA>wT=�ܾ�'d�5��;Gu>MȄ>G�>�T�>MTG>ƺ=N���A�|KO?������3�޾��6h���T<�9�>h���>���S'v�vy��1�D�MO>���?�W�?�ی?g��J�nc�>��>��>�Vҽ���Ք}>�����Vy>b�B;�Re�� G���L>��=aϹ>]R��[������Q����r@+�{O�=�m޾�&Ǿn��ã�L����"D�蟾:�����!����K�V�_����p�� e̾��۾?�?\�y?G�5��J��/:#���A�k�䃘>mf�s-
�b��M�<b�S�t0���K��O��:1���5��i�]B�>	�W��߷��s�� Pa�F�z��q�=��q?9žvI��ZĎ�3s>/�=���;) (�FLw�l���P�l���k?��B?{�����'�"->�5?�16>�>�Ӿ0*m>���>��C?R�-?���E��������J�?���?�@?z�K���@����\����?O>?M��>{2��$�̾����{Y?�2:?��>�6��=��U����>0�Z?+EL��b>6C�>��>����ْ��$�@����~�K�8>`�ԻO5��ng��J=�n,�=Y��>X�w>\�򑭾��?J��ъ��`��ח��Y�s=7�	�&;;?�`,��/e�§�>T>�>�1��o�����=�B?���?���?�~?ݰھ��}�x'X>���x��>Nw>(Fۼ/v���>���>��D������01�L��>��?l�@��u?2���ڿ���]���㿾�♽��}=��>g��=��>fr<=Ǘ��Ad���o>ϼ�>�>7�>#YE>�{7>'�V>����	!�����,-���Y���5S�����=!�޾��S��q��޾���~M1��8�=B1�;79� ���5�L���!>:M�>�p�>�@?��>�S>�/	��3�7�ҾO'��*$�L�*�O���x�"�����B��»X�Y�A�Ƚ��)���"?i��=��>/@�>�n�	�%=C�>C�(�>k�>��>u�?��>�Vm>�!>�7>�f�=�A|>�j�=v�������n�;�?`T���^;�A?3�W��*���5�K��J���9ǁ>f�?P"Q>��'�/���ԣx����>/E�\af�V�˽�%����>�|�>O��=���y�%��/�P^��0��=�݄>_>y�?�r���$����=}��>�{�2<>ٔ�>�\7?��?z�!?W�s=֡>ŘӼL0�>V�<=G�$>��q>�>�?�03?��'?>B�>�>t��0�Q>\�#>pX�����>�.�~�����o��=j,���-=�>?�=6@=ZP=��5���M���>�";?���>$��>ـ���&�n;x�ĥ��)>�A�V5�>t��>��?\j�>���>.ܬ<6�;���߾&����\�>G�\>Y*A�	�t���h�� 5>�X�>|9<?*�M?��=�(��E�t�=m =T�a>��?�?n~�>Nv�=Yq�����eۿ!�CS"�ڧ��Eʼ�"> >���=�]=�!7��v/�Ǔ�=C+�>���>0�>ۋO>�q6>A�`>Ū�>IU#>�Z>N #>��>>E�x<OO�4uý���5��=0ة�T�
�!����s�2�	޽��~��������N?�?��a������I澧��~��> ��>���>�>�>u�y� 2!�K{�B�U��!��	?��h?J��>���q�>sʐ�7�Ｗ�?�k?N�>���9=Z�о:�==X�>B�
?�:�>N���8��2ځ�Yr"��,Q>bX�=S����?�[?��ƾ�!�x�S�P����<�M�\[X<Z�i�8�n�;��`�+��� ����΄��|��'��>��?�O��+�<����"��3���3�����Q�n��C�>�M5>�d�<ɡ���ꬾƼھ�Y���ս	TO>ϳP>X� ?��8?��^?4�D?���>��Q?\$�@�8?$R�>O�1?�v?oA?��+?�r?��=pv�>��ӽ�콋�>���p���һ��ֽO�>�u�>}�>�N=zJ*=T��<W��=�#�����o$�>p�!=��<h�="�>��>U�?��<?�sf�V����_��F���՚��N�>y�>2�~������=�C�>�-?�>��N�CM����꾻�K=�M�>�e5?�B?<��ݩz��x��O�j�M}���H>���3�)��Tξ?D�}w�~��>}>�1�=��>��}?�Z(?��?�����-�(�w���F�ޙ�>���=)���9�<y��=�8�*�
��b�%�M��G��dƾ���r�=��j=� >���=)���r{�>rQ=�+�=�-�>&=�u>>B�>��(>et�>�Ox>�X�=�,B�8�}��U?�*��	�8�]���}���?N��+�=�5V>#��*�>���������Խ��f|�p��n�?١�?�[�?GWR=$���-�>L��>i�>כx�G@;��)>�}H��o�>6Tt>W	��־���=Y���>-�Z��!ξiQ�G���ְ�� M�$[R=HZ����7�I��8�Ӿ������ھ���=!s��,h��sB�K�=�h����VRǾ��ھM��G=�?u�?�����W��3$��5� � ��@�;0�9�bA���m���ý�>��<���%꾤�վ�S���M��P1���>��z��1��H)���������{5��z??A��-�Ծ�D�;�>Zǅ>z��=���g�����^d���m?WNg?�1쾱,U�������>��D?�ø>�?Lڽ���zZp>��[?S<6?�b�jk���[K��u=��?�U�?��??BcO�tvA������
?Ks?�z�>A���};���!�
?	�9?�z�>;���p���@�N��>�_[? 1N��Tb>ܴ�>�D�>B��5���N�"����b����;>�n�Ap��i��>�Gl�=��>:Jx>��\�����Pd ?��渓��vV���2�	��<��6���F?++��B��<�<�ȓ>��:��Z��X7���>G�W?kh�?3>�?z�#?�̾��/�a� >7[�=[�P>&8> �=Z�I��2>v��>�����������>U��?u@�W�?�\����ۿD��ʥm��'U�͘�>��5=t)
>��O���;�"ͼ�!�=q������7�f>A�N>�_7>�*�=ƚ�=A/>�H��ݥ�����:��O�"�W���]�U���$)߽R$����' �k�/p`�����f���z2�����X�Ⱦ��n=��>BK�>��?�]�>�>>.��L��t\��ݬ��В�n������5������t|�>�	{�mi��۬�d�?��e=#���8V�>�U���ý^�>+��=JN�>zj�>�zy>3�>���>;�#>زh�Յi>Q
>?��>e��>x�h��(��<�O�mR|�Q�O>�Q?�疽�(�L8/����%9��X��>PH?C�>���2���}^�-$�>󫇽~�a������򉽤�>�S�>��,>��}=*�<:Iu����P/�Z�>\#d>����8Y1�\���c�=�M?����·�_�>7>:Q�?FO?�
\>��?n��<#?t�N>#�+>q�>o��>��>g?ݍ�>�b�>��M>����� =�1>%���<	 <`L<�b��P��=cPp��*=L���Ѩ>�&>�=zj{����~o0=Hz�=�@�>�'\?�~�>�'�>������i��-�Խ?Dg>�����>U��>ؑ?UO�>2`�>�H�>+�����F���>��>�kI� �r��5���c�>m��>�0X?*�/?��[=�W����I�,=E=��>5Y�>��A?���>(
>x�Q����\ſwB����>`t��כ��`�s�67��
�k>�J]��?�?�i�M��>��>��:=�
=�\
=�$�=!v�>��>�H�<�9�ge!<=�=(��r����=��,;h��w\-=iM�<�ź<9Ù=iV���)�O��ň�=_�>
?�'ǽ8U ��˧��&�_o��9�>�X>�9�>\��>0.�9
!�m_g�Qo\��b���?�,]?(��>��ľ�>�o =��=a�0?;0?_�>ЉW��ҁ��_�X�L�}g�>��B?v��>��(������鋿��,�P�c>7n`����?e�c?/�ga�����f�X�T�Y�w�$�'�PZ�=�N���.��6�ː����ʽT�]��=b�>�Ъ?E�쾐}N=zs�����F`��d̗��>�]�>gy^>˗>��N���C�u��/z�dWL=D~=J�4>��>j��>���>��
?Z�>��?`�ü��?�>��?��>���>�(?'z?;�>�>G�Խ�$&�꙽�셾%���R�;v�b=��J>_v�>*7��<�ٽ�=|.>��=�>U�(<(�l�ɞ^=��=��>[<=ݍ
?��R?L� �$�����+�C=8��>��>���>PT>�	^;!����=M;?SBQ?߭�>SE�=�۶�L;��6���Nܽ"��>��@?���>���#i<����U��Rr�<�G/>R9&�ꙕ��hľ�Ѿy�Խ*9>�>�>��>S�D?W�C?�c?F�	��S��ؐ�`�R�&��>�T>�Xu>��>�(?C������M����N���?�1&�����$�&>��X>�m�����87>ѐ_>��=�&;�i���~j=�V�oт>K&?:?.?r��>�'�������2���*M?��龩�0��Gg��2��
���o�9{�>j����v|>�U��g	t�Ӵ��!n��Jݽ�,�?���?�?�󷽭U��?�>y��>�Q>�4_�n����>����{=�u�>�<�<짾e���+:S=�t>��{�^Y�'����y��\7����=�/��l<�dN��(߾/�ԾO�Ⱦ��=�wþl5н��|��_ =6��N�:� ��&¾�!�� م?hW?=8��sy ��
�P;��f">�Vi���f��:W���3��(���e��_<��t����C��6,�>�����\��4����о�Wn=XM�<ZI6?� Ҿ�"��s�~�?�6>��>��8���{����i� �
�?�!`?S���a\�#�y�<�>��?A�>��%?u��ľ@�>ق#?0�B?�o�ۙ��o;�n�o�6�?�E�?,�??��H�DBA�z��"�ǲ?�t?q��>���ƾ�/ǽf�?�7?>��>����������>��X?�K��g>�_�>Z�>���A���e��0�������,>OL�����Uf��L;���=�?�>�As>�^�4��-\�>h�Ͼ�h��h�ؾ��?������b=t�z>���wK�>ڨŽ�F7�YQ�)����P|�H����5A?���? ?�]?����$M��ľ�ٝ=&�>�F?� �>��л��>q[?� <��^�RJ���K;?=�?���?&�H?q%O���пP��_ɾPe���&>0�N>z2x>����M=��Ի�R�<�f�<�W'>�/�>S1B>ۺ,>�2">,�>��=�$���/�\K��<p��.*I�Kd*���	�!,���2���s��������[��= {�S�ܽ��Ͻ��4�s��2�p�8n	�:{<]B	?�X	?Zx?T��=�w�>���m���B�����/7������z%�����-O�`��1о����a~���T���2%?l;u���F=���>+*���>���>.rj�.>]G>`��=>>�>�c>�c�>���>��#>rƚ>�_:xȃ�����#�2�?�����=��@?����斋��@9�{�𝜾G�>�e?C"�>���@Q���(K�~�>�2Ľ��P�*��.�z\>�ѭ>�v >jƈ�$�L�F��Q$n��$�>B��>�ٿ=ӵ��򵾷U�W�,>:�>�Ⱦ�];>b�>b%?Jr?�0(?`ۇ=>�$�=IV>:�=8�>,\:>�w>�?��<?H8(?E{�>2��=\eJ���h;��]=�Vw�* v��_��mmL����&2<�R�<z��=��=Y1�Gƃ<g��=R��=��>O �=XA?׭?��>���>= �=C���B��L��(���"��6�r>|Sq>�U�>cM)?�+>?(o�>efD�������&:ź�>��Q>��=�䣁����pvD>��>M�?��G?��X=��@���=�^a����=ç?��5?4[�>��2�[�b�0��f˿��`�R����|4����>���<�N]���O>+����g����a��=FN�>��\>;�b=4�#>���=�~��+4�>���>��>�ۅ=��.��1�=������)=StZ={��=ɪ����	��PW�-���j&���%�E�1�tk��yD�=�)?8�?Z���h�>����}z��)4���?"L:?تK?��]?YI�>y�NX��V���7��B��>i�?�K�>��_+�>w�:��&���>t��>�E��H�<?�?�����
+?w�9?e��>�&�庉�J�w��R�� ?���,�,�?8`�?/[8��ʾs����{�S���=-˾�IV��ӳ�9��-�/�Cr����YL��]�>W�-?¸�?
��/os>�0�����*|� ����t����>s�=�@>^��J�¾j����	��@ݽ%�=�>�>-g�M�<?w�+?a��>�ه?���>���=>>�(?��½�?r??y�?�Ĳ=8��=�i��꛺=ɂJ>��E�$�Z��5込��]"5=���<kT>'O�>�<�����=a[$<�B6=����r㜽����A0@=��h�}��=��=:;>��?)�>C��Ȏ=�N���\��>�k2��64�:,y�u����m�;
�<N6�> ?�9�>G{�=�����<Ǿ�N�3�>Ω?I�o?x�@?.���&vᾐ��Nb=U?T=�s�=S1s������J!�ɿ��j�K=��B>����&%v>�F�?�?P&v>�>�nO��ȕ���޽ߤe=���0��>��?���>Ma����/��Z��&茿}+�:¯�z~ľK>[�>a#>�B�>��=�����׼�t��ąn���Yʽ���>a��>WF?���>V%�=���&��?#V?ף�E��K��˰�h=�g?%�>\y��(�:?��!=<s��S���.�#��F�>�J�?��?��6?������	=$G��&޽'�ռ�W;�.}=d-]>�K_>�q�>W�)>���>}�о�
�=]A�>B�A=wΈ�G��� ү����Ì��4QP��������+���L1���[��!%1�wE�Eg����ľ��?���6����!ѽHbC�=k��䝩�9���Ri�?��?i:�>��j>��X�<�&����a]&��H۾�Ŏ�y����ս�_��T�侥��t.��U@�Z�K�ľί>�ł��w�������?#���<��{>�
1?��ᾃ��Z�%��B�\fS>b!>❶�1ʀ�C@���X�H&m?�-?M�����9�=��>u��>�O#>����|M��5U>21>?@G?�?y�-��I���͏ϽPB�?d��?9�H?�M��T-F��a�HOy����>N ?���>I譾�[ݾ����FѤ>�fZ?_!?W~��Ja��:�u>,�?�Zh��k�>���>�O�>ا7�km��b�sSþ��9����<R�=��=���WH���k ��x>�|P=�½Z����>�Cƾ������y@�X㷾��=�3�>����>�?�[I=�#G�r,���sd�0�oX?y.�?f�A?�8l?\��db@��ʾ�h�=�(?�m?�p�>���2��>CR�>,��,qg�,'߾�L?���?�v�?`�G?u<�p
տ.�������|����u>�[�=@�8>{���`��=#�%>�`��K����s�=&B�>��S>��+>U�!>��_>-�'>����*�j���|���@SS��6@��F��+���۾�qֽ����+�m�̾����Ӯ�!��z��͟I�6�=������=�%?���>9I?��4==>f5��>�!�0��ń��� �N�����փ��4���Q���:��� ��G�`�V��>�]<xG�P�?��ڽKɖ<Dڈ>��<Y�>ǸW>�w.=���=�T+>�a>$X�> �>���=y��>�?��d���ɐ��,H�2p��@>�""?��Ⱦ�3����H�| ���z�#+?�9*?1�>�`���R��P�'�(��>������Q����n��d�>���>ȭ>��=�d��O���K=��>}��>���=R��&Ӿ}�D�s9*>�g�> ����~�=�l�>�?�Ȃ?��9?�>���>��X>�B�>��T=���=B7>�>�9 ?yYE?�H&?9��>M�=9�g�:*=Ӛ6=��I�����.JϽ4�����Mh,=z�1��=N.T=��E��P���ڼ�P�;�M�=�8=v{?9[#?e��>1?�`>�8�he�h>��a0=�=����k>\��>�?��)?�0?�,�>1�	���߾՛�<�(�>�0�>�8���6������>g��>R�?�-l?p[>��>O�K�V�˽U�>�?��D??��>���=(9����nؿ ݃��M����M萾�&���_h>b}�>*c����&�#Z>�>y�_=�5�:>	^>7W�>��R���>�^E>vH�=&(�=�8�(��#�����<���<^k�=vW�=96�<7�W=����8��r���;�<h����B�f?�4?�}<�^z>-1���h��-=�+?ykB?��?<r?�P�>�.���uv�.π�P�Y��9�>��?��	?����"O>�tA���� �>ƈK>wR���������q ��c�5��?Y�%?uS�>;�@�ꅿ
�t�\�7��:�>F!����|�?��j?u��E}o���2�W�`��l��a�ZP��	j�����O��DP0�����t�j��>}y?�ݏ?�vR�SY>A�Ⱦ����b�X��Z���i�@+>k��>��w>�a�RYm���ʾU���{z�p��=W_�>
RQ=�o�>�h?ٓ?�k?1�?���>�v��&?~��=�x�>�u�>�=?P��>c�>L�F>�1>#�9(h۽cn�wL��&6�;l~�<�>!�>�~#>����<�O/=��;=���
�����;�=���=��=���=m: >�?��?;�Y<��=�:�V=�l�=�x�=����m���7��������/<&;�>&� ?�?�#�=������A�X0>8�?(�@?�j)?��Ǿ�ּ�[����Ѿ����=P⠽�wվ�H�w����w���=��>�쿽A�i>�?e�?5�>��=X�$耿��N� o>��<�L�>>?�.�>����v>������t� ���?�&>��*`$>,�y>�+>Ÿ�>�=؈λbE��8J���(��Ud��W�:�f> �>�)?߼�>Hƌ=g���ݿ���E?�v��Ս�t-���b��kI>��?��L>���4?�v��/p�H訿��"���?:��?�?��G?8�8��.��f�Wǅ=�������^b�Փ=(.����>��r;ޒ��-������=D/�>�@n>h��yE��O���<�8����C���ν{��嶬����i/�̕� ���w�=�K������

D��DK��3��q�۫���'�� ���ʜ�?���?[�>G<�>��;�l����?�4��;�
"ž}	��k�yh��߾	�ھ���y�;��i�2����>W�Z�9��QO}��)������@>��.?�-ǾR������^=k�&>&%�<
��B[��(e��	����W?w�9?�=�1���2��:�>X�?�R�>��%>L��O�<n�>��4?�=.?�^���9(��tP���?���?�|=?!�����>�U�,�����BT?(�?��>"���.���ņ��^�>��T?z?ӫ����i�{��&��>ͭf?7�X�!�>�r�>��>�
ӽ�O��؀�C2��w��;Q�=��&<wg�=6�!��-x���{<�>���=�s#��޾�ԣ>7�����Ї���,��a����=�:�>[����>I�G���<M�1��	���^w���\�;p@?���?Q�J?��_?�y%�PT.�������<�_�>���>\a0>r���&�>K�2>^����a�{I��iK?��?Fp�?E:R?&�~��ѿ|�����ھ�DʾoU4>�8>�D>p��9��=�)�=��=���=��>ŷ�>`�H>�Kq>V�>��*>��4>3�����)��u��Ƙ���M�������, p�P%��dN��� �c?������ܽ����l"�#
�՞���F=Y(:��#@>�T?�T??4�>�4�=��=�ʾv�����0H�����C�ʾ�Kf��♾����8ز�ȽؾxY��P�1=_}����?�;>�i�:�?D����E=�>��=~�=Y�>��<�X&=�x>���>[S�>-H�>Ѣ>�{�>� �ۄ���2v�Z�+��kp�~C�=�;?91������9�1�5/�����>��?�0�>���١����H�b��>?r���@�N}��%�����>�ܵ>{�=�*i=�������x����Ԗ>O;�>��=�W���ϾR�*>���> "龞p0={9>>�3?�5�?tA??���=���>�|?>ԸG>����yg>�J�>�ѫ>:�?�-?H?��?W	�=�a�$�.=�4
=��V��Ĵ���g��a���#���C�e,����=�?>��T=�"�;̱����½'�7=F>=m?r�?͐�>Vg?��[>&f���%i������ˋ=�`p���p>�>��>�%�>1Y?M��>�!�<���������3�>��=�#m�Ǿ|�jV��x��=��	?7ׄ?o`U?i;�>�0>z���y2�=�*�<g�>l�;?���>y��>t;�%��ɿ�o��K����<1#�=@
j�w���$↾S|ȽռB=�5>�a>j�P>:|'>�Ѧ=�`>T��>�J>PA�>l�y>>Λ<TS��� =z0��G�<���;,��x��t�|����%�)i��T��+��Ǔ��)��l?J�?�@6���8>r���/�� ����'? �T?�.?��`?�Y�>����~��ą����Z.�>9}?�5?���/5�>M��M=�/�>g�>���������<2W��ƊF�Yc/?]�-?�u�>bV�����k�pZ@�i�>�j�4��<��?�6^?/g��ZϾM�!��@�(��>w����l]H��휾�����8�
��g��2���Ih>nZ
?к�?��ӽ�W>!���s��!�c�i#�� �=_�">ܳ�>,�E>�M{�^��:�cϾ��T��v<�[�>�܅=�5�>�Y?ix?}�d?�?'�?l�(�?�s�=U
�>��>Dt?"?-a�>Px>��n>���<s&]��������a}<5��x�=e� >�*>�Ɵ<�'3=?:=[��<)R�λ�S��<c	4< ��<di�=�T�=��>]p	?[��>ߛO���='q=)9�X�n�Yx2���V����y����(��6>�Q?��?M��>JYj<�/��1�	�M���}>�-?
N?#h8?ʧ"�����\X�x�پ�;�n��=���=*־6ݾ����+�-1>9��=����>�ٟ?�7�>���>OY>q0��Ł�\��4a>,b����>S�$?���>Wߔ��>��Վ����mA��V^�y<��n�&>&�j>|�)�u�>��x�C>"=��&=�Z���ni���Ž��*�Nt>���>��?�rQ>GW��敾��3�̯??ȄȾ]Y��5���.�$�<��&?���>ׅ�=��I?:���pȆ�'�����;��U?���?k�?�oV?
t��{���W臽�K�<� J<�����Q=�M�=�gj�>�7>�좽�R+>���g����t>al�=!�ź�ψ�_靾��=Lֿ�>D)�ݠ���t��u�о�MԾ�I�ĉ���+�+tȾMP�o8����lY���z�;����k��1C���k�?c��?Vw�>⩁>�O-��J?��ʾc�=�ľ��+��u��}|?�@����˾���6� �6�:o5����� �>=�Z�� ��;�|��(�ed���A>.�.?��žj���7��L�_=>:'>cy�<(��m_���s����^yW?�n9?�뾳A���߽��>N
?���>E #>	ߔ��7� ��>��4?C.?\#�����8��g��wP�?o��?t�>?�����:��
��g�D�"?�?2��>q*u�|3ؾ�񄾌��>��R?�?����/�k����v�>X�X?��|��_>�G�>Ӏ�>|��dh��Z,����;Q�V��=^d^<Q@�=�g����f��
P9�.5>>��t������>��Zƾ�����K��� ��rμ�>���r�?_l��A;�a'��*��ͭu��b,�3?9ޙ?�<?JsY?�����M�L�Ծ��=AI�>9*�>S6{>�闽(f�>�A�>-��ᰁ��}��%J?��?V��?�6M?v�l�}a迥;��G&�L¾��>��K>���>bo-�?��=�d=
�&�o�<�2o>[�>�>>Y
>�;,>�>�4=���4"�J����h����M���!�B0���y����l�@�t�������?���Ž�4�w����"���>�H��(�y��M�=��"?�r�>���>���=�^4>y<�������̾�A¾�� ��r;����������A��������	�E���>!����>�=O�{=(�!?�\��]��<;��>�L>�p�>#��=�>-w�=V�=�N>��>"ӫ>{>rg�>��܋��[����C�-���=*?dϗ�Rch�~�"��K*�~ƾ�2?bY-?환>�������v�Z��a�>J�|��2�X-ͽ�1)�g�=��>��<�9=Nu��t��THɼj�>��k>��'= i<�A�9���n��=���>�T���<[�_>;\�>�V?�K?1_>���>*l>'��>�H�<�+`=��<�c>�A!?%�4?��F?R��>Qm�=����c�=��<�R�7�T��%�������>R>�>"�m=���=;9彡5.�%�=H���=��;��>U�?��>�^>Z>�𵾮ڌ�a��$}�������u>�>}�?1K"?�2?�J�>2�Z��-ؾ�;��>7�y>G��3y��M��0�=^��>�x?.>7?�h�=��<��,�+�-��{*>�P ?�#=?�>� =p���v	��7ӿs#��6#��Z�C¢��x�:<DG�fP�v�C��7&�A�ɽ !F=@kU>0�>��[>Q�.>:>��E>���>�Vj>j��=;�=3/�c;�no�a�@=F�Q���;_}��������򴲽�'���v�4\���9@�?_ȼ X?�m?n�5��2>�}��E�Ⱦ�)~��?Q>M?N=!?�{\?:��>+c'�m�X���w�N𡾨��>M��?i_�>�!�3�i>:ż�q����>���>�
�:�ߙ���=�o�����Ә?Q;?���>5$��v���[�� ��?	������`<�??�u?Y��� P;�N�[��������"�\G;��5��%2��^���%�����:f>R?s9�?�����W>k;ؾ�]w�D��>{#��}�>�}>�(T= �7�D���H����H���>�h�>L*�=���>�M?W1?��u?\R�>
w�>TZW���>6Nt�64�>���>���>�m�>:��>��E>� �>���=9��+	�5���`��;�N<NVK=>�V(>L�z�2�Z�v�=�=`l�e`��	�����z�<�=�jP>\�>'�?��?���ϽB{_=@}�����=�4>6.>.~?��d��h�{=V=��?��*?�
?��=�,�����e����>"�?'�H?��?�A.�e<J��}ƞ�X'�W%	��ɛ>)�w������G���	>�H�>q��Vr>d�?�0?C(?�h�i�*�Z�g�H�^�=��}���>.�>Tt4>l,��܊8�<1|�?4g��/�j�=.]��i=�B�=���=�9>�l�=4��=�)=�J���4��� ��n��>1��>>p�>'<>�S6�($��+��f�B?�޾_�,��� �����(�=��>}b>�2|��<?���F偿&ή��'��
??�l�?@�"?f�6�_6�3�>Sb>1��<�6�=�� >�ƻ�;����=�Go��i =E���褼��"?!�>�V<�=���)�BԢ�̿��D��
��
���`X��Gɏ�%�ϾC�H�>#��U�A��Y�������|����?��z4�Q���"�Ծ8����~�?���?5��>�A>FF�7Q8�!q�T�!=�LҾev�����kk�y��v-��W�	Y��4�e%�j׾�ś>��Y��@��|�|�3�(�ӥ����?>�0/?�bƾUʹ�����g=�e%>��<^#ﾞ���{���"��]W?��9?�?�}��F���>��?(i�> �%>����U�4�>�A4?��-?�)�A��f6��C$l�?v��?��:?����@�Xd���Y��b#�>�1�> �?��½�Jؾ�M���.?�WV?�l�>ï��}����0���>�Go?�NX�C1|>��>s�X>":Ľ�D���!���V���ý$��=���*�	��2���
�>��=�t�>&�>6�k��lþ>#�>rȟ��V�"�޾�:E��Vؾ��>��>Ui����>{	�&�=�)=�����)x�����]L?(��?!,I?a,j?5n!�{"N�:��J\;>���>xy�>��t>{[���t=ť�>����]�k~۾�B;?�g�?ڎ�?��U?�l}�ݿe?��c�	����� J =P�>���=66�i�8>8n�<�1?=���<�\]>l��>�QM>&�6>^Y^>W�0>�+�=����g�%�R��WP����J�9s��h��I�E�U���[V�����t�ϾY?�����N¥���h��.�p�m�=�`X��>
�=?#8�>6?��>�c$>iY���u�G�ξH�оՅ�N��_�(h}�=-�������޾|�4^��T+��?��>q�> OG?%4��W�;?l�>��=�˱>\�M>�aS>�VD>�-->��>�G>CI�>�$�>@��>��<�}��Ɖy�K�A��*"�c;�=��)?�n��O�����/�m����H�>��!?,	�>�;
��ޒ�u"h��)�>�[���U����866����=J)�>M��=~��<n-P�Ső��L �e�W>�zv>���=���ʖ����ｐ�;=j��>��ʾ�^�=Jh>k�?�Ik?voL?k&> c�>�>g�>��<��>�K�=J\>YG?Oc8?��F?��>I�=aW��9�	�P.=of����h����N;�p�=��<�X>�xv<��7=�s?��^M���=9Zm��I�=��=���>?V�>��>��=�ዾY�e��}Ѿ��<��}��>�F�>A?�-"?��?t-�>N����lV�JQb���>���=Ogk���y�$ߪ�:�Z��x?�	p?��L?��|>a�=3 Z�Hn���#=>�>:�<?>�>�R=������	�޿I�V�+�_�vǬ����>�ӽ����>7>H�H<�p��R���>��>�ql>�i�=,u�=���=��V>�P�>�N>�=^�={8�=��$�9J�<�c4=��-�n�@<����<W��jV�	ٴ��I�'���U���@�=֜?b?A`޽���=��O������..?�g@??�fj?�ۻ>T0a��Hq�3�}��镾���>
��?X�>/E"��`�>��̽�z�:���>�B!>�����`��0Yt�婓��˔�L@1?��7?,��>�hn�υ���e��;�kl�>����-)��?�-?��g�}�d�'�0�b�<��\�>�yY�.{	��ڋ��O��d2��>�'� �J�l��d�>E#?��?	�^��>t��<5��]�Z�,��tV=*U�>�>�V>���� n�H�y:h��;��	
>��>k�=q��>�?]bD?W�u?h�
?��>�z�	��>��ʼ %�>2��>!��>���>��>ë�>d��>aѢ=��K�Cy���u�6m
�ef`���?=�D>,�D>������=¹�;�l<0�H<�ې�X��9#����c���1>YQ�>��=�L	?g��>�W�w�p��<��*���IǼTW=��n�m�����⾣������;ɸ?�9?��?��=XH��E��5�c�b>��+?��A?�)?� ��9HA�����C�A�����J<9S�>��+�u
 �8+�Q���o>s4<>sd��?u>﹛?�?OH�>a8�=��+��`i�����.>ޥ
����>p�+?}��>`]��UDO��5������\)#��L=���f>wA>a<=ҕ> ��;���wֽ�2��=� ��]����6���->��>�(?u� >��e�ш�����aE?@ջ����_ɾέ�%�=1�?ƻ&>@r��a�?Z���D��Op������?�T�?��?J�;?>AF��nؽ:��<�� >�U�=�O���*�ȓ��趽���>Z�$=��(�f��DA3=.�?��>�D>*���m���ռ�����)7��۽�������Ծ6L۾\�������t۽�䠾��on��%-�\���s��%R��0G����+�MZ�?,/�?5�>;j>fxC�_,��Gľ.��; ��i��R:���É��W���O��
���@��?� ��>	��4ƛ>��Y�]@���|���(�X鏼��?>//?[fƾvִ����F�f=k^%>���<� �w���z���:%�G\W?��9?4G쾲 ��,ὄ�>��?Y�>K�%>�%�����g�>6A4?S�-? �켋��h9��(ܔ�1j�?���?ux=?<��U
>����������>�?Mp�>XG�An̾����;?H�D?ɢ�>���-6��ʛ#�w��>Z&]?�&j��z�>.`�>F"�>-���-@��+�}�����K��h�>�r
�0��^�Q����8��=!��>�W>�L^�Tr�����>��~�N�$�H�P�������<��?e=�/C>��h>��>n�(�p
��d��������L?莱?�S?�a8?XR�������=lͦ>+��>��=���U��>���>&��cr�c/�ć?�G�?���?�dZ?�m���ڿ�I����%I쾬=ϵ(>�>�>�� �χ�==k=�l|��ē�-!l=���>-��>��>���>p�8>7uj>�G��\9(����6�����H���U����L�W�̾��S��'~���ꩾ��ƞ���q�;�<�¤��\��2|(�3z\<[�&?D�> ��=2�=�>�$����;�>��{����W��d���g���E�������g���t̾�
�PM%��5
?�ܽj9?�i�>��E=���>�S]>�
>�@?
?��c>"p�>J�l>���>��>���>�r�>s��>4�<#薿��f��K��$�A���>���?L6������ ��}�g�9��<��y=]�>��>�x)��ڞ�z����r�>����nG��>�<��$g����>��>\A_=<��=w��<)�򾶡�}�ݽ�"�>�!>*�>��Q���>�=k��>�MH����>�[>��4?�PU?}�B?#�ѽ��>�D>�w�>8Bg>����l�=z9=���>i�U?��A?�?��=l0������a=��A:���2<�X�����<��
�i����=�*�=6s>P�<������<����Y����}>Ѕ?l<L?V�=��?�^5=����X�u�=�9V>�k���@?���>L�>��>?���>0�A�z���G��@�ͽv��>7P>��(��Ww�r�y�� �>���=��>��\?��>$����v%�*���>Y}�>��?&��>��A�J�>����⿴\M���^�:O��0fO>�%Y>7Kr�8!ս!�=;u=F���*�S>Y�>��#?���>��>&�q>��>�1>6B�=3�<F��<�>�O�Cj�=�4=��8����k<�(��8N>i� �B�m�����j&=H l��?��?�&(�y5/��0���ھ������>�>jc�>��>tL�=�	�xzL�iH,������ ?#�i?��?W]D����<����'�<�S�>��>سN>�H��y(���
���9�=u�>��"?ʽ>Dcc��;Z���g��!��إ�>b�G������?�$_?���WY���U���w"8��P�<�����:s�D�½��6�&�D�g���<ñ���Y�1^?n��?b����<�=D��f��ᶃ�D�h�_=�7V>�`�>���<_p���3����I����F_T��8��֐>���=�:�>"U ?�A?Q�m?�I'?:�%?����;�>#�<ӻ�>�>�ݴ>?��>Nq>��$��l�>��>mKs=���ׂ�2q�<\$m��J�=��]>��W>�-�=���=��=�@������>yѽ�˓����<�L=��>���=D*�=��?�c0?h�g�Ќ��U�Cr&���ٽ`m>���><�=�ɉ�G-������
?`�6?���>�t�;y�ξ:�S�6^־ M=Z�?��7?K��>] <Rr>C�վ��V�J>I��>��4=��Ͼ�h�3Ak��o#���>Ġ�>r�<��G�>d�g?�?�u?��=g�9�Sw����W������h=�S5>�0?b��>��6�e�3��0d�`-[���,���>='<4����=t��;�/>�O�>��=}>��=dL��t�_���>��Y=��>ݼ�>�??�:W>q����d�׾[G?'����%��餾زd�����נ�J�>Az�>'�>�r=�R�}��p�>���)?X��?P��?7��?t;��C���*=Hh>��>���=腱�g>Py��p~���<�ؕ=�u���ט=e��=Fj\>G����u�LM��X
F�YU����k��M�=Ρ��;������<r����=����0.�-X���;����W>�Yᾄ�k�WQ�����a���Ͼ Z�?��?l�>j�s>�1����{��v�=.갾��]�̲ܾ�釾'��a���)ξ�@��P4�sC���E�)H�>4�X� ���"�{��@*����߲?>�g/?��Ǿ�������V	S=	D'>X7�<��ﾥ̋�y��N��%U?�t:?c�뾥y��~M��>�S?���>�(>N��oo罪��>W�3?̏,?3�μ����3ʋ�Ά����?pS�?��<?9�B���;�y�8��&?�
?�!�>�˄��pվ0��x?e�2?�G�>��0���v�OI�>��Z?��S���[>:��>��>�@������ż���[}���s'>�-<! 
�X��m�5��3�=�ǎ>�kv>�'9�����1��>cP龺kN�"H�݅������<��?co�%�>�*g>� >�)�Ě��������m�M?d��?�xS?��7?���G~��ᬽ7M�=QЦ>�9�>���=����$�>���>�w�/Eq�����?��?��?>Z?�(m�Կ�A���������)>��>�dQ>�MܽM�=��<Т�< $ۼ"�=w}>Wq>�S�>�Q>̂r>��_>������+��Ơ�@㐿�f>�U���8���_�i��:��C���lƾd�žF�ֽǵ��t�̽G�u�p�{��ս���@�<,��>�O"?N�4>w��=� i>������=`��I�X���xa�2Z��i��L�4��Uy���G���!�}o��?�u��y�>@�"?>���>��>��O=�ր>$�.>��+>�(�>Qʭ>_�>
��>�>��1��a?9�0>�ا��M��|����s���/>�V7?�}$��?<��h���5�����ɵ>>��<��>�r �2~v��+u�+�>ȷ�-m������x��>N*�>q��;�=ĭ��߾mۿ��`��ͥy�
�=p;��$¾�p�/6>�'a>z
��qa�=4����"?zW|?�V?�L�=�u.?��Į=Y>>�C��)���o�>r:�>�AL?zM?"JE?q�y�N
��}r���
�co�S������US~�{���i��=��=5H>��#> ��q�><�$>J�=�� =�#�>��M?�L�>ڝ�>Y��c�{�)�[���� {/=�Ƚ��?+X?'K?��>F��>��s>�>?
��iᾯC�>�e\>�92��D�L?I��0�>TY>S�)?�=H?�ʆ���؋�>�=�R|�W>Am?t��>CW�=�nf������޿de"��'���M�X�<�I�<w�v�O�����=����ߥ5�Gv��z�eX�=M�>}Vh>!�^>��{>���>%> ��=�l�=�C�X;��1�]>K
���a<�s�<��	�B� =��mO�b�e=6O<�Y�c��@�?�g?6}���Q��8�˾Uat��:�>��>�	�>.��>�=�;�U(V�	�-�m�I�P7?�q?�>\]����<�i��!�<n�>���>���=�ڵ�#+�������߼㟞>��>&��>"� ���a� u������>��<٫G��?�7d?�_��¾�.�|��l�6�Er�=�7������a ����h�&��\�j(�^��G�"�5Ӊ>�?�?\����W>����e�������	������<��>��>$ <L˾.�&�j~־��y�z�M���>؄=��= ��>1/�>�bM?-�%?�U?G�Ծ'�?�>�4�>N�>���>��>p�>Q��<��b>��>��>3���ĒA���ռН����/<{�=D��=dy����<�r>I�3>h��9�4�c�=�+2>��<WW�=b/�=(��=ժ?<�>?��>�JI��2ռ����R�����>��>U���%���h<8>	κ>.T?`}�>��=u'��~ţ�ֱ��N�н-��>8.j?�
?Bq+<+զ>KZ������pn��#�>�����*ʾ�;�`e��V�>b:?��>�>l�k?y9?��?ru	>��"�<����;�:"Q�G��D��>���>f��>Ԫ׽*5�s!��?�J�_���-�*��)!>��=�ڛ;zn�=U=��%>Hq�����;9�<B@�=HO�����>�>?��>��c>�A*>����bB���+F?�✾��>����žQr�H0>ō>>��ؽ���>��	���s��Ȥ��;=�w�>��?}��?��g?�S7����H>`4K>��>p��<.�D�=1b��g���a3>�=�bz��������DKG>�)u>���f�վ��ᾲZQ�Q9տ�|�d'�>�eҽ�|5�a'D����AGм^���}ֽ�^�y+�����<����|F����"繾Ě=�$��ɤ?N��?$B>���=��;��X!�����/��=��󾍨*�v�������1�=�
%>x!����L�2������(�do�>f-f��D��qr��=�a�]�{I>@�$?�ϾW����#��Y���
>�/=�n���C������j�.��@?��7?��Ᾰ�������8�=Ic?F��>r�	>�a��c���m�r>#+?<%?H|�X���{N���&��S�?�ݿ?'y??�S�Y�D�ܷ�+61��?/�?�p�>!u��8žZ����?�65?0��>^u�ݔ���r�>��>��U?+W��cb>�E�>E��>�^�8��t.g��Ԝ�m��jU1>��lW���^�� P����=�Ǖ>�	s>]�i��M��2��>�9��N�ʡH������=܏<��?���a>�#i>�1>�(����̉�NH�9�L?1��?[�S?�f8?{Z�����������=%��>|ج>o��=���U�>���>�h�sr���t�?�F�?9��?�SZ?��m��Fӿ�
������A��"��=B'�=z�>>��޽˭=_�K=�ј�"U=���>R��>o>,<x>a�T>q�<>%�.>C���V�#�ʤ�#ْ��[B�� �&���vg��{	��y�J��Oȴ�f�͘������Pϓ���G�g���R>�J�<�wٍ=�?��?z'�<ɞ��o��>��^��Rʾm���}	�"1�r(�L�ϼ�z�F�־�V��dw���߾�����&�Ԩ?���<屘>(��>���=��s> �>��>l��=��O>��>]��>�lm=�?�>G��>Wd�>��9>��?o��>6������J
n�a�?=�{A>F{P?�#W�-n�_���1�l���L4v=a	�>��>��V�㠉� �p���>+"�>�վ�=캸I,�c	>�_�>e$p>�8'>���;8��2�
���;�=ء>fl�oٕ��3����|�\�>���sYk>̦ιF'5?_f�?5?��<7�>X;�<bӎ>�{�>�$�|Ƈ>#��>*�y>z:?Q?�K?��1�ΉU��+`��������˶<r���.�<� 0��3Ľ��>�5*=�B�<dƽ�ϼ�~���M���L�=�A����
?�CC?k��=]�>�z�U�q�_�P������B�=<���k?	�)?�j?�F�>��
�t�>}��=#bƾ��ľA��>�P�>e7�yƊ�)~��K��>��.=�
	?��]?�u�������nR>��>$��=�@?��8?B0>���A� ��ƙ�5O��W+�P	[<�d=?���/�䨣=QU=N�罣.���8O>A[)>3�2>���>�>o>1>�~�>���=�O%>X>>�B=<k>�$��g3>���;o0�>e,u=�� �y*�<}��Ԩ�@�1�';<��=m�E���?��(?7��	60�	mp��߾�n��恋>�>I�>�?���=<��Lu>�&�<�R2ӽ�3�>-C?ޜ�>	p@�Q�>���G=�M��>Aa�>w>Je����W�� y��[��3S>#��>�#�>4KϽ�X�RM��OZ��>G�=Rs���?d6q?:��J���u%/�G�ƾ}Y)��,�;�_�=u׼�����j��(C�|���=������,>:��>�н?1D��=H�i��ԓ��N����4�d�=��̾���>nŴ>'9��s�SfT��K1� W����0�TG�>���<�E~>]��><D�>��N?E?پ?�j���/?J7G>V>�>u)�>��>�_�>��>r�>*�#? ��>��>�����SӾ.d�T�ݼ2*>3d�=�,�=ֈU=@�=� =D�=��>$��;��=E�=�A��!�=c�">���>؍?0^ ?����n�=$`b��������=��¼J�����}��i�t�<B9e>��&?�߼=�D������� �)��<��?Wa?���>��\�
�N>\��Bm�W�P��>즈���t�����þC���>~��>ݰU="�s>;"|?y�?��>� ���k<�l��J8��=�~�j�>hh)?���>{U��j�Z�	���R�rjI�Y�3;��w��ԯ=&�=-�=J�=�@*<C��=�V�ZR7<c�=�i=nV=�c�>uO?�3)?,�>vAe>�J��Cu���I?����:���桾��оY����>2};>�B�ge?H(�]t}��ۥ��=��>r�?���?��c?�JC����.]>ۙU>�>�V7<�(<�S��⌅���2>�F�=1�z������7;J\>h�y>�̽��˾����H��ɿH�N�[�>Aܼ���n�\�j�kv�G�G=C����>�x�|������>%R ���;R�������)Tw�������?@+�?��U>���=_`u�i�-��p�O��=֗��`�����m�8���S��h�]���ǹ���X.�he�:����>��X������|���(�U���� @>U/?}�ž�������0c=��#>�q�<)c��墚����B�V?Y9?%!��	���Oܽ�.>`S?[Q�>F]'>T���.��ґ>�4?�g-?�t޼��M���ƍ�qP�?{��?��;?U�A���B��C	��'�b?��
?L)�>h z��X־?���r�?~,*?٨>����v�����i�>sJ_?�eJ�I�Y>��>�N�>p��\���-/���������� 7>�e�;�:�<*b�/�8�@�=���>�\>_�]�4���6�>~��OO��H�w��P��ֵ�<'x?0��>�i>��>"�(�n���ˉ����^M?-��?��S?Zb8?-��A��L���k��=��>�>���=�N�ۀ�>ק�>�l辗Kr����r?"8�?ų�?�`Z?�dm�s׿]����վ6�پ��n=�֔=EA�>&�G�9=jr�=��<�qv����=��@>�E>ɩ>q>�>��z>A��>Kj��iN)��h���0���oH����Ӗ�����7�ԾE�׽�
� b������2�$�:��*�w�l�%�����E�<�k=)�?�*?��>KJ/>�W->�6ѾT9�)�[{��r�����2ž�rQ�G�����]��׽ҒŽ?�6�Q۾�D�>�C��t��>���>x���sY>%H>�>Xm.>�1>��	=������Y>��:>
�P>�?��>q�>�NB>��v�a:��[k`��Qf>?��>T�d?���<7���C�d�|~1�GS��>��.>/�[>j�����I��Mb�B��>�f�����������r�A��>��>��>(=+w��|h�IX����>ϐ�=`�C>Y@L=Ot��(�
��>��ﾺ\�>U5�>�,-?!8n?7a?��r>~�>��>iR>6F�=:@>���>��>��>�?��?0��>F�=Z6�C=�=�c9=;�1�cm�9
�l�=M�
;"2��,�;�_e��b<�����9>�#>ܯ��*\/�m%K����>W�=?��>^Ͱ>@�J= mQ��-��Ԡ����>=繽˔�>��-?�6?���>��.��<�>r}���Y�[L��ۂ�>N�x>HV+�K�R�����>�{�=\8?	7+?����9�����<2$>-,>��C>}�
?�?i�<k�ǽ�#���aap�%_�RO��¸�Q7�>��:���%>;��>#8M�4c/��䇽�@>Y�>�|@X>z?�a�>%��>���>��=�"�<�_>a#�<�>/}�=��>@E�������Ҙ�2�_��������������=��=�;>(N���?� ?�*ҽ�?��
彣�¾�g�F^>3?���=�m?���>�?3��qX����U�7X�>��S?��-?ݚ-��U<=�W��%����>��>p�=$S��;A�+�d���>���>�A�>���>�}�d%�*�7���ھ9u�>7�]=�>��G�?~VW?B����̛�ʕ���&��g'�iT=���=����Ɨ�����̾�?��P�&�GM��c�=e3�>m�?И���=������˴���߾�6�>�/� j�>_��>9��;�m�O3�^�a�����{ܻ>3��=%�>h�.?ؼ?�\?��?�?���%j�>N�h>I��>�S�>��>�?��
?��7>��8>P��<<K��>p � �|��~�==�p�г�=#I_>�*>��>�(�<-o=-/=C������I�+=_��=S9����=� �=�u�=1l?Z�?��:=���=}��y뉾|��:��Y>�?�=���nec��E���p�=^��>��?�ɶ>j��a�����)��C��<9c�>[W?ǭ>��>��%�=;7:���ܾ��?�칷>Z��<�ž���#(�q��W���s�~=]�}>	�p>E�k?��<?c,?M ���-���Z���.��y� �K���>f��>
UK<\������7l���\�b7�ʺ��,O� �	��=ME�=�ی>�>R
>�ʼE���<������CQ�<T�>sܠ>���>�n>�T=�W����H}I?8��� ��F��!׾i5�� >�EQ>�%���m?�?���O2��P:�E��>D$�?���?�o`?��C�H��"^>�_^>��">C	�;`�M�LZ+�v����P5>B��=
xt�6z�����;h�^>�E}>��ƽ.Ⱦ!��!�:������Q�2
=�����h?��_$��t��ԣ����׻:�����ka=�㡾)��l3h���2��#�<�t����?��?G��>�0q��T(�����a_þ�Ϊ=<��۽ֽ�0���\K�:s�=B�<��9+�/�	���e�͎F������>��X�����|���(�뒼��?>�$/?{Qƾ�����z���c=�l%>��<Қ�ȧ�����Ũ
�\W?3�9?=M�@�����ը>_�?���>�%>妓��i뽬��>��3?�`-?�H߼:县(���	���>�?���?�A?w��!/?���-�`�!<�e?�Q�>��>���4�������>���>!I�>��̾V9���2��6��>S0??�AU�=��=�Ȼ>l�l>ʂ���d���P
=�M��T���%�=ə�<.W �}g���8��b(>���>�|A>�R��e����>;�Y�N��H����)�����<bm?���>
Ai>�>8�(�v ��U��������L?���?�dS?Qj8?�7���ѧ�5�=T�>�Ĭ>���=������>;=�>ML辗Ir�)��?~G�?
��?mWZ?c�m�xٿ����X@о˂����=,9���=��O���=*�=e9�=�U3<�}-=p�>A
�>��>�X�<6K#>%�>\���X+����R���'G������U�����'R����\���E�w�E�|�ga����	>��i��{��m���e�>
�?�?��C>��e>*��=�ڼ]7������*v���)��^㾻3��ˮ����(=�����d�:3���%�?�C�MVǻ(lo>f�==ͥ�>��>��|>և ?t�h>Lē>}���NM>���>�?v>�	�>O!>s�>
�d>�/���6��m�|�����"��!1?�e��p>~(h���?��A�#��>Ε >�`F>ܫ�"J>��4��>ޕ/��́�a��<�7��Q>�l>>[ڀ>�Ms<R%���Ͼ]�.�������<>�If>����y�y�=J�l�:��>�=̾�%=K�="�c?E�|?�~m?�	�<��>!9�=�T�>�e�>�)���ݽ[��>�
?޶�>}Ce?}�K?�4=|<�5-���C=�I0���Th�I�%��8�=S 4=#,0��5�<L�<	�>���=T�>��ټ����d�>�L�>�u6?���>f8�>�8� hh��u[�q�ip\>�h]��L>�?��?�|�>���=��;Ț4�M���־�q�>�S>�1�$�r�Ӳ�=�>�>�l4>t�=?^N?#7���+㽞���~�<T�>���>�<?3�>T�>΂ >(����忻<H��98�>��
�=���=!�;1FL��7�<���<�a<��+;�ޙ=Ė�>5�>��>EfO�漏>��>�F�>� >��l=!��=bO>��<�T�<,W�o�A�x�h�;v�<�ډ�iK�;�YȽ�Y����>m,g��ʾ���?�o?�LF�hYA��KW���込���B�>�S�>U�>���>�k�=i���uM���1���E����>+c?���>rTE�ߙ=���+�K��%�>�-�>�>7	�����ћ���o)<�H�>!/
?��>�F����J�5i�x��̂�>¾<(�|�j�?�Fd?y���y׾hK�g^����u����=�[�o�Z��� ���׾<T��6q��5�K�-��/?N��?��W@Ƚ_��%`���H��ͧ���>��X>(�h>j�>�?Y=�ޮ=��M�޾N��)�)��Ҁ>��=�|K>=˨>�R�>�d?��?�g/?�V��?깲���>��>N�S>�E~>G�?u�l>䴞>��>[^L>�+�������Bc�Nw>wą>�J�>����!:���}���f��|�7��y�=s����>]�#>Q�c>U>��?��?�H���1>�[�!G��FӮ��K>
י=!�G>]�����>� >�7?�iA?�ѽ0-�] ��P�'�D��9d����9?}�m?��?KtQ��ӑ>������n�?�#��>��=ૌ������������2;�/�=x��=LO�>�Aw?w_G?H�%?ma���Q�a锿�*�;�Ct�� �>yk�>'Ŀ>�f�Ϥg�3&*�hq9�h���ڭ�NQ=I��=Ōc=DRC�->�=�>�qK<>.R�� ��T�4ܗ�)`�=�)>}P>���=���>D�����Ծ�I?����f�%����Ҿ��%��*>�eA>�:�q�?N���t~�����M<��v�>�+�?���?zd?��C��F��*]>�[W>��><�$<UA��o��G��,�4>�=�)x�OE����w;��]>R~>ʀ˽a˾"�?D��Ŀ;�a��v��o�����O�[�����������;#�G���پ=������y��=F���l��%���x�0u���?g��?f��>��t>Ʀ�/��EA�"N�=u��3�ѽ����	��Ԛݽ����l޾�ϰ��69���ľ���%�>B�U�^���m�z�p�)��Կ��A>�00?�Ⱦ
����^�H=r�>�ؘ<d��0���rq������gV?T :?�M꾌���
�㽗�>��
?���>��#>w����ʐ>�5?y/,?Z�꼫D��^΋�I��}��?��?�Q?W@>�3T��Y�$�X�q?�d�>�]>��<዇��#�����>L�>�?Ο!��sl��� �>�A??eC�z�?>�F�>�t8>M��f�+<�i��n���>#�2�����DM���^����=�{Y>�/i>�1N�!s�i�>�1辥45�J]�?����� ���=願>�����=�SB=ͧ��r�%�\;p�B��Lu���>?�n�?�O?Q�C?���p:4�@�[�!?��>2�>7,�>8���,�>Y�>f���m���ʾh�+?��?�j�?I�W?�N��Iտ��]���v�������	>u� >�(��I�>4��=ey'>m7�='�N>�q>�+>Y�_>Wq�=��B>�$>pR~�w�'��R������b�����Ͼnbv����\�1�����f���M���63��-���u�;�˽�Ґ=]�K�*�H>칸>'Y�>�A�>J��=���=�Ȁ�X���g������9��7��=ž�^���S�N�S��a���̈́��؜�_��Xx�>͂����,>t��>K濽�T
>��>��n�i�=�j>�X�>��>*�>��L>ǹs=Xq>��>�f�>4��a��	y�$�1��Z�2��= ;?�L#��ʾ�S�(��І����>�E ?T�>r�"�����&1J�O�>R��C�>��!*��mŽ�#�>��>�'�=]VҼ���6^����h��T}>���>!g>C�4��x��
��`�>�w�>��Ծ9c�=��z>i�&?�Gr? 1?=yx=���>��S>~��>��=|EI>�ZW>���>��?t�6?��-?t��>�ø=��P�<��<�(1=R9�йp�ժ�����Ok(��Yq<C9C��Z=�@K=�1j;�}N=�W-=?�ݼQ6�:���</��>�?�A�>���>f�n=�о�mB��~Ⱦ�d��X'g��p?�:�>���=�$�>]X?V>z�><��Q~����>3�&>=������Ǜ���a=ay?�&�?�D~?l�>S������y�>M�/>+�>��?�Z�>]2`>�%>#��9ݿ�����'��[��T3�<G�A=(�T�"�~=Ԃ�>l:��
�=��<�>�P>r�>���=r>�/�>��>&�T>F�>gɄ=G�(>�-(<�I2��G���^�=
t���V>~K����5��f�<k�X��=������<q??�&	?=%�=��=o�x�'lm�5v��c�>3H?�'?�$?�[�>�^���\�&�t����^�?pX�?IX�>��L����>�(j=�
>��>�I�>��:���b��B���K�Z�����>�iD?�"�>�5��J���y��X
^�l�>���<�ԽG;�?�Df?Q��i}����Bb8�ϕ
��R=c#���b��ˎ�."�IW2�$���.�����^Ei='�?�?�I���j�<*��܋��Nu�?���o�=gb�<&��>��>T6B�����[������z�4�G=;��>�vo��i�>eo?�7?��;?~1�>�;>�����u>|�`�%T�>���>��
?��>�v%>sA�=)~=�}�<�9r��n�@|����5�a��=��x=CKx>�U%�5�D��:�n�U=hH��q�`N=g6D=�.�=\�/>�f!>�1
>��?��>�R&���<>��>�0��u}�� �b �N�r<#��L���,�>w8P?8?Ue?	G�=���/�'�4-���_>���>V`9?3?��>@���U!��b̾J��=��>� нC�ܾ�G��"���	o���>h @>�����c�=m&�?�^#?/��>\�A=�w�U�c����i?>���>�`?�֣=h.�Q\��Ҕ���~��Ir�:F򾼙���W�=��M>a>���;+ǽZ�Z�T9�=[�$��$*��J�=[�*��p�>>��>�A�>���>���=���a��Q?)�޾;F�v�$o߾t����H$?[*?�7�=lR:?��<���v1���	A��
?��?0�?ʞ�?er�5�����=�ty�"�>��8=�RW�q=q�3>���>�,�tQz���>���=�2�=f�f> �#=U���KĽU,�<&����{��S>c6M��>� #A��`�����0.���E��Ԗ �>T1�x�ӻ���W�F���J��Ұ�8�q��R�?�J�?!��>J�z>4=M�2l���`�i>�e��4Pڽ�Ӿx=������VԾ� ��%�@y<��17�;-'�O�>&�x�E�i��
Z���/�>���yi>��?Wu��*?�"	H�Hs���>�!�=����Q���薝�Kj=�� S?P�B?����+)1��þ?-�>�cY?F��>�
�:���d8�s>��?k1?<�=D玿���/��<Ժ?��?)??K��[�g��F:��о���>�(/?�G�>�S�$꾌Pﾌp�>��Z?�?��$�A�[�)���>RPp?P�!��!�>�`?4Y�>%��׾u��Q:�?aھ��a�R�>Ԝ>��H=T�;��Ȣ�ԛ�E"�>���>ߤs��ڛ�z�>x�Ͼ����X�J��zﾟ��9��7f0?�$A�s�?>���D�=�D=�Ɨ���������N?��?��1?I$?	��%�W�kѻ<ٞ�>�� ?
��>WԘ���8���=^>�SQ��~�;�$?TG�?�?�=�?��}���ۿ|���*۬��̾ >�v�=��>و�e�>�Gg=�"���yu���>^k�>��d>KQ>n�/>;>�1>-ă�xh ��y���׏��96��_� ��e�u��3�b�X�����%��ҏ���̽�N��ɹ���C�����W�s�2Wj>�j�>48�>?��>�w�>�>�f���m��8����<��1~��)��u�ľͬe�&8,�|�'�����_��������>8�B��Z�=���>���J>�s�>��a=�*>��.>V�=X4>.t.>-#M>�.5> e�>+>���>"���lf��៿#�e�'��u�J>���> ��<.�c�i�(Z���{���?�G?N��>߫ʾ˓��l��/�>�E��7��\�e�U;�FQ>��>b:>7+I��-.����|;���>���>��2>�"����оR7(�}��>��>�f־�F�=�	�>R�?~p_?�*6?o�A=0��>�~>��]>(=�)_>ՙ~>���>U�?A�-?�7!?���>_�=�|�Z��=mS�:�	�c
$������$���b��;ѥp�]EZ=���<��5:�*�=}+�=���<�xv<O-�<8�?4�?iy�>��?`���Ee>��6(��z)����=�đ��ʸ>��Q> �>�B?���>9ot>}��=w�����ھ17�><�c>#�@�Rq\��-a��r>�+�>�Q`?�2?�=_�F�GR=#���.�>y?��*?���>�'>��_���E^ƿUH �)B���+���=z夽\2^�hr�>+�}=�vg�->�=m>�H>��>�+O>͝�=��<�A==�K�>Ѱ�>3�>�(<��`�����I��,�=��Q����X�l��`��jü�ڬ�������˼�
�}���aM�<l?{�?%<>�V�'�O#��������'��
?���>�f?V<?ev�>l{���a��m������B�>�#�?pb?D��[��>5���v�Ž�=�>>c5>Z;�<�y������ؾ}��c� ?B	?�Q�>G	��l���m����\�P��>�'=��Kl�?��\?k!�r�����#���C�{��m1=]ݽݩ_��Y���� �;{7�e����U�H=y�M��=� �>m��?�4����=AI��=�����������Vb=��h=���>k*L>��7�eۢ����T׾��O��@�<�Ę>����b�?n��>��?.��?dp'?�	�>���<?���m?��>�N�>���=�#�@ю<0$����<�o��2u�D@��2u{=�2�`�= (
>*c�=���g�(>�i=����ˌ��u=�Ϣ=��=z	>g�>Ȁ0>��	>[/?(L+>nŽk۬>�� ��J��==������@>��=`���Y3{�>�I?&?2�?��">�¯���Y1��[>B��>Y	2?�#�>��<��P��[žT��I����>�:�������ľ�<��u���ٟ>��6>\1Ľ��>_5�?+�(?���>4����3�0�0���UW���4Q���?�^8?->��߾y�q�1�������i�)#��N��L�=ދ,>H�>��>��=�D=�	�< =>���$��U��!V�>g��>�?㲌>���=�͘�o/
�P==?�P��<},��ꏽZ4���N�=]��<���p�<
7>�+���<�P��;�z>�>)Q�?���?V!�?m���nS={����@1�ń��uľ'�3�a�>ߙ�=a �>�`�>��>/��Ua>J*�>ob>�aR�X���h���n>#(��$���l�>���Kc���8K�K�(����=@߾n������4˾�"������%��`v�����)'Ǿ-�Ǿ�t�?�?�V�>aw����T�^�	����>%�+���˼��Ҿz����~/�l�ľ|����'��d*���	�af����>̒���P��v��RHQ�#f�_3=%F=?:d�珋���2�����0�>��K=�˱�kʌ�ï����z��A?(E?C���<����T<�Xj>e�??k�>a(�>´P��:�'J�=�h?�?,z�S���yЇ�����@�?v��?��R?3B���6�:&����ƾY??U�s?|��>t�2�x��[�v7�>�l�?]I3?wn4=�N#��A9��=>j1�?��^��V�>��>�J>���.k�c��->��Pl>��0>W�v>�T>��������{����_>�f$>\��5��ge�> ���Cʾ�=�=�;&X����=�'�>�g�8��=�X��)�����L���������(�:?/��?��?�@?�������m�>`��=��>�t����U�>���>δ�>t�����O���O'?���?���?�h?^*�ؿ=诿k�þ/�h�k�]=�~>z0�>ިe�H�=>劖><���Ϥ=�"?>���>H,T>:�>��:>��>r5>C����(�񰖿����Ai��8��H��������žOn��a3�(����Ė��h:<��=�g���qA�,]��\��h�k��4�=r�
?�	>��>j:�>�=�>֊P��*���� 4�x5羴t���#ݾ�;�q��PH^�@�^�g���ECz�:4#�RK<?]�=��>�s�>�=�>C�>��=2�S>U�=ե=0�h>��t>�>��k>��>y�#���>`��=N����z��/7�cmg��c��o?G?��P��n��Ǭ/�F�Ծ/����Γ>�?��F>�)*������S|�z��>c���[�U�ѽ�U��]z>ԝ�>t7=-&��D���yy����?(�=L��>��>��躍냾�:���f;���>Lu־���=�mw>ұ(?��v?+'6?�x�=���>��a>C�>���=iTL>z�P>R��>4�?��9?p�1?f2�>5.�=c`��&=�1;=��>��W��o������'��<��1���G=��r=h<W8a=]cB=��ƼU�;=��<�y?�a4?e;>��>�=��?�~IJ��R���=>ѳ~��z�>F��>]@
?[�?Q��>�>ۋν\�;�����>0�>>0W��*t�G 7�caF>;._>_^A?�!?����Et�`]�;���=��>G�?C�&?��>��=8+����򿿲��e�\o��:��:���=�>׾�ޣ=�So>�����t�>b�>D�>���>-:N>�8�< I>lӷ>�ږ>�=�8T�-
:>��'j4��<>����ｺK�=6�ؽRbC�e^���r�R���]ݍ;Ļ=�I=G�#?���>�wL���)�6*���V�{-��G�>���>d��>���>k��(�����E��zZ��x!�sȄ>��@?� ?u3 �{	>�s����½3�=7'>3��>�}F>v����g��b>J)?e�^?_�=?�v���HM�;�r��uM���p>�����*=С�?1=?��?��1�[E7���M�i��<�>্�BȽ���k���������ľ���4�"�`�?Q��?al}��V};�̾t��ƋM�Bj��$7�}�p>�>x�>����L���R��  ��kԾ�IU��I�>�����
?:�>��>���?�=�>�,�>*'��	?�=h�%)?^�>1��>�_?VF?���>P�ʽ��V��긽O��@_�0�������� >k[)>q>�����=���=*��<���0�����!���~f�=R
>�24>��>+{?�8?.1�����=�x�����$�-�kI�=�a>�G���uR�~�>�G�>B�^?|�=?�*�>�y9��uD���n����m>L�?��7?�K�>�Z#>?�=v�$(���!'����=�>��똞�%������_�ܽq>��>Ȣ�=��p>[�|?�#=?5�!?������.���t���!�А"�ּ{�>7�>7�=�ǾC�0��io��?a��_4������M���'=���=@�>�B>7��=��>ޮ�<�����+�*)I�5ڼ��>�<�>�"?3,[>��=�"���A�2\N?�y5��{���/><���$�>�2�򁁾"
M��7��{�;��s�տ/f��>��?�L�?A�?⊘��]����g>��=3�O>��U�6y�V/A���`={�/>&�/<��<����+�М<<�>b�G�x���h�w�c��<8����$�Q�>�¾�9��=�	�8x޾B�W� ����{�����-~��!὾��;6��p��O)5��䔠?���?�ó>ۣ@>77r���S��Y��;7>!�Ȍ<�����m�j���%��횋�������0�� ����Ҧ>v�W���V�o5x��^�H��"#V>:"N?M���!�=y�O�*>+��>�ڃ���D��Y������GZ�'7?@e?s��^�X���ξ�6�>�q?0�*?�J��&>�j�y�h>{�F?�7?�t�<�>_���Q��ʥ�v��?�?4�\?:����Ma���8��z�����>S�?��?_�3��#���uQ�m�.?ST?:��={X5��ax���"�F��>��k?I�>��z�>R�>�!l>��c�	���'��Ͳ*��p��d-�\?D�(۬��1�����C{�>Zc�>�	>�-�G�A���>���nJ���8�q6/�ᄯ���%>Y4?���w�C>̣�>w�>�4�2a��NN��*(����S?�?ra?�<?%��$B��g���"��=H$=?�\N?Y+2=����>gz�>��9�v���@���?~��?���?C�k?�A��Կ<����)¾�쾊;�:{��=���=@�k�7�U>Sj>ȁ�<��>��>���>x�f>VMl>/%>¬�=*M(>�`��E�#�>8��R蛿,|Q��1(�I?��z���о�Z~�� ���s�Mh��	���+�ʽ���3A���$�\O.������>�??8+�>��?���>�/h>������6�� ���P��ZO�������� ����s��AG��m�S��NW�r��*��>�VŽ��8>.�M>j؋� �=Ǝp>G��0�c���_>5H�=$ >	 �>#RU>*{>���>[>H��>V���I��������E��D���K>�?K�a�%�v�+U��m�៦��K?V|9?E��>	i��M���z@�9�>&D��Ҩ��&���%@���#>	�>���=]��=�QO��1���'>uu�>�Ƒ>/.=r8#��f���E� �>���>�IѾ!F�=��u>�<-?`Ux?"�/?f�<=j�>�G>N��>M?�=�0>XnB>p�>h]?�:?�1?s5�> ��=s�a�@s�<��L=W�=�4�z��eʽ.���⼝Ō<x�?�r)b=�(]=��<I�=�@=A����G�<t3=�2 ?D�?%@�>E��>�N���1Q�S>~��K���=��ؽ�w8>���>+J?O�?>�?7�\>�ֽ��¾����V�>r��<�1�� ���t�0f�=h(w=z|(?D�;?婯�^,[�e><'�<��>1�>��?�)�>Slh=�G�=����ο:�=�-�z=��т;�!w��bվ���>g4�<���l>�Y�>��X>oR�>dl�=B��z��;��=Ej�>>6�>�91>F�$=~G���2�3�=����\�I���<�����t<B�0��#6<=֑����0���<�J?\
?��콈�j; �T�t������:?�XT?b�E?(�T?�t�>�)ƾY�k��uy������e�>���?(�?�\K����>ү�=yG@�}��>Η=��7<�V���$ü�nd�|=Y>;�%?~TX?H�>&����#����%V����>	�>=���&��?��\?��������}.���E���	�r��=5�˽.H�ɉ��%@���0�T=�����~�q)Z=�?*S�?����ľ�=�`���ꚿn�������3�=��=ߧ�>�XX>�[*����}[���˾,�[�L�<�ϖ>�$�h+
?6? �?���?^ ?��?SÆ�B)�>e�P=(�
?Gs�>�U�>�E>�1�=Dn�P�k�Wĳ=BI¼��g����7=;ǧ�]�W=���=�9�<_���%�=d�l>e˙=i�<���=p�1>]s�=��=0XT>��'>�'�>�
!?x/|>˄�h�>�)�� ��sg�ey��쿼�2"�����Ⱦ��>��_?�lQ?��4?X�">�m۾�U�3-��6�>��?N[*?���>)�=J�>��Ùʽ!�=G��>x!���߾ǉ
�����ӽ�z�>U�j>(��>��?��?:�	?���=t���a #�qf������4>�,?�	 ?�>��׾��I�A��vo�RK;�4;���L��O>��>x�I>��#>��=>� >��м�@���u���T�$�h��)�=��;>t��>W�Q>\z�=�ͱ��A"�+7R?0Ý�v�6@��g<�>���>.��=򝸾a��>�^���9��#���f�O��>�6�?�O�?S�r?�8�h��s/=:^���T��:b; ��<C�/;���J��>zV�>bs������l>&A�>4̭>O�l�yx��e�����d�����W5���>~������F	��I��$�R�Xq�1o�<��&*���9�,�&� z���@p����į��p��}�?!�?��!>�W>��M� �C�>"�d;z=gd��/�>�W��@{�i������f�� ��!V�!���M�>����㬔�&*|�ÓA�:"�y��=�?��g��6��	�%��v�=J^�>)t>����l"o�ړ��C>@�d`S?^"4?�Oؾ]���ۊ�"�=�J�>on�>1^>R s������t�>}�<?d�#?��h�����Ā�u7j�3��?�-�?�YB?i}o�5VI����s�`��>�n	?I­>g'����Ⱦ��x���>_�A?��>��Ӿٞn�\��u��>��p?�X����>ij�>^9�>�Ђ�A혾�9���#��)����=�ME=Q��Wy�7H��GW�}>w:>��B�!C����>��Ⱦ=}T���j�PB������$>��?��x�?>3�V>:yJ=yIO��۠�Doy�����R?�C�?pU?g�M?6�/���H�P���!Wa>�1?�b�>RL��m�ѽ.+�<CO�>�`A��5�����-t?��?7M�?��y?�y(�~�ѿ�Ɣ��K̾z�ϾKx=�~�<���=��&��d>;��<�aF=j�=Q�Y>57�>wg>�K>�4&>P8&>D_>�o��ʿ$�����5����T�KA$�*��V������������(屾VY���������x��!C�W�i���_}^�5�>>v�>��>��>�;>{N>޳���@���Ǆ����\���?��Ҿ�{��w�>�������(���q����	���?	$<���=Q��>���$����>�=��>W�#>c":>Es�>�M>��E>ԜR>�
b>�B>��>������4����:�cӶ�	`>�@?ۮ���Y=�.qN����ds��&��>�
)?�>�����Q����K����>�m��d�)�" �J
:�H�>8�>E��=S*�"L=DV���j�=���>~>>̉=��Žm�ʾ�9�U�>�\�>��¾!\=��\>�1?�&n?�?*]=��>�6�=Q�=�9Ｊ��>E�>e��>:�$?��	?�<+?�	?3�=�Ss�6�;�T#=o$��<���G�j�s�<'��z)���<�w=9R�&	>S��=m��Q�'=C�=���>F��>���>R��>Y�"�����G���ɾ���:rPսn�=��">g(�>��%?�y�>��e>�s���¾@������>�5�=��s�������1����>��?(\t?V3^?A��=Tʃ�7D+�O�S>>DO?�"�>/��=ݹ>VRn�4�Gҿz�\�
�R�f�Yg�;�?�������>���=�˾=�O�>U4�>K�>���=�4�=%si�.�N>5�=݋�>n�4>�q9>J>�	���=�d�<4G�=֡=H\4>��qj���]@�|M����l;Jy�<gꑽ/hI���=f2?��?�����a^>���=�;����ݽ>9>9��=���=*p!?��=~�!e�ZK�Y4��,9?���?dݺ>+z��6>�X	>�R����>��5>�"켹g\�@*�̋��g����>�0?�A�>�k��Mh�����*��b�J>VH|��:�ز�?!�Z?��4�ݕ�@9�B!%���4����>�%���$�m���$�]�������FMY��j"?癝?��4�oe����sޣ��$h�_���`]𽁟j>/��>D�>0Rb���e��*���m:�ۘ��:eD=5I<Z�?��?H\L?Ĥh?���>�f�>|{=�t�>L]@�u��>�N ?��	?���>ϒ�>��s=}�t=�M�_\g��4/��ޓ����<�o=���=��/>uJ>��=��x=��=��=fEc�á��2=��b<k�=?�=�Q2=��Q>e?���>�)��X�w 3>tXk�����D�R<B��>��1��!'�0��؝0>�w?HZG?��)?g�����y�;��Ⱦ��>�??�6?�*�>����W)��j�����~>�v�>�>�"Ծg羆����&��<�>CD�=�&��o>bY�?�	9?9*!?�Do>N ���v5�i���dkS������?�+0?s0 >f��(�t��\���Kb�5��a�ܾDb��0ӥ=��=f�=_�=(y=,18=��>�Բ��F�[����FU>K�>#��>)?�gi>UY���Ⱦ�-���5N?��N3T���ξs���̛�>��?��>�! ��Y�>yk/=�(������v�$���>R:�?>��?�.f?!��=\Uֽ
�W>V�>��{>q}(>L����l��Y�<I�G>�@/��Z"�\����A>�S�>%d<>�"���b��8r��v:�E	��Q@�YSq=�����H��R�ھ��ھG���N⽧O�=^�������w��TA	�ah�ٶH�o����ƾ�ν�-�? �?�Q�>�>c �f�T�r����>���Gb�=���/u���c�ϗ���檾4�-G�J�G����D��>U��e\�-�~���N�ťz���=1-?7���Ә�e���@&>��O>����ھT5�����.A���I?�XB?��������I�1ls>� ?:�>�%> ����q��>��?��>KK�9y���8���@�<�R�?���?��??��V�*?A�6����ER?T?�i�>�l��*ƾG�:�b��>6�;?�A�>��u%w�J��e��>]W?@�M��qj>��>Z�>Y�ɽ����ҫ|�N=������B2>T��\뽻�L��g�d��=/g�>x�T>��I�i}��r�>����s�	�k��"�N��=̱�=xL?Qࣾ�w�>crV>���>����܌�ĭ�����5B?��?9O^?-�y?=|g��(�tG�nΚ>�?���>
'�>��<5��>�F?�V�`��@�{��>�n�?BJ�?%7?L��l�ؿ:^���\��*��i�ٻW��<���>Q>z=��]=7ȡ<i�[����:4;>>bm>��s>0�>��D>�]L>���=
t��/�W����{���I>�������p��9۾�I{�Y`>���������@�Խ�X��q���pd�E�0�l�O�
���-=�(�>.�I>|}?LǕ=�f�="���%��Ŀ����H�>��H-�����2���P���Ƚ��F���=y���Ҿ�)�>����� o=�>�m0>
A>P5�>uq!>�j =`�=S��=�'u>@P@=��<%��=�	>�rջɑ�>u��\q�V�i��m�8��*<��]?KU��0����B��Z�3�ݾ:�|>#4?`��>��1����c�K�_��>��}=�Oҽ�+*��×��ڨ>H�>���=��=��~��R������
>v�>���=�E��i}��K��Ć�=��>�Oݾ���=��V>�)"?$�?R�5?©>���>��?>+��>�,�<�3>�R_>Q�>��?R�$?(?� �>��=��O�n��<~��=_�M���b���ĽK�B��A���
MA�Y�<�ő=u�<<�E��';}�\�P3�<j�<���>�[?m��>�J#>g����*!�*��'C����=f�����>Ϊ?�?
	�>�ʲ>���=' ������<�S5�>���=x�O�t����z;�M�>��>��P?�^?���=q�����>4ؼ�?�`�>,�O?[��>~��>��=��AͿ��2��y)�!�n�z��E =�� �����W�xս�t�<��S>���>��c>��%>:�>�F >A_�>t�R>Ws�="k�=�-�<�ᢻ=���a���'��==%�~��2м�1E��c�ǿx��ؽ�_ֽz��������?��!?��H=k�&<�5	��e��վ�)ٽ��`>aW>��1>66D�5^&�<'�sR��˳���?���?�U$?�`����=��S���:��=*�Z>fĀ=Z���dS>�D���=>O4?`,?��|>��B��f���s�;��"��>�=���6�?*�O?>Ծ⁾F��)�:�,�j�*�2�F���Ҿw�Ѿ�`-���>��C��}��;cC���>][�>��?�����S>3�U�pI���ƅ�u%��7j�|+�S{�>:�>����	�>%��Y�J�<&�r>���>p�-����>�Vg?\؈?��P?��=?l��?���J@?��\>=�y?��/?.�f?�u?�?H�>��>{�>��^ �
�{��,���G�����=��|>1j��d�<�Y�<G�;��>�w�K�f�
���!��=�f�����<y:'>�>�r?�?o�
=�I�<�9>��}1�9��=��4>�%?рB>[��0��<�&%>X($?�"?��>��^>�飾�@��>��֝�< �?IX?�?��Ž�gJ>^=վ����U	>�8�>��B��N6�����h.R���z>,�f>�>Z�A=V|?�W!?���>�!���}��`�b�L�Y�ٓ��J�u�h�> �=���>M��?41�].��;�l�h�D�=�;����I>]|%>���<���u�J=}�t>5�>r�q�������=���ץ?�8Z>�/?��>������]�G���g?�]T�j�v�m��.(>�½=B0����>�غ�fv�>���L*3�����ݝ�<�?r��?α�?yj?+r��P	��3�>5$d>2 >��<9���B-:�8���=@򝾓*�ݧ������>F�?�0�=2���H�@��=�=ٿ��!���<��~ؾ����K�	��]��$Z��w�׾R�ҽ��<m7���W�0�ٽ@ý�ԥ�.T ���澕S���<�?�c�?g��>�F<����`"�p���|G�,��i�J�8�-�l���Ǿ�������N1��~"�n' �}(����=�a)�U?~���{�:�*�-&����=��>�Q����������</=�=E�>-�<����R��X���b�a?�WV?�k�U�{Ȓ��=jJ
?�:�>M?�>�f����5=�>��,?C�?a�8�����0.s�ӊ=�`�?��?'�??�R�͎@�t��2����?��?��>�l����;Q(��~�?@�8?�	�>=��ޙ��uO����>�]Z?�AN��Sd>.!�>,�>p2�����b-�h������M7>����k���g�S�?����=�%�>Qcy>�Y��ŭ�L�?fiҾM9��3PE�$@#�ϼ�"�x���E?�'�Ib(��W�>m��>*b-�Ӄ�����$=��b0?�ɳ?=�?�?�+u��;i�V;}S����!�&��>2<��(�|Ҏ>�B?k��֌��h&��I�>?��?�K@�͇?������ٿ�)���^پ��о�Ԭ=m��/�E>kr���	>��=ٵ_=1X���f=Z,�>#�a>�)>o��>�D2>De
>�e��C�!�"���ޔ�;B@�]�+����E!ڽ��n�>�y7�Ƶ�J���]/�=�X�࿕��o����R���/<N�2�ˢ+>,��>�D�=���>d��>:��>R���Td������&'���(��j�z�Ծ�������n���h��?��m�$��'?���=��%��h'?�z���=���>��>�_"=}��>��F>��>kt�>�=�>�a6=��.>�>P=���>ާ>�ᒿ
�M����6����j?Q����W��cM^�Aʊ���ھV!>N�>���>��S�ѥ��p��?�"�X�Ͼa����=r��>ʉ�>�m>A����=U���zž����d>2�>�!�<7ž�H/���&>�l�>��`�Ȣ�>�7�>69?���?��Q?2�=��>�M>���>��=I�>ݴ�>		?�
/?�^?B�U?/�>���<�5_�X=v��0\*�������3�兽ִ���R��� >A��=�m={� �Z�r>Ǎ>(K���=�=9x�<y��>�{f?���>�r1=rWӾW�0��Z�'T����=�=#@>$�?]��>-]�>��e>�sb>ae��m���a>�0?;[=�ד�X�����=�q/>��*>4}�?�c>?��>S3��]4�=Y3��ۨ> ?鯀?7��>�T>�N�=�����˿*�%��oP��־ф��0=qF�;x�3�'���s*=;\�
=0*>\�>��>"7>�,e>-B=O��=�;�>v�Q>���=Z>.�s<E@�=�|��;�g<���� �Ũ���; �<k�<�ν��X� �;���
Ks��?y!?��<�A�L��׽����4�U��>9\�>���>W�>�Z����@�H�X��%<�-�Z;8;?ȯY?k��>��Ͼ%U�;��K=S>>9?�^�>5��>�\��dま1�)�~�W��>C�C?g�>e!��S�{��pq��=��Li>���=��g��Ӏ?���?�������$������y ���7	��Sf߾�W征�� �k������S+���,��>�O?R8�?:��l&�>�r�E����$�����c8}>���=�Ð=��>�A�*�Q,�&,̾ݐG�QDʾS2�>��(>}�<�7?j�-?��?�HL?�S:?�s>݄O>��>z[K?�E>�0L?:�"?�":?+�A>�@>���>�!n<=	���h�����<�Ȧ�<��=���=mx�='�<��c�E�O�Y׽�s���z<��E�N�D���
=��Ǽ�t�=��?h�8?�d�}{}=E���B�p�8�=�N�>j*�=`kK�c�&>�d>���>3�?��>��>����{� � �4�2;}�?4�R??g?�|�=Z
�>a���$���5��L?>��;���X�|���W��'�o��>��o>�7�=��>���?�@�>إ?��<{�� �������C?�����þ��>|���R�3�\�e��K�&���g�� ��-C�F��>N�'>?�?���s=0�F>��t>^d>:QZ���=�0g>����ٸ�>$ �>5*�>oG�=5�>������h�9�]?�;ż����  ����UF����ޙG>�|�=\fN?�X�X�n��H���P<�a�>@��?�J�?�[?�VH�~~2�1O>>�2�>���>Z�>dD���k=��*�2T6>��<��4�����������=��=YB]�V)��sڲ��P�=Fڴ�YJB�^	��Þ��/)���۾5���n��a�P�V!\��F;L��Y�l��.�����Ty��놾f����y����?<,�?�Ό>bo> �A. �*�*���[��>��F�H�↾K96��ԏ�	���.���6����,���\��d����>��<�!���6)��n��� H,=����L?���S�D��3<��*��0�H=�L�����p�J"��L�žKua?0�??Y���������3?���?���>���=d�E��2w���?Q�=?�J?d�Z�2������O��=d,�?���?��??�O�D�A�o�����-?�?c��>u����;���K?'�9?S��>���g��f=� �>��[?�>N��b>��>0S�>S��Ώ��9�%�!/��rH����9>[�� ���*h�)	>�" �=��>gfx>3]�� ��L�?fiҾM9��3PE�$@#�ϼ�"�x���E?�'�Ib(��W�>m��>*b-�Ӄ�����$=��b0?�ɳ?=�?�?�+u��;i�V;}S����!�&��>2<��(�|Ҏ>�B?k��֌��h&��I�>?��?�K@�͇?������ٿ�)���^پ��о�Ԭ=m��/�E>kr���	>��=ٵ_=1X���f=Z,�>#�a>�)>o��>�D2>De
>�e��C�!�"���ޔ�;B@�]�+����E!ڽ��n�>�y7�Ƶ�J���]/�=�X�࿕��o����R���/<N�2�ˢ+>,��>�D�=���>d��>:��>R���Td������&'���(��j�z�Ծ�������n���h��?��m�$��'?���=��%��h'?�z���=���>��>�_"=}��>��F>��>kt�>�=�>�a6=��.>�>P=���>ާ>�ᒿ
�M����6����j?Q����W��cM^�Aʊ���ھV!>N�>���>��S�ѥ��p��?�"�X�Ͼa����=r��>ʉ�>�m>A����=U���zž����d>2�>�!�<7ž�H/���&>�l�>��`�Ȣ�>�7�>69?���?��Q?2�=��>�M>���>��=I�>ݴ�>		?�
/?�^?B�U?/�>���<�5_�X=v��0\*�������3�兽ִ���R��� >A��=�m={� �Z�r>Ǎ>(K���=�=9x�<y��>�{f?���>�r1=rWӾW�0��Z�'T����=�=#@>$�?]��>-]�>��e>�sb>ae��m���a>�0?;[=�ד�X�����=�q/>��*>4}�?�c>?��>S3��]4�=Y3��ۨ> ?鯀?7��>�T>�N�=�����˿*�%��oP��־ф��0=qF�;x�3�'���s*=;\�
=0*>\�>��>"7>�,e>-B=O��=�;�>v�Q>���=Z>.�s<E@�=�|��;�g<���� �Ũ���; �<k�<�ν��X� �;���
Ks��?y!?��<�A�L��׽����4�U��>9\�>���>W�>�Z����@�H�X��%<�-�Z;8;?ȯY?k��>��Ͼ%U�;��K=S>>9?�^�>5��>�\��dま1�)�~�W��>C�C?g�>e!��S�{��pq��=��Li>���=��g��Ӏ?���?�������$������y ���7	��Sf߾�W征�� �k������S+���,��>�O?R8�?:��l&�>�r�E����$�����c8}>���=�Ð=��>�A�*�Q,�&,̾ݐG�QDʾS2�>��(>}�<�7?j�-?��?�HL?�S:?�s>݄O>��>z[K?�E>�0L?:�"?�":?+�A>�@>���>�!n<=	���h�����<�Ȧ�<��=���=mx�='�<��c�E�O�Y׽�s���z<��E�N�D���
=��Ǽ�t�=��?h�8?�d�}{}=E���B�p�8�=�N�>j*�=`kK�c�&>�d>���>3�?��>��>����{� � �4�2;}�?4�R??g?�|�=Z
�>a���$���5��L?>��;���X�|���W��'�o��>��o>�7�=��>���?�@�>إ?��<{�� �������C?�����þ��>|���R�3�\�e��K�&���g�� ��-C�F��>N�'>?�?���s=0�F>��t>^d>:QZ���=�0g>����ٸ�>$ �>5*�>oG�=5�>������h�9�]?�;ż����  ����UF����ޙG>�|�=\fN?�X�X�n��H���P<�a�>@��?�J�?�[?�VH�~~2�1O>>�2�>���>Z�>dD���k=��*�2T6>��<��4�����������=��=YB]�V)��sڲ��P�=Fڴ�YJB�^	��Þ��/)���۾5���n��a�P�V!\��F;L��Y�l��.�����Ty��놾f����y����?<,�?�Ό>bo> �A. �*�*���[��>��F�H�↾K96��ԏ�	���.���6����,���\��d����>��<�!���6)��n��� H,=����L?���S�D��3<��*��0�H=�L�����p�J"��L�žKua?0�??Y���������3?���?���>���=d�E��2w���?Q�=?�J?d�Z�2������O��=d,�?���?��??�O�D�A�o�����-?�?c��>u����;���K?'�9?S��>���g��f=� �>��[?�>N��b>��>0S�>S��Ώ��9�%�!/��rH����9>[�� ���*h�)	>�" �=��>gfx>3]�� ��I��>�'����`d�l�\��Ͼ����E�>�����J>^��=>�x>�;S��*���ѝ��G[�\tB?�h�?��A?g�d?&zR�r�O�K��=}��E�>�?C\>bF�����=s(�>O���hw������?���?�!�?�bY?b|��߿G������E�˾���=�ɓ=�m>|��<���=��j=8d�<$���8l>��>��>_j�>�.>Y>2d>I%��&z$����G���V�%�@���[�T����۾�,�ҋ澮���)䦾�1���Z�8��T<¡� ���s���1D�ë�=X� ?F�g>�`�>�L�>�]=��#�����p���ϑ�:$������;K��Zb�X�d���ھ[ޚ��|;�f�)��>�
�=
�;�|�>P3����>M�^>�V�>���=y'�=b]*>���>hh=�H>f��=��9>��=��>w+������0r��!M�rT�[[�; ~?�%C�ڝ����H�9�/�:ꤾ��>\RU?���>ě�����̭����h>�7>z@�<j53j��L>�`�>%5�<i��w:�&���Ѹ0���+>��>\==��h-��2w��ن�=�M�>ؾw=�=wk>��&?��w?ķ3?���=��>QMU>��>䓚=R(D>��E>�x�>щ?�U6?w+?L�>u��=KSg�=;=t{�=v�K�%?N�U֗���޲N�vv<��;�o6�<��n="��<�.+=�:=�U���;<lV�<&?�.?Yf�>?@�>mN��<�rE�u	:�_s0>p�#<Õ�>j��>W?���>�˷>1>�z���$ľT/¾[��>��,>;�W�G�r�N���>'��>�E?D�6?x���������<5�>���>�g�>�.?{S�>$�=�;�0����ֿ�	#�s�(���=�a�Ҽ��;�D ��ϼxu�<�'��*峽;`>=y^O><��>�~>��:>��3>\K>�&�>R{A>���=C �=��<��%�+Խ��׺I�L��}<�n��26�<v<��-��O���@�$�ܼ2�μ�����X?�J?�qý8w>U񌾙/���9ﾔyR<V�>!�>٫�>�Պ=���O9m�M�W����y�>��~?պ�>�Qj�f�5>Z�=:�����>��>,>W>	�z��`E��¾���>W��>���>V@e>��<�㐿�Г��;����>�������<�?:�>�}i�� ���E�$M�ȠD�7��>�ʐ��#���"��S%�֡F������/e��������?��s??������y��9d����i�t������>��>�9r>�fD=ԙ��� ���'��Ҿ`�h�F�0>e�?8�a��(Q?D\j?j�\?��,?��3?��d?���Y�?n��>��:??�?�XX?��B?Z��>�p�R��=��&>B�->�.�}�'�N��<f�l�
��<�m�=�a׼���;���'C�=�'=�X=�瑽}���f=�%�=2G;=nR>�} >P�?S�>`88�"]�W@Q�Jꬾl�o>�~�>_�=!�����ܾ�"þ���=gy�>�3?Ԭ�>G��g�(�q��b���%<�>�%?"�1?HL?�ɸ�4�>Ć!�8��݃��{O>@LF���ܾ)��`�Z�;��}�>�	!>O�����u>uQp?�15? {?P����	bc��/�H�޻�J9�y��>Ip�>
nF=���w�,��Iz�NTa�<z0���(�<3����;�>. =�y>B>>��>�1�=����˶<����H�H=�I�>F�>��?Cǃ>_�O<e��2���qS?��*��JO���(%����@����x�=o����>m�|�t���m�W:�QU>���?�H�?�e?�k���,���=t��=�&�>dW=�g�w�X�!>���>�)�=�4(�<á��>2�>Cw�>#�=���῾Z�'>:�̿je�Е�=���[�>�ƻ��[�&n��'�3�GE��A���8>;��/����-,���N��ϾE����	Y�?0��?�>��ƽc���tWݾ�_����z��	^F����lk=Ө�V����N����C����Q��U�>�ړr�����d�����b'���x�>�
���c�<�����L�=HȽRq����������G�޽!�]?q8U?��¾�:E�4}-��A�����=�;�>皃>T�=SO~��ߑ>�S?c/E?P)l��ڊ����Sn\���?_��?�V?�F��=��B-�1���� ?�?#�>�>�$������4?Pjl?M�?�� ��Ą��2�T�>�?OlF�_l>�E�>o�>���ψF��%�=���=�c=��O��R��;��A���V�=F�>�]�>k;�>um� �3�L�?fiҾM9��3PE�$@#�ϼ�"�x���E?�'�Ib(��W�>m��>*b-�Ӄ�����$=��b0?�ɳ?=�?�?�+u��;i�V;}S����!�&��>2<��(�|Ҏ>�B?k��֌��h&��I�>?��?�K@�͇?������ٿ�)���^پ��о�Ԭ=m��/�E>kr���	>��=ٵ_=1X���f=Z,�>#�a>�)>o��>�D2>De
>�e��C�!�"���ޔ�;B@�]�+����E!ڽ��n�>�y7�Ƶ�J���]/�=�X�࿕��o����R���/<N�2�ˢ+>,��>�D�=���>d��>:��>R���Td������&'���(��j�z�Ծ�������n���h��?��m�$��'?���=��%��h'?�z���=���>��>�_"=}��>��F>��>kt�>�=�>�a6=��.>�>P=���>ާ>�ᒿ
�M����6����j?Q����W��cM^�Aʊ���ھV!>N�>���>��S�ѥ��p��?�"�X�Ͼa����=r��>ʉ�>�m>A����=U���zž����d>2�>�!�<7ž�H/���&>�l�>��`�Ȣ�>�7�>69?���?��Q?2�=��>�M>���>��=I�>ݴ�>		?�
/?�^?B�U?/�>���<�5_�X=v��0\*�������3�兽ִ���R��� >A��=�m={� �Z�r>Ǎ>(K���=�=9x�<y��>�{f?���>�r1=rWӾW�0��Z�'T����=�=#@>$�?]��>-]�>��e>�sb>ae��m���a>�0?;[=�ד�X�����=�q/>��*>4}�?�c>?��>S3��]4�=Y3��ۨ> ?鯀?7��>�T>�N�=�����˿*�%��oP��־ф��0=qF�;x�3�'���s*=;\�
=0*>\�>��>"7>�,e>-B=O��=�;�>v�Q>���=Z>.�s<E@�=�|��;�g<���� �Ũ���; �<k�<�ν��X� �;���
Ks��?y!?��<�A�L��׽����4�U��>9\�>���>W�>�Z����@�H�X��%<�-�Z;8;?ȯY?k��>��Ͼ%U�;��K=S>>9?�^�>5��>�\��dま1�)�~�W��>C�C?g�>e!��S�{��pq��=��Li>���=��g��Ӏ?���?�������$������y ���7	��Sf߾�W征�� �k������S+���,��>�O?R8�?:��l&�>�r�E����$�����c8}>���=�Ð=��>�A�*�Q,�&,̾ݐG�QDʾS2�>��(>}�<�7?j�-?��?�HL?�S:?�s>݄O>��>z[K?�E>�0L?:�"?�":?+�A>�@>���>�!n<=	���h�����<�Ȧ�<��=���=mx�='�<��c�E�O�Y׽�s���z<��E�N�D���
=��Ǽ�t�=��?h�8?�d�}{}=E���B�p�8�=�N�>j*�=`kK�c�&>�d>���>3�?��>��>����{� � �4�2;}�?4�R??g?�|�=Z
�>a���$���5��L?>��;���X�|���W��'�o��>��o>�7�=��>���?�@�>إ?��<{�� �������C?�����þ��>|���R�3�\�e��K�&���g�� ��-C�F��>N�'>?�?���s=0�F>��t>^d>:QZ���=�0g>����ٸ�>$ �>5*�>oG�=5�>������h�9�]?�;ż����  ����UF����ޙG>�|�=\fN?�X�X�n��H���P<�a�>@��?�J�?�[?�VH�~~2�1O>>�2�>���>Z�>dD���k=��*�2T6>��<��4�����������=��=YB]�V)��sڲ��P�=Fڴ�YJB�^	��Þ��/)���۾5���n��a�P�V!\��F;L��Y�l��.�����Ty��놾f����y����?<,�?�Ό>bo> �A. �*�*���[��>��F�H�↾K96��ԏ�	���.���6����,���\��d����>��<�!���6)��n��� H,=����L?���S�D��3<��*��0�H=�L�����p�J"��L�žKua?0�??Y���������3?���?���>���=d�E��2w���?Q�=?�J?d�Z�2������O��=d,�?���?��??�O�D�A�o�����-?�?c��>u����;���K?'�9?S��>���g��f=� �>��[?�>N��b>��>0S�>S��Ώ��9�%�!/��rH����9>[�� ���*h�)	>�" �=��>gfx>3]�� ����>�微3J���B�S�	���7�v��;���>0i��q��=�pD>P��=:E+�o򍿬z��<}���D?>�?�]U?��/?|y��fݾӟ}�L��=���>���>ɣ�=N�0N�>�`�>E���9l��R���?;�?Ր�?(P?��l��Կ�����%����5�>!��=�8�>�����>> o>r��=Tqý���=Tu�>KC>k�3>Z��>Nd�>}5�=�a~�n!������s���Fx����)Н�DI���нgD�NZ��y���gI=�ޞ��hh�� ����Qp���[����=�B? U�>�ZY>�#>̤�>�m��������� ������
�C>��X�"Y4��Jf�0�ܽ}#G��k���;?,�*=��>�?��=Y�z>���>lp->S��=�Б>�i>�>2-m>�P�>N��>�/>k�3=Lͷ>�T~>>ׄ��܁�cc&�_t��@R�̓2?�%�
�j��)��т���?�	��>��?­�>R���ȕ���~�7�>�ؼ��W��XT�=o/o>�#�>#�=A�V=;�=�0���B���q>��>NI�>�>��P��H�w7G=�s�>���?��>�a-��uF?�x�?	Z?�e[>�_>�7x>�=炊>`P1>�K�>�ސ>Er&?�9?,�?i��>+0>��ɾ4�=�%ͽ��o�=�����=_P��<k>0��2>�R7����+;>�@����ݽJ�>q{>b�?�|;?L�7>aY�>ȹ���J��IR�ȣ=?��=���V�?1�>���> K�>h��>d��<�i!������;��� ?�0T>��l�n@��ge���$>��=�~+?�D2?[�>Dw��{�4>lbv>P�>3��>��\?1 �>�*��c��?���ٿ �H��|�aO>�>��z>BZ��Co�>��>�%�nG����=�3?2��<�3>�
(?�po>u6���%�>,JB>/�=n�	>~����[�ڄx�a��= �{��>�<��+=֚����->�Sʽcｌ��;>SG=3o7�O�Z="?ۤ�>�.&����-�۾�!����X�?���>�F�>��>S�ź�&�19`���R�����7h>x�R?��(?�?���>�w�,.�;r�>t��>���=�t[�q�e=�����3���^�>KΝ>8s�>�z�_q4���l����R��>(��=�z+�֕?6�c?���������c��	E�nK�=3������Wľ��2�=�,��*��k �|;>��*>/?��?N����r=�\
�gT���en��=o�K)�=�̽-R6?��>ML�L"	���8�5��XԾ⨢�L?�>��=p�>�q/?N��>�ӂ?�\E?47?�c,����>��u��Z�>�?l�?o�?��?�<�>ٞ�>�mc��/�����h��y��݀���>�;o>S<=>W�=j�j=R� >�B�;��v�e���<�Ž�7g�,�=  |>���>� ?G�A?ؽ�p��b�X>z�w<����0O�kx�>�x��Rڽl��>i+?M/?Ȋ?�Q?D� :�!Y��@����U@R��!?�?��?V\>rk�>��Ծߴ�?��ǌ1>��f�� >�}󂾌���wY�C��>��>c�o<��>$o?q�>�};?8p�;
���k���-���2�������>i�@>�$���! ����eL�4�����Btt>��g��UҼ!�G>��>�8�<	su=�$�>��=�eV�;@b�Om��@hN��U?Bl�>��?۰<>�o�=3�����)�I?����i�.�sоWZ���>1�<>���?��s�}�g���H=�>��>Y��?���?�>d?��C��)�E�\>5NV>��>|;/<՚>���䈅���3>��=5~y�����F�;P]>�Jy>��ɽO�ʾ�1�H�*���@c�.����
����{���Ǿ)Խ��¾�u$=����j�ξ�鍼��<����v��I~��W6���þ���?�W�?�k�>)���U�5�9�s�.���>+�$��%a�@������V���)��&w�n�(�P)�����Nm����>�\��琿1|�)4��ơ�>�/> �;?�.��V���2���=<�>��߼�� ������<����Խ��]?�15?G�߾�J����޽	�%>��?.ӻ>��=�As�4�$���K>��4?�H?��Ƽ�H�����=�D�L�?�o�?��F?I:�6�J�|�
��O���C�>uZ�>���>|/�b�������>���>Fu>d�(�:i��E8+�=�?��w?�����c>� �>��>�H�=��8�`S[��
�r�����	>�mC�NT8��|���n��=���>�W�>�N�S����>mӾ�������&��7��u�=�b�><�!�� >�M'���G#�a���â������W?=��?��V?��_?k����<�|���� ��>�>�O�>�_e>�9�>O�F>ؚ>?az����2�������>�?h�?D[�?}�R�߲տ;)��k׽���ɾ�t�=���=��q>��>��~�=,V=盯=sa���5>��>ul>O�>��|>>%9>T+>�3���!���Fv��!�;�W�! ��y��,����b��8�¦��õ����E�x�c����w%��:���;}1A�e�&>f�?�>��w>r}>�U>�Q;�'c�C�������m�qb.�n~��@��c���[}=�V��u7��`����/?ߺ=��P>�}?�t�=�|?=��>c%=��+>-�\>�i>���>��>�,�>؈>�r>��yj�>���=镅��ꁿCi1���7��'���A?�H�����Ԟ,��J;@!��1��>�?]�f>�Q$������~�>�nD�',`��[���߻��>�>�J�=�¼)�ּP�p���ڽA��=*�>�>�yM�g���<�%=�=Y!�>���ݎ>f�f>��#?��?��-?'M��nh�>Qu>*">�N�=$��=T�F>��X>��?��3?��4?���>�>>�閾�AV=��=���Z�<�R���Խ�4ѽ+_Ͻζ׽==�x�=���͜�=�<w;-A��5�=�=w�?�[?^c>�?�v�2#���E�&�����>��/��
?r�%?ٖ<?��?�+�>�7>��u����$�t��>���>�N���߆��=U�>_�_����>'�?�
�>��&��>#>�\?�?7O?+��>@��VJ������,�ſ����e���<I E>@��>:c��X�Ｐ��=|U=Z%��鰽���>���>g�>��>��>���=�-�>�$=���=���=���<+�<�X�:Y�=�g=�բ=Xͽ�߽c�/�p6��Ͻ<C�ؽ�;�������֦/?d�>Z�����_�����w�%�?���>��>U�>q�������i�T_�����*��>FP�?e�'?>g��ػ�>l�G�$dK<(�>�7H>v��=�TM�߫�������c�4�>b�`>��>e����J��T��a�P��>���=���w�?�-]?�s �?|��:��0�w�H�0�="��t������>-+�(03�Qb,��"���J�y�X>�W-?x�?��达�G>�v�-����mw���;�K9���7q��>��I������ $�,�v�> ���Ⱦk#=���>����6>\	?��?��_?�~*?Bp)?[�M�)m�>�>OZ�>t�>�r�>�k	?�9?�Ѱ>_*�>���<�ۊ��N��6y���=��W���	=̫�=l$'>����,��=g�=�����W P=��=i�(=��w=Q�8=9�>�WN>ϫ?�Z?%�þ�о�<?}t�=���b��>��O>�	>��0�;�?��1?�\T?�Ga?��6?��A=��A�fp^�b�����Ы?���>��'?Y�b�`M|>NwB�6R��\4�=�E�=at׺۫T�������S�Mz�nV>�w>�>+:�>�{?c0?%�M?���<H>�[�K�Et־D
�[Y�o7�>T��<E�����ž����`��XE������8>�e��D���*>)�>�uV>�]����>e�>��>�7I�S�� �=��?�M�>�I�>_�e>l>J���M龲�J?Vf���,�?Т��վ�<�>�@>ij �֤?���}��<��5P?��;�>KE�?M~�?�'e?��;�E���U>�I>�^
>��;= A�g"�:CC��?>���=�g�������;Il[>�^{>]�ͽ��ʾܾJF9����7�S����ҾҾ����O���RXf��΍��0N��[����4�"���W��z��<=�� n��Xž_������?A��?�΍>�g�=ĄW�{�E�����<6����<�-Ѿ����_��Rb�K���%�$�L�'����(�r��Λ>��Y��?��W�|���(�����b�?>9/?F[ƾ\´� ���Bg=�H%>/կ<PJ�懲������
��bW?��9?�H쾈:���S�)�>��?�v�>	�%>���"�<�>_;4?c�-?��뼏��s8���p���i�?^��?B?�(�oB�uv��H��T�>���>,9�>�!��Υ̾Ւν޴�>qz$?R��>5�����T���.?��`?���LN�>��>c��>�Ӈ�]n����*��ݤ�����=\꼣�)�����s�-�h�=��>hY>N���󉡾l��>M��YXL�G� ��mc+��,<F]?�����u>Cr>0�>��(��\��4{������I?<�?�~Q?S�;?������id��A�y= �>�.�>hҥ=^ �F��>���>,�is�5��N�?¶�?8��?��[?rci�BGӿ����������=�$�=��>>��޽�ɭ=��K=�ǘ�Z=�p�>}��>)o>K;x>p�T>ț<>��.>o�����#��ʤ�.ْ��[B�� ���wg��{	��y�����ȴ���6�������,Г�y�G�e��U>�Ɍ���\<�u,?e�>��>�.y>�`>J�b���-�5��E�8�[����L��$��n�����d_�Kdӽ"�����C�P���m?��K=l�d=W�?w��=��㺪�F>A~���J>��=,@����>��=�f�>й�<+�D>
�=�a��>���=4����~�7)@��(o��`<���-?G	.������b��>žH��΅>#�?j&U>�\#��ȏ��Ӂ��U�>S%��w�-S���%�t&�>���>~�C<uͻRy�;T<����Y�=��>��.>&�y<�}|���=�i�+=��=�}��t%�T�F�┅?ZӘ?�y?�>�A�>�1F?��>D���,�>�g8?��>졽>�)�?�! ?�ǭ>��9�#޾��X<��?��8$�н;t�0����>��*�3�=d�
�Sޠ=��X>�>���>��=�<>��=���=�P?�P??�>q�>x㤾%�`��sD�����>�����?��?C	?ߣ�>�U�>�z�=� 6��S���.�Rp�>0��=F(v�����%u
��% >I��v~?Ul$?�>��m��=��<>� ?@}&?ͳE?蓴>u��<X�㾿3�+߿�@�v���;c���,�M�=ϟ�6;��Sڼzth<�tH�4d�=X6>�]�>�«>�Z'>���=v�=3��>?�.>	��<�/4>�K��#g�'3�82
={���I��xP$��6�Ӓ����罕ʽD[��ڼ��%�ݽ(i*?Х�>l���'�݋ھ��˶��m�>tZ>�:P>���=�=�".�#b��F\�[c�p��={A�?��>?^}��%zC>v&>U>/��>���>�:c>��Q�[��ľ�ٵ�]8�>�?�!H>N"�>Q�a�6��	��>Q̙=�2%�?��?T�Q?W��ʌ����;���:�p��U�d��v��o��@�5�&�@���(����<� �=�O/?�X�?� ��N�=:��Bi��4 }�[1�rƒ>���=
�?_�7>&�
{��ǂ$�{�Ѿt��}�0>6��>��=i�>�Y?v�?	j?�$?f�?Գ"� �?��1>��>��>�?�z?P��>4ۀ>�5�>��w=	�z�e<�귤�lQ�;�J3��s>��;>S�<>��;�LH=W�=�E<�����޴�<�QG�k֊�7��=%>k+>�?�]?��� lA�U�="�F�h��ʺ��a?�4�E��C��>H��>yN?�b?�]?lҽ˳k���9��7������>�1?�]&?��A>��]>K��������<d��=���r���axQ��K��47�e�9>_h�>�/D>�v>�z?v�M?�w?�k��D����۾S�%�[ޣ��N^>���>��8=qN�&rK��x����d��/��m>ɭ���j9>Nȏ=�
8>�_l>>)�VtT>�|1�1z	>�)��BiĻ���=��>t��>�P�>hb>7��=�+���߾:�I?ݚ���j��|tо�a�?�>��<>����?���/�}�8��tH=� ��>���?"��?�>d?2�C�M%��\>�FV>��>/<�>���l���k�3>��=q�y�����Ԟ;�]>_Cy>n�ɽ��ʾX/��xH�L���tkP�{>�w������㾜����jQ��"*��t�i�ž^���b����=� ��0��������ᾧ1�?2��?��K>X=qR�b�'����{�>�8�O����]����0���>"�'z쾁\2��K����|�͞�>Zk\�;���b�z���8���M�>�H8?w���&�������<�=a�������Ȇ��̓�����<
H?��B?�߾���>A�A�>��?@|�>��=�e�W���.>t�;?j�?��ż ���?����	Q�?P'�?+�E?�=��dI�� �j�M�~�>;�>C�>�vm��x��>�2�bg?s?�M�>E��6���D��?�b?�(��ٻz><��>W٪>):��W��ߕ/��`��DF����>*��ʢ��`C��k2�S��<ʍ�>i_�>��C���n��>m᾵mP���F�����C��7=�=?�W��L>C�g>=��=c�*�����sӉ�4�{�;?zҩ?�dV?�:9?)K��r���.�~&�=9��>��>���=۲����>͛�>�徒�k�����R'?�=�?͓�?�t`?��W�	�ο�	���S��S����6>nj(>�;�>�ýM�d<E��F2D>��=>�
>���>9�6>*kV>��w>r�>>6�>��{���'�VT���u���/�60�����>x�s���a��S�
���Hܭ��	:��̽�M��hh������a�%����=��C?��\>1�>2�>gz]>��۾�kپk��W��1���J+�����z��� ���Y���ｰw8�b@�_U��x?3=���>�5?@e�֕>x�+>,���w��>JV>��M>��>@>b�l>c?>�(i>n�&��֟>.��=����7�v���G��^���J���J?��B���@�N4��Ѿ�����A>�|�>�8U>~.��s4[���>���)�|��:%��C8=䄥>���>n��=|��=/��R9��hA��C�=��|>D�*>�C�=@�V�􄽚�2>5�>�yؾc�>l�i>Ň(?`�v?)�4?4j�=��>��]>�T�>C�=�?9>S$G>� �>�%?�8?{D/?H��>M%�=��b�hU7=��K=)A��>�q�½���Q�y�Ż&y޼��F=�i=�t�;��M=.�<=��ӻw�<X��<�?�N?d�!=��>�`��uC��i��>.��>ph��9�?g�?|\"?E5�>�>t�/>�짾�V���.B����>TG=>'�l�|��&�<�rO>�w�<��F?�2T?�B��c��A�?J��>u׾>#�F?�bv?G�>�����S��4Ŀ���4�%�Z�>�H�E��>Z���]�>���=zb>C���#�G�"�>�"�>$�>+" ?��>�[ۼβ>�Z>|	�=P霽뽿��<�_H�CN�=1���t
0=����9�޽�6�<��нAB�=��<�B�=0򞽖�</1$?g'?��<��+��Zھjw��5&�>�e6>��>�Ѓ=]F�ֵ"�q9l��iV�E ��0  ?Ȃk?5yS?𬙾�c�=m0O>�Vd=��>���>�K�=����F#�呙�]K��k#�>���>���=�_���U�?�H���Ծ�+R>�8>�\�z�?
NF?�j
��៽����u8�E�O�o�Z�xF�A�˾�ܾh^!�ռ7���n3������ҝ>s�?:c�?s���\T>��#�p�\���w�N�x�=�Y�>oa��� ���}���/���ܾAp>z��>�_=�X�>�+?��?Huw?Q�#?	 ?`:�/� ?Q᧼���>=��>2�?�?��?�'�>~�>W��H�����N#��>�>I��B��=ތ>��>�>�eC��;��[(n<��4N����VY=1��=%x�=�޹=�?�9Q?����#��<��>.\`�0$@�k�_>MV!?L�#�t�˾��>@�&?�AE?U�?��E?Ɔ�RL�q}�Xg�.�;N'7?G�?Ά�>�O�=�U�>~�`�D�I��=f3>%���ݳ�����ج��NU�hM�>?��>N\>DC�>��j?G.?�Dq?)r�� |���i�[8�3�H��<ɽ���>���=mY�;�
���2��!}��"Z��l���.�"+^�+�=�EH=��>�q>i-F�X�:>	R�=�5=:��=��`>D�=/i�>ׂ�>��>�F^>��K>��쾣���I?Ah��\f�� ����о�"�;�>��=>M$���?�a��}�����f=�f��>�M�?���?�$d?�B�wP���\>r�V>��>�f=<>$>��8� �����3>(J�=�%z�鋕���;�:\>y>ۃɽsʾ6���E�UE��5�R��O���~꾺q������I����<����ԛ�맚�^dw�g��I-��U�b<����x�c�M���gw��Ts�?�W�?�;>�>m�J�a�5�����>���S�=+���Y�O���}��[Y龲�.���%�=a#�Z���L�>��D��9���@o���?��	�bA>ۋ0?A�ܾáM�R��-�6�1U�=���������g藿���~�U?��D?��������8��3�=U?(��>�g0>K��h���tb>�F?d?c�Լ�����Ey�����z�?�^�?�sE?�=���$�#��l���m�?qʿ>��>4���5Lξ|��"��>V�?:��>$��`���A*��/?�Ok?�gI�Ԏ=>!Ȟ>�2�>�c/����0"H���`���:�3�/>���<1�!��펾��>,�>AP�>:`������%b�>�R�)�M��'H�Л�Pc����<�?����ţ
>h�c>g�>�c(��5���܉��
��!K?��?#�S?�r6?���ʯ쾧ѧ��N�= Z�>���>O�=y7�ú�>]I�>�G�U$r�?��O?HA�?Ӷ�?͎Y?��m�}ѿ�@��=î�Vɲ�L|�=�[�=��D>4齙��=�u[=�J]�\������=��>Xc>�s>FS>��:>�C*>�ہ���#������{��FB�dl����EE��!�	�g�}�@k�O@����������&��3�����H������0��嶾��<��?O��>e�6>��?>Hl>l#������W�R	�P�7�����#�����?]���5n�=�W������;X��H����>?}t=&ͪ>�y?A��=;��>���>T��� ->��<���=K�>��.=�
�>��> R>}����>;�2=��l�pvz�%J��%���� �j�)?�Q�gǯ����H��p���Q>{F?��=�� �����J�q�y��>�щ�
�j��J�;����M�>���>"ǜ::�,�[��;��\�6`�!���=2�Z>w�Z<����IV���> \�>���:B>]W��+e?��?n�_?Tמ>��_>t�Y>�w>��>���>���>5'�>ׁ?6�t?u�?"k�>Q�>O����w������G���އ=ð��v<ʙ����>�����,>O@>�F�<Y���1�=I�Y�(q	�n���^?b%?�+>>��>�-Q�iC�P��bS=�a>~ڹ�6b?'�>�i�>к�>-T�=<�>�~�������`�����>�U2>p6y� ��8΅�(�~=��>t6?c�\?[�<�q�|~�>�b�=۹?��?FQA?��6>�_D>��ʽ
����Έ�&��/�	�<?�{;��>��ν<��/�����G|>���=ٛz>�ԧ>�+�>�!n>��->�W�>��>{P+>v������=��<��:�d������=B�e�ͧ��D���x��2K������� ���g�k2��g<�����?���>��E���=YbɾG��;{쾚��=�>�@�>k�>9B��:�5�1�c�cf4������,�=�d?64
?��?��=�~����=c��>C�y>��v>V���u�.�����=��{>��5?0�>�dn��!$�R�=����[��>Z�'>�֔��?�fg?���a�
�?��t+���/<+<\��sH뾪 ���H�QnL�ן9��Y����,>��l>��?ef�?nG����=����옿�y�������e>�a>��?�$�>�B��ߢ����K�� �zw�>�5�>{����x�>�VF?x%�>)>�?W�4?�eW?E=UC�>h�^��X�>���>788?��(?�?��>ma?<PI=�L����A}����=���1M>�6�>φ>�	�=�?O>v��='C�<����#�֣���
���হ<�,�>���>�"?�b?���d�=�����_�Hwɽ	+.>:��>��f�?�ü _�>���>�'?!�*?�ME?p��=F�C��� �"���=�c4?��?e�?a�]�i2�>"Q㾜�o��W�z�,�p"����$G��-��=��<�y�>��=/�Z�>b?�B*?%t-?
�U�%�DIv�012��I�1~<E��>��;>�a�5D���7�y�l���m����c��<Q��h<�Z�=��V>D�=>Ie>;�V>չ3>*x:��W]�;�8=��*��?<��>x��>��r>u�Y>X��`��I?p���k�6࠾xоP[���>O�<>l���?���%�}�^	��<E=��~�>F��?��?/<d?��C�
-�b�\>oAV>��>�/<8�>�[��MY��x�3>���=�py�+�����;I]><My>�ɽZ�ʾ�9侚�H����9��G=_���|c��Y?	��1��$����%]��Z&<,*��ߎ��d[�!�׽:�>�8p���	�]"l�z��,��?�\c?Yy>�ȽM�r��_�//�I��<�td� �b>�+Ѿ�馾 ������4#þ�G;�xS����Rj��,�>��R�����u���)�W�d� �>�?�ʾ��������o=�>\�Լ�s�z������������^?�S(?}��R�͆Ľ�K+>�?Q��>���=	�����ɽ`�t>'�.?�0?$c�S���:	��DZ@��5�?V#�?:MS?m��Wc����T4@�%>�>HF�>��?{���t帾�$(>��?��+?-��>:����a�3#��l�>�F?G�B����>��>v3�>�	��tv���MǾ�k~=CS>r��������y�ԽB3�>�(�>Ťg>����Bо���>n'�W�N���H�z��	���<�?̑��>�2i>35>.�(�-��6щ��F�T�L?��?BzS?=w8?�_�����i什��=�>��>���=�����>���>�辁nr����?A�?E��?�LZ?Ƌm���ӿ�娿n[���̾��D>��>AE�>Z�ǽ��=舵=C2���!����>'��>��i>��>�ͥ>犄>���>�B}�Z� ��f��[�t�X�A�������� 	��=�'��fw�(��6�о�i���=��9����@�=�V
˽��C�) ���Q佃��>F�*?n�>���>��>1��½x�	��<�b�.+P���`��^ƾk̾���E\H��W�ݗ�U�����ﾜ��>��Ȼ�T�>�v�>�8��X�>	��>��<��H>}p&=9�����E>�����>0�>�K�>�>>�K�> ��=O5�����BU��$�hD�=��H?����ƾ�h��I;=�9�>�_�>�uϼDW�k����-���
?Ե���Ͼ ]�=*����><w?�y=xT=��>F���LN���>�<�>�A?]Ê=o�=�gǒ�}�="_�>�\���8/>���>z@?�j�?%T?�h:۱!?�v�=V��>�,�>-E�=0*s>��>H�*?�&_?�"?��?�cD=#5��6c�=�3J>�`=���=[�I�N���ϼF�F=},� ��=af�>x���=A/>݀[���[�)=��>��Q?�
?S�>�t���@�-��� ^�u��8j=��>�!�>��?U��>I��>���>�k1>T����$��
�>��n>�Z�����+��{I>���>9<D?J{)?�Ň=f�[=]~���V/�8]>d��>�^1?���>t��>.P>Ͱ	��ֿ(Q)��K�7�O��Q�r��<��N�w�w�^���i;�I�뽂�<"l>7[�>,�v>�FJ>�,.>�S>a��>v�S>?5�=ױ�=O	������1���e�<`|t�3
������"��<݃]���½"������]���7����`��?W`5?�u�<_.r�M���p��?����8?O{?e?{�B?��=�<��}N�I0(�<˽̠?䭋?�0?R�1�"=��B���=��c�>�׿>j�>>��=�}">����Kq= �z>-+�>�՘>�H�2�Z�uP��n�Z��>�t;�`���[�?"H?��Ҿ�m����.�HA2�H`���@�Y�l<�`��:����"��BJ����hS���B��M��C��>��?�~������8��h�h��[޾��`��=�	?$��>Tu:ޡ\��z��-�f�j�(��P=8��=�LD=w��>F=A?�5?��`?�S�>}_>�7��6_?E$�=Iپ=$��>IK?qA?�?��>�"�>��>f��=$6� (R���<������>9�q�ō�=l�=m�ѽҿ>������j1>^u���s=�&>C����E>M.>�F�=��?H?�-D�,�=9Ͼ���?ֈ=���2���^=�lh�ؐe=6�Z>�Л>b�^?D�^>��3���w�V� �=�)?�.R?��?��=�(��a(���'�iǎ��=~�m��<��޹�S���ƥ>��>�ܡ=�$b>��}?}B?�!?א���"/�$�w���*���ü9���r�>���>�I�=&�ݾ�7���r�T1a�G1��eS�A C���	=���=��>�>>=а=��>�&(=L��M�ս��Z<2*��a�>���>�t?�%[>�=�ĩ�� �~�I?�נ�M�����EDо���+�>J�<>���/�?�
���}��⥿i=��)�>���?���?1;d?�B�t�I\>-�U>��>'�7<:=�Z��⧃�ٺ4>���=L�x�	H����;t\>�|x>�Ƚ�ʾ�9�kbC���ǿ�	h�P!����׾�P�[r���:�j6����ξ��ƾs޾�T�������aXA��b��૾�����=���M�?�N�?���>K�(����՚,���6�3c�=����0վ3.���.����%�����8���q�� W�2+g����>]�S�>o��rC}�~�'�;߼�D1>�w.?%Fɾ�C��^���t=�+>�<�+�jc��SA������T?	�:?e��������
>D\?�1�>M+>d�������>;^1?�%+?0���͍���������?�}�?�W@?��O���A�f��Bg���?�?-��>;c��{�ʾ�n�Q?��8?4�>�9�o����"�>�Z?F�O�a�a>3��>�ՙ>^a�����1��r��)d��o�7>�	�#��,7d��NA�'�=A�>Now>�]�{I�����>n'�W�N���H�z��	���<�?̑��>�2i>35>.�(�-��6щ��F�T�L?��?BzS?=w8?�_�����i什��=�>��>���=�����>���>�辁nr����?A�?E��?�LZ?Ƌm���ӿ�娿n[���̾��D>��>AE�>Z�ǽ��=舵=C2���!����>'��>��i>��>�ͥ>犄>���>�B}�Z� ��f��[�t�X�A�������� 	��=�'��fw�(��6�о�i���=��9����@�=�V
˽��C�) ���Q佃��>F�*?n�>���>��>1��½x�	��<�b�.+P���`��^ƾk̾���E\H��W�ݗ�U�����ﾜ��>��Ȼ�T�>�v�>�8��X�>	��>��<��H>}p&=9�����E>�����>0�>�K�>�>>�K�> ��=O5�����BU��$�hD�=��H?����ƾ�h��I;=�9�>�_�>�uϼDW�k����-���
?Ե���Ͼ ]�=*����><w?�y=xT=��>F���LN���>�<�>�A?]Ê=o�=�gǒ�}�="_�>�\���8/>���>z@?�j�?%T?�h:۱!?�v�=V��>�,�>-E�=0*s>��>H�*?�&_?�"?��?�cD=#5��6c�=�3J>�`=���=[�I�N���ϼF�F=},� ��=af�>x���=A/>݀[���[�)=��>��Q?�
?S�>�t���@�-��� ^�u��8j=��>�!�>��?U��>I��>���>�k1>T����$��
�>��n>�Z�����+��{I>���>9<D?J{)?�Ň=f�[=]~���V/�8]>d��>�^1?���>t��>.P>Ͱ	��ֿ(Q)��K�7�O��Q�r��<��N�w�w�^���i;�I�뽂�<"l>7[�>,�v>�FJ>�,.>�S>a��>v�S>?5�=ױ�=O	������1���e�<`|t�3
������"��<݃]���½"������]���7����`��?W`5?�u�<_.r�M���p��?����8?O{?e?{�B?��=�<��}N�I0(�<˽̠?䭋?�0?R�1�"=��B���=��c�>�׿>j�>>��=�}">����Kq= �z>-+�>�՘>�H�2�Z�uP��n�Z��>�t;�`���[�?"H?��Ҿ�m����.�HA2�H`���@�Y�l<�`��:����"��BJ����hS���B��M��C��>��?�~������8��h�h��[޾��`��=�	?$��>Tu:ޡ\��z��-�f�j�(��P=8��=�LD=w��>F=A?�5?��`?�S�>}_>�7��6_?E$�=Iپ=$��>IK?qA?�?��>�"�>��>f��=$6� (R���<������>9�q�ō�=l�=m�ѽҿ>������j1>^u���s=�&>C����E>M.>�F�=��?H?�-D�,�=9Ͼ���?ֈ=���2���^=�lh�ؐe=6�Z>�Л>b�^?D�^>��3���w�V� �=�)?�.R?��?��=�(��a(���'�iǎ��=~�m��<��޹�S���ƥ>��>�ܡ=�$b>��}?}B?�!?א���"/�$�w���*���ü9���r�>���>�I�=&�ݾ�7���r�T1a�G1��eS�A C���	=���=��>�>>=а=��>�&(=L��M�ս��Z<2*��a�>���>�t?�%[>�=�ĩ�� �~�I?�נ�M�����EDо���+�>J�<>���/�?�
���}��⥿i=��)�>���?���?1;d?�B�t�I\>-�U>��>'�7<:=�Z��⧃�ٺ4>���=L�x�	H����;t\>�|x>�Ƚ�ʾ�9�kbC���ǿ�	h�P!����׾�P�[r���:�j6����ξ��ƾs޾�T�������aXA��b��૾�����=���M�?�N�?���>K�(����՚,���6�3c�=����0վ3.���.����%�����8���q�� W�2+g����>]�S�>o��rC}�~�'�;߼�D1>�w.?%Fɾ�C��^���t=�+>�<�+�jc��SA������T?	�:?e��������
>D\?�1�>M+>d�������>;^1?�%+?0���͍���������?�}�?�W@?��O���A�f��Bg���?�?-��>;c��{�ʾ�n�Q?��8?4�>�9�o����"�>�Z?F�O�a�a>3��>�ՙ>^a�����1��r��)d��o�7>�	�#��,7d��NA�'�=A�>Now>�]�{I���S�>����U�^�)�X�=��JZ��ؽ<f� ?�g��f�=��>h}=ʴ �C���\���ٔ!��1?��?x�*?��C?m���с�Q���㻽��>y\�>��n>�"~�1�>��>\T�e�|���W�>��?���?n�a?�9e��Nֿ�K��V�̾2/ھh�>z]<�c��=��H�V޵=�5�>�>�P�=f��=�"P>D�>��>EIJ>A">��?>����S�!��$������
L�R��ʦ�Y������׶)�O����X��۾x�פ!�,�����s/�EVV;P�$���=��>ߪ�>[ �>�\S>sf�>Iu� b�������(���"0��	��پ��߾R��Gn���l��Wu�AK���B�d�!?\��>��8>Q��>|��>�����>�On=g ,=v�a>O	>�Ӓ>�d�>;�>
�ҽ��>&	>5�>��5>}�����G�l�z�P��Y>���?���'[=�?Ï����6'���,N>u��>72>��5v���щ���>��	�'OH�����1V�SO�>'�?$�d=�Y���\�=�l�kՌ�g�(=A�>u�;���=�������3=O��>}N]�A�l>C��>�<?�*x?�G�>�j<�{	?�#s�\��ClL>�F��%�>!�>��?x%?�P�>��?Y5�=|�5ࣽcP��w�߽�j��uٽ{�伷�+�F����=�Y�=(>q�>0�ǽ�a�w�y���'�6�>����>��M?$?��>L~�UP�R�-�H��I�	��#��JAV>�I�>�;+?�K�>��><[�=W�j���J�6v���>�˙>� p�>x�K�ƽ� >"o�>�AJ?�]�>��k��4�3�+���T��0�>́�=�5?�!?f��>P&�=5
�u[ۿ�7�kJ�r��<�[\�L���<����>5:�=i����]>��E�q�ս��E>ʬ�ً=�_�># �>���>v�>`�=[
�=qC\�k'>=�����B=b�=o�˽�"�=E�>��;�u+=j7�=9o��r��� �K^�BE?�a3?�O�=�����-�g���ɽ³�>C��=%��>=2�>���bA���:���.��<x ?صm?�f�>]$����u`���Xq=�?��?-�>G�>,�>w:��A���!�>od�>٬�=�� �e�^���c�}K9�u!�>r<$=�9��Vȕ?�ZS?x�򾩩��7�%���>�������;��]��<���S���p徊*�
|(��cz�"�ѽ���>L�?������=U�.�����~�n�����c�٭�=i�>���>��=j@���I̾�f��@6�]�
>��>��4>|�G=T>�>��$?�	d?��U?bȺ>N����4?��&���>�?�w�=,�8?�Χ>r����b=ⅾ�>����_e����C�;���4�D��=��R>�:мU�,>	Ԫ=��==ھ<_\���Ǫ�Z}�<�q=�T�;�>��5>��?4I+?C��=$N>:w����m�˄<n��=���=�<Ž�G�������>�n�>�d(?F�
?��{=���'��������>��?�S/?��!?�%���=2۾��g�q�|���]>�*=�B���UP��ɠ��ܾ�3�>B�Q>�=W>�dX>�|?�I?E�?v���?��Oz��i(�R�9D���>G�>%�U>���[+���p���i�,�A��y-��(1����=���=n!>�fl>(�=g�>��K=�Ni�� ��R�=\)=��q>�	�>2��>#<�=hZ�=-������Z?g��+�R��M:��+���?�>�e�>�澩�?��>P��h����a���=IF�?��?��<?���3u�e�>�D�>d��>jR�;a5|�^e"�.�9�F�>��>J�ɾ�֩�kPn>h��آ�>b��<b���w��9��=벿�b��g���̾�q��lU�����Ń��vG�qq�=b��jj�����윽�M�=V�=�K����k���������?$�?;׷>��ܻ` �	�?�D�^ͅ�����櫾<��Z�׽��#<����R����;'�BQ���W�^,�>r~K��ґ�(�}�|*�1���J4>H�/?[ʾ�ִ��D��`=`y >N��<R��=0�����>��~Q?��<?8�뾁���G��H��=5�?VV�>vE>�J��V�ݽ�;�>��*?!+?!���I��ػ��t��P�?E�?(@9?(]Z���=�Ҿ����v�?K�?I\�>���W�ܾ6�����?P�,?9�>�'�	���Z�"�[��>�AV?��>�â2>F�>+am>(����=����ǼJta�hd��=�+>�z���
��N7�E�NI�= �>��U>=��ܕ�EF�>�쾹cS�yR�"ž�S���K�� �>��ľP��=�Ww>/�Y>4*2�����+�l�E�E?��?>jK?�<?���/��aS��4�=>6�>�`�>G/�=�U��>���>��������K��n?P}�?'(�?��<?Lr{�t=ӿF���¶���6�=Sr�=�>>9?߽S$�=��K=�֘���:��>y��>ƹn>	x>�T>9�<>m+/>+����#�@Τ�ߒ��OB���ɠ��`g�9�	��y�X��L������������f��._G����?�.�����q>Z�>�P�>1N�>�|+>�y�>��� ���EX�6}����cO�� 2Ӿ�"�_���X1=+5��Xx�H��2�O��>�u���>j�>��<�����>�ѐ����=��=���=a�>�^=��s>&>�e0>opW=B.?%33>q���A���퀿"���0�>��?��8�X�P�MD��c�T͖=�^ѽf��>�$?8�?�����צ��HT�>�5C�4۹�!"��,� ~C>V��>�N�/ȼ��>�}̾��ȼ��=fq=�l�>��޽Ќ���ϼ^z,>(��>�O��W��W��?�R?�	�?^��>����zl�>�}T��=.<��>A��=X��>����;9�>�?��>�>�@=����f�1�n='��mk<�>k�v м���3a�'5\��'4=�-K>;%>~W<�<߻�k��>�<��J����>��F?���>{�?N���MT�@;���a����<�ͼ��0>�s>�?��>�c�>�,�>�4:�P�l�Q_ȾE�>3��>d�o�G^w�e����Z=c#�>�y]?G:?�c�>��ɽ����H�L�5>���>��(?�N�>���>��m>\�
l߿~
��)�rU���i�O�Ev9�j�>���=Ak���(����⽛��>�A*>:l�=!�\>��q>�X>���>���=�֠9Er�=��i���>?Gֽlꇼ_z=���=[���ub��׷�����=���<�1>�[r<�b<!�= �>��8?��>!�ټ��1���7�l ��?(>� ?�n(?B��>��=�<8��!��Nl����F?�ц?DDC?u�r�[�;�ϼ\
=�w�>)�|>�8>]G+=��1�T��"И>�l7?DȦ>Ʀ>[���";���XI߾�>!����i��?'�\?
7��/���?5��L1�`z���?�O�нd����:��c�t�6��Q¾�2��
���#���-??����ü;���.����o���˽��+�>cg�>z�@>��T=U腾��Ҿ��B�B�7��S�{��=���=�R$>��>-&�>Wf\?a�?*��>�-s����>L޼)8h>�?l��>���>��d>E��;���>�H�~A�=�n�������_�(m��y��=�;>;C�=kj��>:�=ˎ<���ob��h(�=������5�+g=�%��d>Z�=΄?k?c>��>�a��VF��y�=���==�,���󼶨��<[��=�>�>�	^?�Y�>e���-/�����(81��ݕ>/?�?$�#?��q=��;�B����=:e�=3>�8x�-Ӿ�|��M)����8ϯ>��>?{T>�A>Kӄ?��U?��(?9�߽��;���W�p!�}r�<�>??4�>Ώ���ʾ��������)�?g߾md8>��b��V���>G�O>��k>XC&>�j">��<C��M釾� �d�>�LP>�~�>���>slN>~�">5���`�w0Q?�<��
R�ᐶ��u�[ג�̎Y>JZ>)M@���
?i��M�{�Û�k�H�wE�>~��?���?�W?-�j���ˡH>?Id>�^>���;�y�̽T�����<>�Z�=��ɽ}�iSi=Y�>�e>����Ҿ�|��s��ÿ�sS��j�@(���]��g�{��ž���S�������&y���ݒ�'ۈ��w����ß߾�~����ϩ?��?_Ԣ>�o�<�Zf��/��4��:> ��A��lBb�l�A�7f�%������ �;�_�>#b���+�{ʛ>��Y��?��!�|���(�� ���?>5/?�hƾh˴����b�g=<w%>�c�<�7﾿������"��SW?a�9?YQ�D'���"�`�>��?gq�>��%>3)��� �>d34?S�-?f�켂��06�����i�?���?4?�䞾��G��ᾪQ�==`?2��>�K�>�w]�*�־�{�qI.?$??#?����(v�,��U�>�:9?k�`���n>V��>���>	Rɽ�o����=�o��m���P�=�!<H�C�=o\�Q.���v=K�]>�H> Ψ�(���S�>����U�^�)�X�=��JZ��ؽ<f� ?�g��f�=��>h}=ʴ �C���\���ٔ!��1?��?x�*?��C?m���с�Q���㻽��>y\�>��n>�"~�1�>��>\T�e�|���W�>��?���?n�a?�9e��Nֿ�K��V�̾2/ھh�>z]<�c��=��H�V޵=�5�>�>�P�=f��=�"P>D�>��>EIJ>A">��?>����S�!��$������
L�R��ʦ�Y������׶)�O����X��۾x�פ!�,�����s/�EVV;P�$���=��>ߪ�>[ �>�\S>sf�>Iu� b�������(���"0��	��پ��߾R��Gn���l��Wu�AK���B�d�!?\��>��8>Q��>|��>�����>�On=g ,=v�a>O	>�Ӓ>�d�>;�>
�ҽ��>&	>5�>��5>}�����G�l�z�P��Y>���?���'[=�?Ï����6'���,N>u��>72>��5v���щ���>��	�'OH�����1V�SO�>'�?$�d=�Y���\�=�l�kՌ�g�(=A�>u�;���=�������3=O��>}N]�A�l>C��>�<?�*x?�G�>�j<�{	?�#s�\��ClL>�F��%�>!�>��?x%?�P�>��?Y5�=|�5ࣽcP��w�߽�j��uٽ{�伷�+�F����=�Y�=(>q�>0�ǽ�a�w�y���'�6�>����>��M?$?��>L~�UP�R�-�H��I�	��#��JAV>�I�>�;+?�K�>��><[�=W�j���J�6v���>�˙>� p�>x�K�ƽ� >"o�>�AJ?�]�>��k��4�3�+���T��0�>́�=�5?�!?f��>P&�=5
�u[ۿ�7�kJ�r��<�[\�L���<����>5:�=i����]>��E�q�ս��E>ʬ�ً=�_�># �>���>v�>`�=[
�=qC\�k'>=�����B=b�=o�˽�"�=E�>��;�u+=j7�=9o��r��� �K^�BE?�a3?�O�=�����-�g���ɽ³�>C��=%��>=2�>���bA���:���.��<x ?صm?�f�>]$����u`���Xq=�?��?-�>G�>,�>w:��A���!�>od�>٬�=�� �e�^���c�}K9�u!�>r<$=�9��Vȕ?�ZS?x�򾩩��7�%���>�������;��]��<���S���p徊*�
|(��cz�"�ѽ���>L�?������=U�.�����~�n�����c�٭�=i�>���>��=j@���I̾�f��@6�]�
>��>��4>|�G=T>�>��$?�	d?��U?bȺ>N����4?��&���>�?�w�=,�8?�Χ>r����b=ⅾ�>����_e����C�;���4�D��=��R>�:мU�,>	Ԫ=��==ھ<_\���Ǫ�Z}�<�q=�T�;�>��5>��?4I+?C��=$N>:w����m�˄<n��=���=�<Ž�G�������>�n�>�d(?F�
?��{=���'��������>��?�S/?��!?�%���=2۾��g�q�|���]>�*=�B���UP��ɠ��ܾ�3�>B�Q>�=W>�dX>�|?�I?E�?v���?��Oz��i(�R�9D���>G�>%�U>���[+���p���i�,�A��y-��(1����=���=n!>�fl>(�=g�>��K=�Ni�� ��R�=\)=��q>�	�>2��>#<�=hZ�=-������Z?g��+�R��M:��+���?�>�e�>�澩�?��>P��h����a���=IF�?��?��<?���3u�e�>�D�>d��>jR�;a5|�^e"�.�9�F�>��>J�ɾ�֩�kPn>h��آ�>b��<b���w��9��=벿�b��g���̾�q��lU�����Ń��vG�qq�=b��jj�����윽�M�=V�=�K����k���������?$�?;׷>��ܻ` �	�?�D�^ͅ�����櫾<��Z�׽��#<����R����;'�BQ���W�^,�>r~K��ґ�(�}�|*�1���J4>H�/?[ʾ�ִ��D��`=`y >N��<R��=0�����>��~Q?��<?8�뾁���G��H��=5�?VV�>vE>�J��V�ݽ�;�>��*?!+?!���I��ػ��t��P�?E�?(@9?(]Z���=�Ҿ����v�?K�?I\�>���W�ܾ6�����?P�,?9�>�'�	���Z�"�[��>�AV?��>�â2>F�>+am>(����=����ǼJta�hd��=�+>�z���
��N7�E�NI�= �>��U>=��ܕ���=t����P���y�GF���R�a뇽���>4p*��>�2/>.�>���N���Lt���_���r?�Y�?K,H?AiC?���[�ھ0�=;�#=/��>��>�żA�Rig>��~>+&���L�n/�'z�>#��?S��?]�F?0g~�g�z���q���3��)
�=(��<^�>��J�l��:$����A�/I$�1�>�T�>W!W>��D>p��>�9>Z�>}��f�"��I������A�A�+L�����{��G	��l�M���������������Z=�$����A"�%�?��1=��9ϼ}|�>\��>��h>�=�=���>�2�=c-���۾��
��D�����W������j���D��7�>�/h1�����n<��J2?7�½�K�=2q ?��U�?�>���>�������>~�7;7ZV>��>�Ο>U�[>��a>䜬>�iC>YR|>N�=m��
|�u�;�X^��#�<�oD?Ϟt��{��47��Bܾ�c���v>l` ?��7>l�(�NД�� t�s �>�[O��q��-ҽ�c6�j�>���>���=�����@�%�q�c��=���>��>p|�������9����=\��>dTо�G�=}V ?��U?zR�?�b?���W`�>3&?���>v��;���a>��7?���>L$?�
V?j��=<>p=�Z��O��&V<�{ �Ro�=Zaq;�:f=
�;y=Fa��X��=Rͧ�Z�'=��=�*E�۲��l�?=�F >�?'�c?�"?�/�>�W���r;���c����5�`>�i��A��>A�?�?O@*?���>�@�>)��=��	�i$'�ݺQ>�i
>����z[�X�.=��>R%�>A�M?}"G?�E�@wp�"B�W1�;�>���>�;?�|�>S`>hJ@��$� �̿F�{0��k�G�U钾�SC�aFS��UJ>�e<������Q=t�4><�N>9�>
qW>��>��>-d�>yD*>&li<�N۽L�n��^�=m0+>��=$D�=�mP=���=i�:��eRr�н���A���.=x�=�~?;�
?P�6�<��=����V�7'f���>�Ax>u]�>��>q8��	���d�+^��Ş�C�>�C2?s?|���P��=�'<|s��0��>�s�>�U�>W��G۾(��|?O�k�>�V?z�g>MW6��"A��xT��$�=�>>Z���g�?ۚ(?~I	�dYw��M�dF��s�:��cϽ��¼W���2�q�,�oaD�z���1��c��kؓ>��>*�?�>�S���4�R.��1~��%]��a�=�>�	?��>�<�������Z��0������!�Ӕ�=\�=0|>͚�>n�?	�?+�R?�?1���h�>�8Z>�?[�?��^>zV?"F?}�?m�=���>Y��e-9���{�V_x��>�=0��<��ϼ�H>Λ:��m���N��&i����\���=�z^=��<(��=v��=�#�=�
?�jI?v�8>�����+���1���C�p�D>�m�>��.��+�t�>��>�3�>�0 ?�0?��c>(|�C�"���ܾ���="��>և?9K ?�>H9>	�羭/ �y.�>��Y>*���
���0���Ӕ����#�C>��>*)�=wM�>���?��E?�^�>�5�	A�Ģ�����0%O��:���>�>�ƶ>\a���/�dJC��W�o�3��#�K=M����=��A>YN+>�ǔ<����=	�\�
n
>����e��=�0�>��
?��6?�Z�>��p>�1˾-�2�Q�G?�a��-)��Q��'hž�*ʼ��#>jn1>Q� �%�?���[�������];�|��>
e�?���?��d?�0J����M>>gS>�>�L��40O�r��j�7�Wn4>-��=a	}�=���,���
R>w�>�a۽|���Lv۾��7�5]���5.��� �z��"a��Ϙ����I�I��,��@�=ɸ=�L���� ��Ӿ��<��ћ��׼=~�¾-Pо��?�j}?`~^<I��>gp�%�8=׾�P.>�_5��� �+i���C��߂�k�b�����ēE�9�i��N�����K�>�'��۵�ɉ1�p�^�tV���=��F?���$-�� �8 #=���;-;��(�r���#똿W�߾�Y?M?�򳾕e��>N�>A �>8,�>�q�>m����)��m�>Ȥ%?��?pX��(���c�H�&�.n�?��?��<?rSw�~$T�|�^��� �f>�m?�1?V&¾~���O�+�_!�>OP?X��=�E�ʿ���7��^�>�_�?�ㅾ�Q?>��?�d2>4�ԼVоDz������Up�n��=���"v�f8���8���>�ٲ>#MZ>Zb�c��-%?�!A��i�$3~��hE�M��e6M>ț!?�0��6�>�G$=�P�����x��Y��Y伾? ��?2eE?�?����[d�#�f=��;�9j>^��>�E>]������=t�> �k����s����.?���?`��?�O?����מ�y��7�j�c�B[>:
3>��V>Z��)&>�a=���<����>�.�>�}>��h>�a>�>��G>y(���a�	����7U`�G�?��*�;�U�:�"�vX��\��"!��o=־��#�~����d�)㐾�.��ձ��B ��0#ܽ�с>���>N�>�;�=2�>�*���������4��a-�E�q� �����[��1=��D�<�N��#�<Y#�lV?����uL>�j?PW����4>w?_>�����>H��>nO>9θ>�G�>��>f>�O>p�=�{>﷊= �����z�9�X�P���;}�C?��Z����O�3�bH߾>q���I�>��?�yU>�''�����y�*}�>�GI��pb��nͽ%j�߉>�F�>�~�=X����j��x�W��S�=�ބ>��
>��k�A	���'�x{�=���>ټ�ڛ>��j>�1$?�x?�	7?|Ư=�l�>��1>��t>�	�=�5>��<>b��>��?�<?��3?�A�>ɩ�=�?��2=)�=&=�C[2�{罉o��q���?����O��i/=�:�<�
=7�=�M=���N��:rs*=i��>%�U?iU�> ��>T �:L�N�f�j�n���>�F���>k��>f�?�&?�?�Z�>\(O=���q�F���>#�8>�;��Hl�W�> ѳ>D�R=�G�?3Ls?�� >vT���l�p�߼n�`>L�?�=??�ż>l�v>�������fӿ�$�s�!�{���0�К�;��<��hM���ٸd�-�.������<��\>_ �>��p>�E>|�>�D3>~Q�>P=G>G= �=3�;;|
F�aNM=���t�D<�>Q�)l��yCƼ�ʗ��"��]�I�O�>��P�x�׼��?�
?�۽�R������o���u�<�>�c�>!I�>��>��<�g��e��+K�YpN����>R�c?Nr�>�~]�&�3>��!�1�=s�>�v�>0_:>���C��๜�����λ>��?��>���&T���v�p�/�>!L>�/B�*��?�>X?���{�$��D!�?8��i��k�C}��t����.����٭0�����ǾN��<���>-��>���?"̾\U>�����\��}̚��ܾ>�|>�>V<?��>�(w�����Ĥ������7�½;�>�Q־� �>;?.E�>�i?NN?!�>���<�4?�����>A��>�EG?L�'?�a*?��?�?'�N���`�����Tf��=�=C5&>NE�=�<�=V2n>dKX�Y�I���ގe�uܜ��鯻�(<ĥ�2W޽`��=�R�<O��>d+?و+?��ڽR��9"=�������
�>2Q�>ߦ��[�V���P��.S>�?�o??4
?M��=��þ�=
��t����9=�?�?��>���=��R>+���烾?m�= x->�v�<�C$�����������7�N>!J�>�\T>���>"4l?��?51?��~�Bg.���w���^���Xi�$?��+?��K�<��9;�u@���l��y1�4k���\�>���=�=~��=!��=�B�>��;hD9����b=�ҋ='�?;�?�.?`M�>u�K>����!=�j@?�Ӿ0&��c��y���K���p>|u�>�e�k^?D�<���x�봥�̷[���z>4�?+�?�4h?�`#�~D�L��>A�|>�v�>~O'>NM�5sj=�;4����=�����ž�B��x��[DH>z�M>{�ȼ4YʾfR�-xZ<Ϭ����L��h�N׾�����پ�j¾��s��g��yܼ黾D����Ÿ��A"�ֵ������:3ܾr�w�bx?�R=?kp̽e�h��`��7.��h���i=0Ծz"*� ����l��1�v��+�AR�8����=�-��ľ�ڏ>��˾1꛿����fv?�؈7��>ǉ?9��/D��2	���V�K\>zE���&�N�������#�}���u?1�i?���/�0�����!����>���>Q.>/���؀��B>p?�d,?��������؆��+��U��?�ٮ?��??��O�ңA��{�H!?�?k��>(֊���̾aF�?/�9?>>"�e���2���>ɗ[?�AN���b>c��><L�>𽺪���0&��;�������9>���Z��,Sh��>�Q(�=��>��x>_9]����u`?�������^'x�-:9�+"���=��!?�[
�B(?�@?-�þ��9�w��V��+���b0?���?�G?J�?�@���n��5��h�ƽz������>P>,�����>��?%����8��~���?b��?�6�?&R0?�x�@ տ�դ�و��W뾢�>��7>[>+5��f�=��<a��i{�e�<>Ol�>���>(�a>���=q�*>��%>[���O/�:L������kd>�K��3L�
W���,�m����6	���������c�<�n7�����m����6���J������>���>��><j�>��.>D`P>z~V��3���6��������|L����8�۾�<��h/�}�5�t���$������~t	?�$мw��=���>����d>�\�>6�$=՛=>[6>��6>�C>Hb6>i�Y>9+/>��U>~߰=��{>sH�=*��m��{n:��Q��;�C?��]�X����3��q߾����Q�>Ԗ?��S>!�'� ���t�x����>A-G�&�b�{�˽f/ ��^�>B��>���=��Ȼ�b�νw��U�(�=���>Z">ۗk���9����=�>�̾��>M�->y3?<�x?J�I?��=�@�>��>���>Uq>��A>�7c>[��>��?�77?5�%?6�>�"�=|4�I�=�J�=�d	����<ʌ��$��y꡽Ғ���܀=;�J>�g�=�c+<�MY=3o�Z;��k��	<���>�IW?G_�>���>p�½��@�0�>�֣A���>|Zk���?n��>͂?�+?v�?fC�>hǼ�y ���*�h�>oTb>F@�G�}��d�=S!�>�a>ɶX?��h?��=�Ǟ�X[X��5
���$>s�?CK?60�>�7>Pe7�sW�\z�l�.�Q�j�����Y>_v?>����� <�v2�m��fؤ<� >DG>���>�&�>�WB>��>@��>���>ߢ>�=a��GX��m�<�o��X&�<\��;�E*>��q=C`>s����>��L�յ��IK =�w>�E�P���?��>�胾/"�=!�_���WG�D�)?��>��#?O�>��콯�3�5�^���H��Ǌ�q��>%�e?�/�>��l�;(>��Z<No�=t,?g��>�=��0�ʾ\�	�Ջ�&�>q�?���>wD����p�$m����S>%����;���T�?��j?i�6�!���j7�\Lg��G��0~<�)
��ξ=7"�'L�\�H�x�J���`��>==�"?���?*���_>"���4늿�hi�v�R�]H�=�=��?
��=h~��uU��h|R��̾t�p�Gbz�9z?CP��ξ�>�:"?7�>9�?)�D?��3?�{۽�C"?���'@>�?��)?�*?:&?b�>[�>����>�[��T����=Y����zf����=�rS>�'=���=�9�<v�5�obн�K��kP�1;<�2�=�`=`�=Yt
>�q�> LE?�ܽ����]>ͪ;�Zw�K j>�=�>��;�	��4y=^�J>���>�9=?+x*?�g>����y��v��ڌ�<�z�>�&"? �?�2�=�c�=�a۾�)L�⳦�B�9?�=A���[߾mѾ}�_��AZ>,��>pn�>I��>?��?;\?j�?y�n���3�ޙ��S3��Ʊ��T�՟�>!h?x�>ۆ��V�Q�-^���*�+ܾ�NV��5>���=4>�U>s��ώw>Gtn��{ټ��<��=��>�"?�?�W?Ce�>��k>����m��5T?Z�����(�57��}���*f���>��>K�����(?��{=^d�����	�P��_>�{�?2$�?L�r?3W���7����>��>>�>9�B>;�����&�<m�4>�e���ž+r彔'+�oʳ=4��>_/���e����ȟ��V��F�K��k=c��uM���͵�V3��m-׾2�����v�e'�������5᩾g�<X'�,3��������>���?;b�?e��>�Kr>YCe�-����͍��־�[�ʄ ��$׾TC޾�;پ�X�!pD��$l�#WK�eA�p��>�,O��?��a�B��G�
ne�h��=��(?)��Op�~��3J��n齦
��!�'�h^�����r��Gf�?q^?�K ��F�% �%�=�0?7{�>*��>�����=���>FY�>&D?r><����$i�ɖ2=T��?樞?)h>?;Le��rI�_ ��i�3�"�>�?\?*	���	v��	����>��?���>�8�.�R���?�C?�$9��h,>�4?J:>��T��x��x�/K��D(x�=��=Q�u=��*�v ���^�G�=ʹ>&�p>0�B��%��I9�>��x�Y�^I���
�K+>�U��;�9?�I;G>�Vq>���=�#��/��]�����0�8�8?�"�?|tb?�B,?���ھ�+ؼ��^=݊>�P�>�z\=~�?�>ݥ�>h־-;y��&�ڥ?ǻ�?�n�?7R?�m��Gݿ?������N㾬? >�2�=��y>�i��Q�=�j�= �<��d=�<w��>���>VPK>!�4>�X>�=�=F��U�%�Q)��<��@�]�����*�����������Sܾ�q��̾Ʊ���8 ��=���Hjt�r�n��!��{7>�?[t�>Ϟ�>��>>��7>˼v�q� �'4u����O�x����\��Ҿ9(~��4�j�\�����D:��o����?�U<��>r��>�:�O�
>��>�Ђ=,,>�K>��>&gS>�XN>�IY>jQ4>!	X>���=��{>��=&+�����ty:��Q�aQ�;]�C?��]��a��N�3�^�߾u���v�>�q?�aS>��'������x����>WH���b��̽���v�>j��>sA�=b������Q�w�y�M��=���>�_>��e�㏾�K�,��=�L�>f1���f>�D�>�:?ak?p�>?A`�=� �>��>�ޑ>I]�=�$�=&,>E��>h�?E�;?��'?��>o͛=ԍ(�7�=!��<L�0��A������� ����̻ļP��#�=aN>L|=��=
:�<�'޽�$D�8��<�	?l�Y?#��>�>Aì�m��d4a��+��,�'���>l�?� �>��>?�9?�?LV>>w:�쨓���4����>�}^>~d.�̀(��V�=��>��->�??��G?��������j�5�3Y-����>Ci"?i|l?��? ;�jE�Q5
�py޿�*��!�5�,]��Z�W����=@�3�aJ=��5��rn���r�rF��P�=*�6>)�9>�H>��@>{t�=���>�q�>��=�(>=����"����ѶJ��Δ����>}9�=j�8>��e>�R,�����������b�<��><�?�/?X?u��S?��@�����-7E���>��>Y�?��>��q=����v��d�Q���9y>�(g?�?s�����=K�a=*E=s �>��>�Q�>��o�<B��Z4	��ǉ�ň�>C� ?&g�>_^����Y��Fy�n���|>��|=Դ���?��D?�C���ݾnM	���4�?�Zڽ����ܾt뢾�.���5�SVJ��j+�����Y>S�>�.�?7��^v�4͵��X`����z�����H��8>�>����I��@|K���:�w�M/����|4=@Ϧ���>��>��?��?}�?y�?f� �6?/�ɾ�U�>���>~?v;.��>�w?Ց?��?@�G>�ҽhȽ���w�=
�@����<�^>v�>[��<Q��ӿ�^ڱ��⽭v:�P�H=���󎽁:ҽVA�=)K >�9?bfI?G�4x>4:T=TE����	�뽀��>r">=ڳ�q�>��S>�0(?>??^,?'r�>�1徼�!�����~�<�d�>�f<?4*?�-��>9�ت=("�=~��=�2=�i���a������1���
�>*�>��k<0��>��z?;7D?*�?��[��&�	D~�0�.�g�!��@r����> Ժ>��|>$�޾�0��t��sg��c�`_I��B��	�=�v�=ؿ�=��/>|4r<F�J�h��݄��T߻�=���<S��>��>�O"?���>��[>����0G-�uYD?���9��:ƾC���Cd�=x/�<Pp�>o@<U�?��C=-\���u|H���>�$�?95�?��P?��t�ո����_>I��=҆"=術>�;�)5�����n8�>�2�=���t8�+�=p�=x:�=�"�<��G�gK��6�b=>���[�9�I��=���������bA��qξܗ̾Ƥx�)��=�����:������z���Ƚ��8�o�O������B�?7R�?�$�>ӑ>�j|����d��
���ȾO�W��+A�Wh�c����Yؾ"Ƀ�����r	��)�8��C?o~T������g��:cM�<#>���)?��
�n�:>^U�K.���	a>��@��C��M���y��,����S!?�uc?�(�N�X�񸵾�t�>�t'?=E�>�^?dy�9_>��?��7?A�.?S\&�8 w�۠(�{���tx�?���?�UK?PҾteD��M��*���X�>/�$?"d?���E�V�ž��>H�?m����h�ꎿ�=f��A?�L�?��9�rȠ=ƿ&?�'�>�}|�P�4�fD��K��Y��`l7����=N�q,M��M	��*�>Oc�>���>)��,0=�3�??9�2�d��S:�'w7��5q�ά�>~�-?����6�>·�>�H��/��$���aش�c$'?�z�?c@R?�?f���U��<̍������>EO
?Kq^=�F>c�>G�>��]�
T�����)?���?���?�A?6�i�P�Ϳ-���=&��H���e*>@�>�k�=����2>`��=�	�=]�����l>��V>�\\>��>
�o>��>�A>��������Q���H�*�Ц�v�:�����f�G7C�0-߾P�Ͼ�����_���ž �y=����]ýC���ap��~p=oQ�>1�>"{�>��)>A�>�������R��yIʾ��,���]���Vھ��6��ܳ�W��^�D�_���֧���f?���İ�=��?��^�'f�G�L>Y��+Ѣ=�z�>�=�>r�>�l>߇9>\r$>�E>�>��o>��=l5���@��j�8��
H����:B3A?��U�L�����4��߾�����]�>G�?��X>�#�{t���x��j�>��Q���]��T��c2�R7�>�Z�>YN�=H�u�o�d`}���ݽ��=���>�b>0���풾�H�ˌ�=벭>���0p�= g>�K?<�i?е2?s�>��h>��=r�=h�ֻDs�=�
>]_Y>O6?D�5?�?=?��>���=��w��p�=�H%=�sS��<#oK�cF+�D�pF���ڽ�\)>��E>�n==+�1;�ȼ�{�?�|�x0H<�a�>�>=?T"�>��>6+D���=��N���"��>D(M���>��>�O	?k?2G�>�>�P���Ǿ��ڽ>��*>�l^��p�*٬�0}�>�@�>�rG?k)?�0Ľ�5���`�<=��=y�>�?L�#?�J�>�#>�½�����<��&Zu�����8�="�>��ݽӠ��N�>���]�̾�����#l�6`���A��&?��,?�y�>�"�=S�>uKB>O�;>�>c�)��y���f�<3/i��K2�\%���8�kq����c�R����,;<����̼	!�;����ʣ?���>G����<��G��}����?1�{>�
�>�:�>C�R��p%��L�B�;���;�P��>��k?N	�>�I���RK>0�I�h^ֽ!��>���>�2>
9�=��Ⱦ\[��n]=���>��?�T�>�nY�3Bh��n���PFj>�B>��½�؃?\�L?�t&��f�h6��T���6���U���D��'��徠��6�6�i�"�)�)���ʾon4<�D?eL�?YR[�q�p>o���I��hTV��|��#>A>�>ȱ1?p1o>�Ӿ����D�B������N=�!?&>v�$?N�5?�Y?��q?�6�>��>�_��q?U�<,�M>,�D?�)h?y�Y?L�a?� >��=gԼ�`�L����e�o���h�q��>q>��G>�->��v=֙.>��=����ƛ�7����ٖ��
����=9��=��I=?G>�?d'%?�[��),�cm�5��N��<S��=4m@>�ꋽ(w]��o�<�Od>;3?��0?���>�9=X6޾���w5 ����=�?//?)�>L�B<c�=G���E���r=C&H>6�B�p �����R����뽪��>���>�P�=��>^�?g<b?�s*?����aI�}��l$�I^	���=�OC?'�?L>>��;G�����I��ml�<�1�>�0�T\�m[�=��K=��&>��D>�K�=DE">(8m�����7\ؽ�@0<�9>�'�>�	?�!;?L�E>��>l���A��߄[?I��B^�*�#��������>���>���-�J?���j9���У�P�A�S��>�7�?���?�<w?�0����Q����>s�>(_�>���>�%�Ck/����>�=(E<y���7+���&�*��>�	�>my��q+�߄����7���I�!���
���վ
�.��P9� ��ey���Lξ����Q��p�e������?���Si��A���q#�%�?�)�?�&�>�q�>l*R�����1��C�=���O
��R��)��.�^��ь�\��7%�ZD��5p�N�%�+��>�?��Y��L26�.�I�֗��"�=��D?C��������,̽SJ��@�?�|&�������ذw���?]g]?�p'�)�8��˾I�$>+1�>�?��?c1ľѪĽ�Պ>|W�>��??\��'���&����ɽ��?*&�?��??�yU���>�p����?��?E,�>=����ξhb��J�?k�6?R(�>��~�����;B�>�[?�L��b>C��>���>����w�4�F��Ә���0>Xj߻��	���a�9k>��Ƙ=˝>�
p>�a�E,��;s?�	���t��,���`����>��!���E?�a����=/=?�>՛|��ȗ���p��>���Z?(�?4MS?��+?"���[��ʞ=����`݀���>��>�L����>;�?"�/��H��a�J�S�'?���?j�	@̓X?R8��
�Կ���J������ݜ�>�>Y7,>�k�O��<��;��"*�C�K:�{>u��>�x>\�p>l,�>7�>��>yb���#�7u��N���(h<�>��^��+��hQ��?��A���{��xѾힽ�nĽ����u�L����1�V<G}���>+��>���>��>��=��>�u����:������������O����m���뽖ʽǗ�[M�����<p�ۘ�>��$=4I�<tu�>X�,�>2��>�)�=H�>y�t> -�>ô�>�@�>;�>��>y�Q>k'�=l>�f�:��Y�u��(��F��6<��>?�%�gv��9�&�ѾK���Ȝ>�?��V>��"�>��̼q�Ř�>���������}��F��$��>���>�a>>?=B��3�����ٿ=�@�>��>�)��0w���- �7��=���>��>�$sU��>�?�X?�PM?�1L>�/?��>/|q�c:�=�8�>>'�>0�>�F?S�?��?���>N�'>���;���;�@>���������#?��潒\��
/N�v�<�ZU=rR�N u��>q<��V���"��u�=g��>3O?`"?�־>�P�F�Z��SO����\��=!�ѽs��>���>41�>?)$?i�?��.=`�@��V�u���ҳ>�)^>�A�v!z�c]�=��>y҈<Mڀ?@�P?x�����z�>�>Q�>D�?}U+?��>�t�>��=�4��ѫ�����w�2�\�='�[��y�����G�_�d�$q+�O�d�#p㼰ǉ>�;f>�)>�n	>W�9=��q>i��>1��=�{��1"">��<siV=I�#>cY=�ܓ�wE>_����<s�B�[U-��� ��O<6vK��,<�X���?{�?yͭ����;g���{���@�>ɲ�>ea�>/ݿ>H��<Q4�(�V���4�����>+;S?�"�>7�r�$��=+��ŵ<� ?~m�>��=�[�Lю���{��=X�?�?�ȣ>��{�g��<b����uUf>V��=�H���?!�`?�K�����D��BTD������<K��٢�E���!jž���5�8�K��ȼ���C��=q��>���?����r,�V/������	�x�6!�gi��<f�=T��>]��=_P��L���/�=���ھ�@s�3>f�c$�>p �=���>$�?
�?��;?�?z��>�&y���?�O<���>��>,��>X?�?���>]��>2j�=��ý{��\����:#>�&Ӽ`��=��{>H�>M^=ܗ0>��&=���<����n�Q=��F��^�:��<Y��=�<>($W>�&?
w?�
��+_=5�]������<�@�=thJ>zgڽ��}���=Ub/>\�>��?%��>Ñ�<�X��"���+7>ø?bV?s��>��4�R�:�@���ef����}��H>�p;����o�\ؾ�9�cD>��O>�m�=��I>W�?P�n?�q?�)B�­@������e�����\�<��\>/�j>��_�"�þ�W^�9H]�LA�ٶ��x��^0�^����&�=g�==�Y->�=WAd>�5�=�Ž1�N=��ƽe�ռ�̲>~��>��>L`=��b�~���0ξz9k?@'�����j;�S��'=$�?:T�>:B=��2e?h9�.�������u��E5?��?��?�M�?�l �{m���Ds>k�>̂�>'�#�ǋ��~X=���� 4C=x%> �!�:�e��HS����>�i>џL��:�\�?��L<Cy��}�Z���n�����@�G���5��
�'��B��B��d�����Ad=��7��E�Ó��`~�L���?�Yw?}k?>W�&�~��������>c=~?3��!3�<I��c.��Y؆�S����˾�~���'�
�$�g���o�>E<ݽ�����}��;�MN >^�=ݣM?� �jؾ|'��5�>�z?�h;�E��}���X��z˽U+�?$lE?����V����h�>-Th?*��>���>�Ћ��d>���>ms!?f�}?R�=HtY��m�
�����?��?�lD?��+�_�T��� �z ���_,?9A�>��?k�=�n�Ͼ|���Q?Id?0��>���f*��r�(�v	?�*�?G��Z�7>���>��K>T����/�˩��3���t��<ƪl>�b�<�2�7<{�ô��в�=�K�>b�>�.T�jV���?�"�@�N�L瑿�ྗ!^>Vj>̃P?���~-<[#??>�=<�!�����#N��w%n��|`?j�?}&g?G�G?4��;F�8�K�:>w�?��>>�>�I�=�:�<�?��⾽�9�[�
�	�?�[�?D��?"��?bPr�HVϿ�Y����1����< E~=��>a����=$��=�.�f�<:�>j��>_� >'p>�>8��=�R>�r���f!�0���=[��T�M��)�����ʪ������ )�h��� �����I�U
m�(o?����T}��̬�=��Ⱦ=�<>~)�>��I>�@k>���=]�=�C�GH���ξ�_޾���6���v��⾕�Y�C��;��N������~�~�?���\���٠>˭���h�=]�=9��=�2�=�a/<���$���\.>�#>yuk=6E:>f�m>�Rr>��=L�������8�k�U�;2�;HB?b�푙��3�lp޾� ���A�>��?��M>�?(�z^��i3x��f�>�A��s^��hʽ�m#�Y��>g��>�S�=������w��i���=S5�><�
>��w�?}����m�=�g ?����ߚ=�>�
\?�Z�? ?	_'>�U#?[&�>.�;>���>|��>sn? ��>y?7P?���>��>u:�>�D���^����=�2н��;���ً��GC=��=R�Ex�>j�=�>G"�<U1���]��4�9�#�=���>x.=?���>\��>D�@���7�$�H�#���̲5>�ȼm�>s4�>���>�O�>?��>�c8>�Pj���̾�侽`�>��P>]�H�*�o��7�y25>)��>�b^?8�1?�J����$����O=0�b>H�?�	?�<�>[>.F�W��&�ҿW&6��s��qf��o���Ȣ���%��~�?��;H�/�IO��*�y=�Ih>?v�>��G>?!>g�>V�>H��>m�8>��=&:�=�+����;jм�f=����F(�፽ �A��[H�ҵƽ����l�)�d]e����4���D�?��?m���y���yg�:g̾�S�F��>˦�>0��>�Y�>�� =�i	��7V���=�>���w�>�c?g��>�_��6}>EF��,���P?2o�>�މ=����*��ox���&>�l?�?Rܯ>ӏu��l�������(����=Q���D�g=��?ǚ$?+��3p�� '�p�P�F�.�o�=y\Z�z�־?�����G<�t��������`>0�>U�?�};���a=��þ,�����2��\����e>��j>��>�.�=M�U���>
(�Ky��(�<��⽈�?�1>"{�>ny1?Ҽ??��m?q��>�؞>Y_�=�?:� >��>��?��>�c?��D?%*I>�e9>U�/���Z���2�����d�= ��~��<�0>ǝ�>�ٿ=u�=ׁ=؇�=��==>�k'>���!�=�@�=vC�=�=��	?�6%?_=W��r�=]�<Ǐ�JȽ�1�=��b>����Z�{�?�=U�->��?062?���>��=�nݾG�o{�<�=#�>�T)?�?�>h��*4>íy�����,�=og>>�FR��-��cT�Wc��0�ǽs�>3�i>�>L=~��>.ۘ?��Q?U��>𭔾˴����;��>"n�>�>;�=��!>�󾃂J��(.��j�W�>��Ͻt�����<� G>{��>vb�=H՘���?>a�G���E�6�#��_>��?zg�=�B�>�0�=,�<��0�;�ɾ�r?��
�����6۾�+�׃	>_$?���>;��??j�=�������o�]R�>Í�?��?��?.Ӂ��ȶ�O�>��>�>ϳI�g��}>w=��˾��Q>5�=�j��<f�\ڲ�4��>��>>��X�3�Mr ���=����gT^��['�2AZ���G��,����#����*���8׽�Ҿ� >��'>G���c��E�¾F��6�׽O�=N?J� ?D<r| >L៾����D���F�=�V�Ғ��<Y���޾�θ���\�D����羌���/H���~#>F������Tˁ�ow5��v.��L,>�-?;/���U��+ �B-�=U�t>i��?�
����!폿5^��caq?*@?5��H� ���s�靭=F&?j�>B�u>�b0��gQ�b��>5??��B?�V=8J|��(t�Gj�<8�?(�?w�??��O�>�A����f�hB?{�?U��>������̾�M�*?��9?ü>~��`��!(���>��[?�N��Rb>���>�8�>��c����,%��
���3����9>*�b���'h�qW>���=#�>+�x>��\�Z����?��$�=~����k�Ӿ�J�>7!�=#&V?�q�����<�?tG�=����z�����/�����{? |�?�|?i�6?�����|廣�?>�ެ>'L>���=��u<�4�=k��>�����v�y�&��k?�n�?�
@sTv?=%��6Oǿ�;����M퟾ȕ>���vD�=w6�޺��[=!���"��]= Ҁ>��+>J��=��7>�;L>��k>�����%������y|��*4�8�*��N	������`���(m� u�^��6����#��ݽ^q2��������־Î�=.��>��T=�Z>�¢>��>��&����<��� ������{�,�nP���k@�J�'����"�U<w� ��8)?7��=(D��ܚ>�:a��o!>X��>.�1>���>�׋=�R>�>���=n��=18>'�]>�>7�m>��=
��w�~�E23�`�K�wn��A,A?Tm�mޣ�q5�iaھ����IKv>r�?�/?>��(�����v��B�>�\/���U��ѽZ"[�Z��>�C�>���=͘^���׼iy��r��Y�=eZh>ܶ�=��Ӽ������z�=���>�Ӯ��?=�N�>3W7?��y?A�<?�g�=$��>���>1�>C[�=�+g>��~>�e�>�� ?�I0?�� ?�H�>r��=�P�~=��)=�O���ý	��6󊽹�սC'���Lƽ��~<�6=3{�>��?��˽rP���=��>=S?>q?�/�>����q\E�I�"�U{�=U�>��	=���>�3?%�(?��@?��@?��>j2�L�� S3�g�>��>:T��6��@<;�>�����>�@�>�%8>�Օ<�&I>�>�@�>%�>�m?�	�>�r���
������⿊�W��H��{�:��l����ZFu��R��j<�,`���:�������Vp> �>C$>.>��p>�M�>��>�>*��=U�?=_hF;m�d>WP� |o=�X>a2�s?�u��=�/�=�	U=ؽ�����=5��<��ɽ.tؽV��>�?��S�X%��%o���ܾ�8�{��>���>���>V��>v�e<�
�FX�I�B����>�>��d?�0�>k��2O]>�e��RMV��?��>�=E�;��Z��h���/�= �?��?Q�>d	��Z!{���l�H���>p���,��\�??�g?��L�-�8R'�g?t�fcӾ�F;N$��ھDv��lI�x�m�F¾����X>�'�4>=
�>j9�?�����K�>�o�΂��h.�kҾ'�R��>Ɓ>��Ƽ�㐽r�,���)��G���p�����?�\�>��?�]&>�U?�]�?R�>��?p��=4 �>�۳>�=&?!?؆?�}2?�?���=�4>b��*�=��(��u��a
q>[�b����=Dx�=m��=&6�=��n='� <4}>��?�
���"齷;���Z��ep<�lL>d�%>�`? �1?�o��ہ<�H�=��8�n��L�&>��>�λ=�T<#�>}�>ޡ+?^V?���>a�����񾁰�i���5ڼn�>��$?( 	?v�Z>b�p>w�T�nx��2?=��>dg�f(Ⱦ���H����:�h�>���>�N�>��>�gX?:�a?�D?<G��.��w����c��)2>�&>.����M>�$>�nU�}�!�J�U�!�f��NC�.�=�� �2�=�z<�׏���>�Ӷ='�^>��)=�W<���Q����2l>���>��?�?��N�O!�ۿ�����]`?���dq!�����)� �*�#4?k?Q7s=�P?i�;�}���X��+^�w��>�#�?�<�?�?�?�<�ǾA+? ��>�W�>T#U�����pt>S2����O={�= ��*Zc�m�=�0�>nC>�M�,H�]3�]df�u(����^�DZ;;m����4�/Ά=�+��������q�	�G���F��HE����kt�W�P�n1��S���@��=�p?1hw?
X�>/1����u�ۛS��=M������о�\+��Ì��q6�G�۾8E�!2�/.���%�o>b���t�s��r�qN5��\U��F$>��U?�}��˽Ԧ���7�6�=j,=��|�c���p��dkK��n�?� q?i��8%/�5�� ,>o7(?�?h�>�3`�;K���k�>vj?|�4?�_>�RD�o5q��U@>���?�a�?�]@?y-H�a A�,����v?��?���>>����Ͼ��꽴?�S8?wŻ>+��ք�����h�>�[?� M�za>\��>Z�>0��%���-��c���歼ǳ8>���a��1�g��]A�dh�=�ٞ>�ft>YEZ�q���k�?*����|�QG{�����:S&>�e��B9?�ݾ���=�?�#>���Ș���]��3F�e�c?�Ľ?~G?�@?��X˪�>[	>��Ż�~;=���>���= ��i�>��>��&������7�L<?I��?˵�?U�7?,t�B�̿Ǖ�Q�������1�>?M�=]�=4�ʽ��#>:ծ����<W�ν�J�=	?�"�>lxq>dL>N>�=�m>�&���"��{���q���4�F�����i�8C��Ķ�7���t���vþL`�=��?���A�)K����[X=z᡾*lJ>�!?{��>7��>X>� D>�4����$�o��?�����[.�;�޾�_��&N��rޓ�����S�FҦ�`ܾ��>xU���4<_��>�)p�*�!>�@%>(�K>zI�=zݞ<5��=h�<>}i.>��'>��=�=�=?L�=��z>7[�=Q섿ဿ�]:���Q���;�\C?hH^��8��P4�~�߾Ty��ê�>V�?O�R>��'������Hy����>q�E�x�b��'˽�{#�1"�>ˀ�>`�=#.���
�A,x�𽱤�=KH�>��
>�wn�"��F��}�=A�> ���b�=��5>ؐ?�I�?Ҿ�>jw@>~�>E�h=��>���=	R>���>/�>=�
?��(?�+?��>%6>�8���g�>�}>̵�����=E�]�B���S�Z>k�
�u��=�`	�/8>P�=�4=�U;�ͽ?����=x�>?�8?i��>%��>�9�m�>��M����k>O���C�>5�>��?��>1��>5>i�`�Uþ�R��8�>b�@>d_���w�:��΢w>�s>��O?��1?F�h���b�;��<���=�!�>o�?�I)?{6�>);>Cɥ��� ���οr���v8�!83>�����!�����Wh=����I�a�{=#�_>�U?���>��>�X�>&�>�e�>ed�>]>�7>e/==�6F��3�Np���|u=�ᖽ��]V����=ō&>�-�����)3<>L�����=�ٽ'?<,?����B5�2�A�)�ᾖ���3_�>��>�;?~{�>۵)>f����L���8���x��>�[Z?�+�>�ג�B>\^��ׁ,��r?��>		�=z'��M"����*�=��?��?F.�>������t�q$e������>�G<<���<���?��]?�
��䫾�t3�U/A�&@&�t�!>�r�������B��� ��>������������t����>�&�?�畾�I�=mwžF�����R�!���?8�!m�>4��>��M>l� � ����2O��9ؾ��㽹�=�� ?Zn�=�W?#?@?�Ia?X��>#�?��@���>x��TN>p�?�f>���>�;�>��>�Ԉ=���$=���P�5xx�G޼�5ٽ�� >��=�;=<7a>�b��;�@>$�};��=�M>VX>�I�=�6�=�h.>O��=*�
?I�?��������:��e����=�ӓ>=s>`e���@M�ѻ����O>mZ?�,?v��>d]x=�L̾���@i���G>t�?�C9?���>�mE�辶=ރ���I�����=9�5>tS��
2��O�򾕫žy���w>�~u>NQ�=!��>m��?��V?�Qd?]SN���)�/_�7 s����>1��=Z��=u��>�ٺ����I�5�O�Q��H��r8�݂����?�N�E<�~�=�cU=���>O�S>d*�>VM�;�����X��u0��@<=�It>�Z�>���>�Jl=��h�g�վ����I�i?�fҾ�j.��[��x:1����߸?l��>Q)���g??Q=�JB����^��1?�^�?�9�?�}�?D,p��������>o��>s�>R�ý�zk��ػ���r��>fg>]�����K�C�LU�>��>��	�F&���	��q<}洿Ӽ0��;*=�쨾R���D�þ]<�G�I����aڭ���U^�Ž��?�����7p���̾�Ҿ�+�q.�?q>{?���>��#>�-$�ځ������PM*���Ͼ3O[=m�ű����?�������!���O��H���#��>􅆾l����u�$�_��u/����>�E?����3ɽ!���Lr�<3�>D���.8�C���䉿�ᏽ�b�?��j?���]����"��>C�Q?%�>���>v�#>Wx��'�"?SyS?foT?��k>@K=�ɮ>�`Gp>p&�?��?�sH?8k�P2R��$!�DʽO�#?L�?Oj�>6ٌ�#jɾ)<}9?�]\?~�>������#N��Z?:be?9�%���N>)��>�т>J���$[��6
��7��c�z;�l>+@��2x�~Z���i_�?��=��>�z�>�\齮j���??Kaؾ�du�O���*ԾI��>j�1�?��
F��#?��7>����$_�������b���6?�2�?�FW?�9?z?�)U����<���=��K>��=͵=B�
���>��>)F2�N��!F5��?XU�?��@�O?�[���mӿN0��L����8���U�=�4�=�I=>ӟ����=�E=(���Ot���>d��>�%q>��x>�AU>�=>�d0>Yi��B�#�����͙��jB�Z��t���g���	���x�����i��+���Mϥ�6������wQF����ˮ:�]!�H��>�X?�H�>ӊ�>�>HyD�\���=v��w��v�ڤ��!�Q���`gd�b��b�޽��f������&��@�徲�>�����+=��>_u0��R>{F�>4��=�~>Y��=ö�=��	>��=�A�=�<w= ��=���=͝{>sP�=)%�������A:�"nQ�v��;��C?�(^��x��|�3�U4߾������>��?�S>�y'�������x����>� G���b�P˽� �M;�>��>}(�=�dԻUl���w� ｄK�=O��>t}>�l�⏾�#�_{�=�1�>��̾�1�=[ف>�*?vq?�2?�b�=��>\�L>n�>Ҿ=��<>N�Q>��>x�?�9?s/?�5�>���=�ca���#=�R=};�jR��Ͻav�%�8��%;ʆV�n�<I�=iw=�-�=�5=Ʊ��{ ;��<=�x�>�L?:��>L��>��O�;�1]=��10�Z�e>�NĽ?J�>*��>�?�=?D��>g��=�@3�ŝ�#���q�>�+>T(L��@k�.����k>�R�>,�F?ˬ,?�E��L�����GP)>~��>�[�>��"?繱>�c_>6������Կm)&�[R�fV�g=�B}>a<��E>�}�B����2�>��=��"?���>{��>P:8>���>菱>�t�=��=�d�=�k���=�s�<�->����F�����V�>��7��=�� �XB	���	����F��]��v?��?�)a�%�l��TF����U�G�&�>�I�>�1?��>S>!�C-Z�V;2�ȡ�HF�>�X?���>�r���{�=��"�H{�=o$?$֯>T��<��{�����o�~>�ӡ?2?���>|�D��yw���f��<��n>w��+�0��h�?�%G?ef�1=ľC,)��E�������=nf�u}�����e
�xM�����q{���N��?W8�?�<T��,�;/��{����\���F�H9�= �K>EA�>��S>3����{���*�Ɵ׾���/�'>}�>��#>��?���>]y?��d?�0�>���>�%$��*!?l.�=(�D>m*�>���>?�?�?�?>?�m>Q_��������t��
���˸��>�>���=G��<K�,>�..>ϔ
>���é�)�����;5�f=e=>w��=1��>h�?S�?f\��=j>{Q>z��r��K]�=>��������4�!��w$>���>�u.?��>,M�=́����߾� ����=��?��?B6�>K��	�)[ؾ�D��23#=��x>7ઽ�I&��͔�T8��?�ʨ3>��G>&�>��>�w?��m?8�I?3QT=2L�����jE_����=@��=�q�=@5�>Ѻȼa�{�">�v0`���;�SC!�QŊ�jr�����<�y_=��>�l=>���;�&>�8����l��)�<Z�=�Z�>]�>�?��6>\��[��R�꾵�f?�碾����˾�*0�w�R<���>?J��=�<?Q�a>"p��Bܳ�5f�!��>�C�?���?7F�?����ܾ�ֹ>^��>���>:,��5�����='���=�8�>ڬ��+��=���>���>Ԟ�>� ������c=𶴿�T>�Er=�G���Qp����������|�������X��!ҾT-�{R%�^����<ӽ�]f�"r�G��%�����?x�?�/�>�@�O8
�O�.�ʺ �*�þ҄=�vϾ{㞾ښ׾;�6S �߆'���.�?8�q�!�@Ǣ>��޽�fu���o�e�?���b����>	X?"���2h��Է�/<n>na?��5��4�� ��t���ɾ�q�x?�S�?�*�ahf�=��B[>�]?��>�>ZT�X�ƾ�J?-J? 8L?P�P=;n�{0Y�I�	����?B�?��??N�mmB��j����?Ig?���>O���c�ξ����?�2:?A��>+���������8�>>�[?L�p�]>�
�>Jڔ>��j���@�#i����o��3>M-������i��_<�ȫ= ��>]�|>oOW��O��W?��������S�ҁ��T>���=`�?{»��n�;���>SJ>����!p�b����#��F?K��?u҅?�!?���#�Aм���(7'>F��>j[=��$����>0��>L�/��=��@YI�{M?���?��@�u?���\Կ��� þ�.�1�f=C��"�4>s�ӽԽ��]W>���=wB��*>z�>��l>Oo>�EH>�W>m"\>���k��F��]���35�*�1��� ����PU�:b9�\�꾐;��_���v$�h@�����:3C
� �o���5�i[��:>�§>~��>��?��>{!V>����(�#���.��x2"�ݳ�S � ���"\,�,2��§�xִ�����6�Ҿ ��>go�=?�>}9 ?��K=��6>o$�>?�=�I�>��=�@6>���>ݭ�>w#>�V1>C�>���=*�{>��=�ф��ˀ�0:�r
R���:;HC?��\�mw��S�3��޾]����߄>ԇ?˄R>{y'�ì����x��$�>�I���c�W�˽�� �or�>���>��=�wջR]���x�����=���>.+
>,F������w���Қ=���>��Ѿ���<I�>��*?ȋ�?��L?g�W=Y�>� �=n��>Uv=�sk=��>���>�v ?�@*?~}!?ګ>;�$>U��L>3�D=�`��Ŧ���U-<m<��L1�=w>�<m��'�e=o���Vn���p�P��ԽS�޼��^�D��>T�a?F��>�?g���$j�_�f���=��>���;�$:?�v�>�V?o�?�s%?W�{>�a���*���>�bi>�%Z�,f���7x���>xf�W?�0g?�f��N��¼;fm=N��=K��>hz?���>���><Į:����dҿ���B�F�Gh��7.�J��<n�F���v�.	�>�dM<1������G>��>�>�H>J��=� =���>T2> >C)>��e��	>%�9���=��<�ݘ���5�8�$=��n��+i�
Aн �}��s޽����\�?��%?l �Iu�^̞�;���yn��d$�>`�?ɗ>~�>
>'�վ�mI�f�El���?dT?�õ> CU�D�'=�4���1>��	?G��>��\>ڦ)�x\��z("�<����?�@?xwq>�ှ��n���t���#���>�y�<Mn��΍?�6?�G��(��80'�W Z�?���OE�Z��*g�`x��o�C�I��%�r�a?��_\��W�>���?��X���-�����z��wqx��&���ѽ�m�<wM�=
���U�Q��>O=�h�׾V�ɾ�EüI�>J�=�C�>q83?�9L?$�z?��>bM?�F�=�?{�>:�>t�?��0?4 S?�Q�>ق�>���>��<E{�=F%)�z�žr����_ͽg-[��|���J>�X��=��8��='t@>�s�5~8��Ձ�.ׅ���ۧ���,�=��]�?�?X�0?��4��%|>��>*���綳����>��>0[�A �-0w>Y�?u�)?�&Y?�m�>��a>�.z�l�����5��<ُ? H?S�?5��"��>�����޾�`d>��3>��;=6����G꽨@R��)[=�>8^a>B�>҆p>A��?N?&��>��r�������9�a�r��פ��J>r˾= ��悽ir��/�q�?���ݔ��;�G�t�L>��˽�2=�a;�p>�>+>CXY=:3B=;��=JV�=�d���,�=�e�<�{�>�?oS?�cI>2N>vm���O徛%`?����!@/�!�Ծ��H����g��>�xK>���I?����a����Ͽtn\�|�>�s�?��?�W�?�$t�K9���N�>�G ?؄�>���赴��C<�����=�u >�	�q�w� �!���U=��r=���7�sG�aJ|��:���H�&�=Q������\�ξj?��_��-���������)Ƚ [*�EA\��"�S�c�b`��-ھvʾ9~�?Nŉ?�ު>�(�=AﾣT��"�t��v�ʾ+�\��/ݾf�ҽ�+�
Ⱦ�õ�o���S,���5��� ��>�v�ի��$L��1a���P�5:�==�U?���%&�6���>�E>V�����,��X��ٝ�=\���Y|?Cva?���r�1܌���>fd?}W.?���>[��8�u��a�>��*?y�5?;H\>�E~�w�c��u�;��?;��?oD?/YR��DL���
�h�k�?�@?Du�>�z�U޾�2 ��?�<?.s�>uQ��Յ�,�~��>�<k?p�5�̒->G��>�b�>���ʉ�Y8�霾h����Y>x崼���J�x��@�v}�=נ�>ő>Z!'�TȦ��w�>�G/�N}���c��Ӿӹ��qn<��>�#�*�%=�&�>�t�=^O@�����!��1B���H?��?9�i?��?����i�ץ�e���.=�>@>�>Ѧ����>���>��"�HՋ�u�O��
?R��?� @���?wm��Ͽ˓��z}��^��ߪ�=��=��T>�(�⃽�t�=Ht�����<�\>Eb�>��G>MR>�?>�Y->�Z-=cك��D����������D����).2�F߃���dU��<�"�쪾�q��x]�as=���#�����#\�}�c�F���BI>E�>`b�>�?�ܡ>(Q�>�]���(���X�Tu�Ć�e;��R:Ǿh&�������H���������!���?�u�=�U$=97?W�=�*����><'�=x�
>.�>v�>L�>�G�>�f>�ӡ=�V}=ݥ.>~>~K�Ə��䌿�,<�/r|��!p>�s?�ٽ�L
�����׾R�[�O-�>�2?&�>�4�����c<�O6?�HA�C�������=Q��>��>�LL=fi�59��0�6���i�b+=&f�>n�">EG=q�����!�ݐ>�>�f����>�M�>��?���?�nA?	������>!^Q>A��>3��=�>Hp.>Eڝ>Y�?�3?��$?)��>H< >dQ��t�9>Թ�<��~�E������Ǽཽ0�t���I�j�(<FZ�=�h�d��<��o�~���S(��A��n�>��X?���>s�:?���>�?~�
&S��5�=��>��i�Q"?S??=�
?��?q;?D�?���=�.�K��<��>��z>�g;��a�Ѣ���P>�ȼ�z??��S?&#�=���=��
=�A�a�>8��>�LM?�d�>���>	%�<M��!lӿ�$�y�!�����Wc��b�;�<�sN�
�6K�-�0���l��<4�\>"�>�zp>��D>�>�%3>GR�>�IG> ل=��=�_�;g�;xF�^�M=����F<��P�(��2IƼ����G��i�I�@�>�>[� MټCG?u�/?K/���ɽ�Ep����ھ���>��?8�?e��>cQ<)'���?�w��� �=H�?�zk?*P�>jV��i��=Aخ��YR�7[�>3�>���>7�h�>�Ⱦ����}����>�X?���>a[L�%⃿���kz+��Š>�l=#����?`�S?B�?�S�J�W�D���,l����0ǰ�C���O�5�ٴ=��T�����^���= ��>�Ƥ?-�?��JR���؛��͊��h9�)�f��v)>�>�:.=�f��O����	X�Q��q����;��>?�R>`�>�9�><n�>�@?n
?[7?�����?^Hz>��~> �?�g:?k�'?�#?2��>\e�>�4�=���=+D�A����nb=0��=��r=�T>�~>���R�ؽ�;�<�޸�ey,�᯼z�>�7=j+����=j�9=��	>��?ߚ?�)>��)">�(H>qp��:O>�X>���<R�Z��o>��>��0?3'N?E�>nw>���a��A`��;<I+?�<[?ԟ?
�_��>�u���❾Bv�=�}�>�0>p0���,����־�1�:?p>�ʔ>5i�=�8>!�X?^Y?���>m�ʾ�b����2�b5@�*re�5"�>�@-�󀖽�s=�%
��]�0*��Qi�w2�l�K>_w����=�~�=ڿ>�a>>h:=�
>o��=0�[�9O�0H��;�6=���>��>�'?/A�>�s>I���z���-D?q�����&�s~Ҿu�	����e��=:��> m:��l?��p=�֍��T��7�i��ݽ>?��?���?m��?S#j�t����L�>C��>F��>�-˽��?jL<�h��@%>f$>t������м�,>�"P>^۽�;��ś���E�n*׿;�U� !�=~;�F߾<���.9 �fVF�3��|?���6��X����/:�?
�)���ת����M����!��1y?�V?�K\��(��`�$��T���Ep�>	�߽qf�G=�������̾6���"����#� �:���~��p�>"I׾���{������86>�9�>��O?l���T
���վ G8��@b=��#>�@޾�Ip��	��KH`�^�Z?�7N?�>��1���+��tB>]�?Qɻ>@g�=��Y��b��A�>��?���>��='�e��^�Ϣj=f1�?<�?F�C?�D��3�U��l��'�K?��?���>s~��l�پG#���G?O�'?\Z�>��al��`"��J�>�hi?��2��5>y��>�0�>:�Խ�"��3򧽰������Y>Qj;��ڽE���l){��QN=yu�>�>0˽�䞾6�
?�t�"\y��C��b���Al=w��1?x�˾�[�<��>B�V>2F:��}����M���"�Z?5ٻ?�Ah?S`?��W�h�u��?"��g�D[+>i+�=��w>O�����>��0?uY?�E���apb�5�%?��?	� @'`j?�r���@п�����PҾ`eξ�``>av�=�*l>`��4g>���=@c�M����	>F��>V�>���>�$><�%>N�=�$��f="���������`Y(��������78n�y�澺S?������վ��о����q�	����;!C��<��|�������2>%D�>���>��>{0B>��=>�.��;~��[��7��,��O��M�����v���H�c��Ͷ�.r���p��>KD7<��=XI�>�5�<����܄>�1�=�3>=�>	�!>�P">�>4>�r=�1=K>��>Ux{>^��=���%���c:�R�Q�g��;��C?ˠ]��A���3��B߾wd����>=�?n{S>؄'�"�����x�Q��>pG�k�b�q&̽&^!�mW�>���>ʈ�=��ͻ���w�)�G�=�g�>��
>qs�[�����.��=��>񌕾Oַ=[�7>Cr??r?�8?ʃ�={1�>��>\�">��>}��>S=>Tя>:p?��2?�d.?B��>_´=����(�=���=E=�����+S⽽=���a*�}��%����=]��=o}껞H�=��<}��s�ս�[�=�(�>�V?�_�>��6?��=�Ă�qX�iN�;J�>֗M>>{�>�>�?��?G�0?Y��>�X�=ɡ�� I)��o�>�_�>��;�YC�������>	b=C�Z?���?��i>�4Ͼ������>��y>"3�>Z�?�?+�?@���� ��Uɿ��E��7:��{�=v�=�ۗ>�ξ�1�<�Ŋ>x�3������QŽ���>ta�>�/�>�#�>�]=�$>�3�>���>/�>k_=;꫼��k�'HX����ү4�Է@���<�y��kg<�������,�I*ν�/۽8�-���?�?m��^���"���1[پ�S��`[�>}.�>қ?L/�>�h$9n��j�S��x$���@;[Q?Kk?�f�>�y��ԧ�=�(�&��=�m?�y�>B��>�zc��������������>O�;?�)�>���Y�p�����]�+�`s�>seu=0X����?ߺP?�Y��H��!%���t�H ���5�V��,���5ʾqe,��3�V
��!�CR��e�=���>!�?Y���N#�^ʾx$��с}�Ef%���(�m����K�>�]�=�k�;]Q���9\�
:�
FӾ+�t��d�>O�=�>�???�Z?K�?�6?�2��?���=��>��>.�?[Z?5�>��>Q:w>��n=���!��������Q�e�ļ�e�=V
>�2>��Y=_}=���;��</a�d����ae=�=p	=?��<9�=B|	>w�?m=?�(���>��G=:fy�X��=�
h>\��>�U!��ɾ��>���>\"?�hc?�?�B�=庾g�׾�,�-�I���>��i?oe?�����y>m��.���5�$<�>V6�;���_.��J���$%=�1I>���=�e>��j>C�r?�$~?��>��;�@��NI�s�0�Ǧ���!>�{�>�x���H�>1W�`N?���|�+{��p`2��%�=�G$�AŅ=���=Nl$>�I>��
��
q>�>c٘�=h�!�ѼÆ^>���>l��>L;?���>-6>mȰ�},�QN?'���ڼ��	˾;�'�P��<�䱽�w�>�6�����>�&�>+����׼�*{�ᛒ>.��?���?�#�?���zⅾ}��>��> �k>�XK��&���ػ65>�l�D>��>��<�Jv���枽!U�=2�Q>U���@ԾZR����˱�"�"���;' ����)�D��q�վ~�h��پ2�������h�v�-+O��Fý�(<�G�ʚ��pB��C�����?S��?0��>��5=���d	� �����=kB��'����~�:9���Y��H�ؾ ������~T.�,<0����p�>
S8��~��q�˹4��>�d�>2�c?�7��B� ���E#�>1�>kD >��뾺-����v��|�_?�jq?ݥ;��`�̹ؽr͖>��j?AM/?U�>��e�𷏾>K/F?�zF?�~�>�̎��p���<܈�?�o�?V�U?T#оXr�}	��Y >��J?@`*?NI	?�4o����n���QfB?�e??ܳ?'�(7��^���y
?}�?�1̽O(=Tv�>�`{>�	e=��yf^��9ȾKW�)�>�] �I�V��辆���<��>돠>�J��!��Ys?�I�沆��i�z�Ͻvk�=S��=��'?�@ݾ��>;��>萶>�c(�P������i$ὩA?,�?Ů�?��?�ﾧ���{��>�T����>Օ�>����Z�S�65�>ٕ?e�Q����Z%�҄1?�{�?��?�Bj?�u���[οZ��gǾ[ś��>���=�8�>���MY�=U�+>��~��_K=���=S��>]L>�ם>o�>��>��E>g����"��I��Yh��,6��������N��#�l��!��~Z���z羯b^��Hν���9]!6��7<�����3<�J�>�,�>�ђ>��*?b+�>�X�>NHӾ:�"� �׾\:��������`*�������g�ƕ���3�Ҿ0k������p?��!>�	��>���2�����?���>�b>�;>�|;>�3>V�4>[9�=xP=�L>B�=B`|>ʟ�=�!��y���9�PkP��f�;Q�C?�\�dޙ��3���޾@�����>�n?�mS>�K'��x����x��E�>Q�G�׎b� �˽(J���>�o�>��=k���b�KJw�r����=���>�c
>�L���D���X���=g��>.���Ɖ=FWc>/*?/�t?�"?�P�=���>��i>�S>�]�=���>��Q>\�>e�?N�,?�
*?�e�>��=�p����=�m=�a��
�5vY�� ���xL��C�7О߽ۯ =�xG=��$<a�=��:ޝ������A<|��>��<?���>�4*?����Zs�ѵ��GX=YB?�8��/l?��?4?��>$�.?��T>h2J��*ܾ���b?==>�p��mZV��P1>�,'�Z��?�]g?k��j7y�;�&�$-�=[5x>`��>ߡ�>���>~��>O�{>
�󿧬ѿH�����`�r���ϻ�R>�7�(����'�>!�����=���5*?,�a>���>6�>ʙP>�>(��>��b>㛧=@������2�<0�Լ�y��u��s=��;��<���=_�?A��4����PO�GK��Y�?�?q6��`���/�4*���5�����>>��>�~�>Z9�>.N�=�y��7�2��������>D�d?���>Xr~����=�h�O6[��5�>���>Rn1>g�4�����bξ�M��>��8?��>z��5p��Єx�:��a�> J�=�}���?J>?ɲ�����ؾԓJ�g_�A8��Qu��K4��᧵�I�>���\���	�9@�_Pʾ�&��j��>p��?Z{K�Jy���1_�`1�����J����3.���o�`�>�u�=�K㽹�侤�8���B��r��� �>��=��>�S ?��C?�r?�6�>c��>٢ý���>dv�=��?�@�>T?ľ?���>�މ>��u>�Α;���5�������<�H�=�=���=R
>�+���`�<ݾu=�+�=�>�/<U��6ߔ=���=��3=�f=��=T(?bE$?) ��8�o>dE�=��]��6̽��>#��>��˽�eu�~co=k�>��B?�]?���>��=-W4��T�� ��dn7��3A?�2g?��?�4���>0+�����-==�ʫ>��w=�g���/���k�bCV=�"�>Ϣ\>���=Re+>7ww?��x?>�>퍰��p����H�>���'ݾo�=�v�=��n����=�w�L�,���z��%��We��3��
�����=�)�=�W
>�)>����B<���=E��=�������=Pb���8�>�	?|y?�J5>̫=cvx�8U�@�^?������ �d����-�>�?��>6O�U�?��>������ǿ�K�+��>��?0�?(��?���1��X��>;�>y�f>�k=SD��6=�:�� �=�	�mh
��0��)M&>M��>�5>QL!�ׄ�� ��FA�W0���
:�h�v���b�E#ؾ3`ݾt�#�ѡy��8k��|�<�����򽜤ӽ����'��ku�Jԉ���ƾ�����P�?���?>ps>���=�E2��n8�X�Ӿ�q7<�ɫ��,��G����W�\�!��^������쾇�-�#�B��U/��d�>�x½Ɉ�� �|��������g�=�F[?�9���$��[ʾs0>'�n>�����M��B��r��t���s?�gk?�:?�~�C����_W>��?�,?p��>�ӵ��ݻЦq>��R?`p?���9n����X���?>���?�b�?�C?j��Y,E�2����y�	?�l�>�z�>��>�z���>�7���?��J?B�>o��d[{�|��ƒ�>�Z?NI�XQ6>���>�n�>-Ľ/u��i�&���_c��>�������0�s����_��=Xk�>2&f>���Bެ���>$���/a�R:X�������ݼ=��>'����= �>fze>}���(��:��|�<���'?�,�?�:m?߹?��ɾ�ê�f�+=��O�}Nd��o>�%�v��Ɔ-?�KM>��_����,'���>���?���?��X?	�`�$�ؿ���[���D���s�=1t<=[R�>�T���>��=ꍨ�]�ཐ�(>���>'�>�ؒ>�P>��#>vMN>������s��������M�$�X:
�.Ie�m���u��]�Lm羡y⾍?������3Ċ�l�,�ʪ�JD��;���r�X>���>���>C��>X��>��>$`��/ξ�p�#��˾羻���z0�]���\����$9K����9%�P
8� ?��5>=��=��?f�V=<�����>��ֽ�+>���>d�>��>G-7>�0�QR=�Y4>ś�=���>�ݼ[B��\�����p�E���I���	a?铢��f�@� ����S��2A>l?T�>!�H�����I죿��?�u��������5b�=�
?�V�>N��>j��=ݴ���ݼ�D˽�P���Og>�o9>A��=�¾����|��=���>O�-@>2��>u�!?���?M�7?ʁ&=:��>�+>�L�>�>�!">�@>��k>���>@'1?��/?Ii�>^�=
~��a��=��=�Nz�*���Y罎���K8����C��{�<�\2��'��9\=��0<� t�aF �cd�<B�	?r�@?�2�>�T3?T�̽�Q���!�d�P�		�>.�U>�o�>�y>0=?m@?��?%�>�0�=�оy�%��G�>�<=�W��w�l�=s�=2Bq<�J�?FVU?u��=�l����=ZX�=2�%>+�?��s?��>���>�=��Xf׿���8u&��,q�>A
�݊N>[wA���=c��=�k1��n���>7=�gw>�5�>�n>{6�>�30>��>��>&${>��>���=z��;��Y��홽�D=��:��<�)q��2����[<����ؽ)b����V���w��2s��?��?����t�=���8Ͼ珱���?m��>Q�?L F>�e�>�y
��K�z���+ >[#?��o?���>���3�>l�C�l;h�?���>�e�=���v��'������נ?��#?a@>�Uc�IdV��6V�}o'�PX{>F_�=��t��?�b?�	ݾ��o=Oi�aN���ʄ�x�c��f��R�����]��K@����ٌ�d�>t��>$ �?��<�R���ȀQ��y��Z2��w���8"O���>>�>����h8�y횾��A��@���������[�>�%�=��>n�?7d ?i6�?�?%�3?�i1�_�E?(mY>��>�>��?�"?�$"?.T�>��#?"�>��Z>��D��࠾I�>�f��<��d>�@�>���T���U>?���(x�����< }<<-�S���=��L>�R=�> �?o +?Ѻ��8:>u �>;�����0-�>ڙ�>���4�����>1?(�E?��<?��?�z>J
���ջ�x׾"�=���>�E?G��>��� �>$����ヾ$��o�	?� ������<�ӽ�y���q�TI�>F�)>���=5�>>��?o�?3�>�i���Ry�a��.c��Yc��=)ǋ>�">����o��a�x�b��Q~�VB�5��=nC�����=�n=�
>�{�=�3�=E�=3딽��>���z�;��<l��>e��>(�9?��>�W8>酬��J���J?/૾#�d����	��+ҽ��=�&Y> /�~�%?h�۽Hl��奔6?M�&k�>м?L��?��?����E��>t�|>'�C>�d���8��$��e�����=>���=$����W��׋Ƚ.H>
��>p������;0�z	н�Q��"~4����=]���˾����g��M�ڽ�ƭ���~�t��Jd����߼�-ڽ�9-�nw�S1��kU�Yɾ�:�?pk?q�'�����%TC��(�����9�>l��a
]��蒾pd����+��z��^tg�`��`��{B�5�I��#�>S<��w���������Q�>�_>�L?|�þ8�7�g�I�<� >>
co=�ƾ��w��Ԯ�bJ��.,?hf'?/Z��ԝ��N榽6�>g?�%�>�D1�Q�y��� =+O�>��d?[1#?@K��ު��i���=�?@��?�%A?4U[�O,F��P����a?��
?B��>K�����ӾZ~���E?��9?g��>��A���*;���>5�^?�K��4T>��>��>%��:��_, �A䚾�榼��Y>b���9�w���Z��~=�.�>�H�>�	<��e�����>fH��?�קr���d��;_��>�+�>w�G�2�>��(>rţ=F�(A������.���>?�J�?��?>�o?�8��}d��]>�
T�>-W?3i?�=9�ڽ�ӽ��?i�����%`��˽?�\�?H��?(�g?�w�w�ݿL���,��������=�=I%>����=���=��<��;= h+>��>7�4>'p*>	�>(8Z>�a�=΂��"��ƕ��i��x�3�������	���Sc�1���vp�ܯ{�Ҿ1�Ľ�.��+꽑f��HI������~��> 9>=��=�y�=��m>Q��>��辡B@�C���֚Ͼ��#�  �<����T�R�޽�:��0/4�?S��� p����Ԗ?�ýV��s�>Vԩ�zv�>�>f�r�>��� >Z�f>��>�>A^�>>�>�;s>O%N>eSJ=b {�DRw��?�"r���.0��7?�`_�����:61���ʾ�C��׮�>� ?�x'>�-��s��x����>�rP��)_�#I�u���(�>���>�m�=vjT;�; �{����R�j=�U>���=���Ň�S	�ۘ�=��>�fɾ��=�1>�@?�s?V�+?�w�=��>�,>�F�>�d=��->��/>�:�>��? 7?��,?�,�>���=)�~�K�>a��=��P�� ���]'�����=2<��d�Kj��U��<Fe�:�E�<�8<�k=��.�G��<���<0f?�y=?W�>Ϗ>������=�`�>��=���0��>�l>�	�>vj�>o�J>��<��
��g/��
��\�>�3B>L�s��z��)��>ԔD>J�=�h�?��X?�ω�������>-A�>�?�?Kd
?ko2>	�>���?P�k�Ϳ5��~L�_Ғ�YGɽ����v��$'5��T<6A��kL�y?�<��\>���>�:*>�B�=Ҁ
>m�>L��>��>�y>B�={<��3�3�J�3���F��ͽ���X$p��л��.=;DM���<�ɐ;Yl�:�m�9x��>�B'?��<�=>!�ӽh���v��;2�>a?�A�>
d�>޾��q��Nia��lZ�<�ŽYZ ?�T?���>o�W��7�=�䁼���>��>8��=ݵ�>����
�$� ��>�)�>��?��>N���L���+���I?�^�v>&;�5*�1B�?+�0?����o����u`A�E��_��=��𔝾ǌ�@�"���I��d��O ��hl�W>�L�>�?7�E���0=-:-�cυ���C��	����Y=�ץ=�r>Q�ѽN<	�W��=�	��j��1���;>��?��=��?��A?��o?��l?�?�[�>c��iB?[z�.&_?�5�>�o?�L?��>�½u>���=�����U��pI���F�<̠V�4�=���<dL�=�}�=� =`S�=�%>}C�1����<h�)=���<�>�>��>J�?�+?���� ���~�>bt=� ��%-n>^=�>��@�5���#g<,�<��>��?���>>[�ܾˁܾ:��� hW>��>��Q?bc�>A��=,
z�^���A����2>M-�>���=�����x���k0S��3z>�>)S=hT>g�?�3?ubP?��&�ʔ���B��1>I�������>�n�>��>QϾ|RQ�d(u�4K��%V�:|����=�f>J�1>׼�< ��=�^>E�����ܽ������e>���=�j�>k?���>��ڼ�1��ã�~���׹q?&�4DT�x���ܐT>�c?��X=aWǽ�K?Ό��i�ߗ����#���-?��?�?�NY?χ>�G��;�*?��>k��=��=�U���8���@��&�=� >��ܾ������w�>IF�>�ș�������/yx�������G���@>7�f��;1��TW�}�:��2���!����;�i��D�=kpl���`>%�4=�`w�����a���)�	��?�a:?nТ=�|����`��~پ9\�=4����F��˓��
�^l��肾L��&mƾ�A
��B�m�ƾ��>�)b��r����u��-�D(���_>(R%?�Y¾�3��&���K�=�r>҅l<y���8��%���%���S?v-6?�뾦����Z�%>��
?���>��>:�� ޑ��{�>�%+?�O?�����/��aO��yN����?��?�J??\H�(q[������%��4?��?˸U?]�-�E?�׷���s'?�S?�e?�Dݾ������A�SȦ>�?�sO�+.�=�?�>��~>�[�=�<(����=�������=H��>����Q�=��an����>"��>�4�>����������i>� �ħ��u��>�vǏ�_A(>��>9qȽ��>�Tw<H(�=�]M���~��q�.���I?Di�?x:�?<O�?:�(�M�J�����9֗>z:_?>?��>	�==��m�$�?�Z�W�T�'Ѫ�Ue?Aa�?j��?�w?t�X��ٿh������\�����>�I<m��=+��F=�Ub<[ҡ=6��;��$>~�>��$>�QW>S?�>��>>\�_=�у� %������
��3�Ծ�����0�V9��f�$ſ�܍��׿��bɾU������4y����%���?�;l����#X>q��>$W�>�B�>�r�>�E�>���m�I�=����]3%��=����B������~�����r���m���t6�1�?����u#=�״>ٝ���iR>H��>�,�<�>M�l>M�+>۝�>��K>>V�>���>3��>�;�=G0k>�A�=o����7:��R���v:�e=?X�i��S��'g9���о����Ԋ>��	?p<>/�-�:�����s����>�$��^Q���l�)����>jn�>�/�=/�H��m#�\~�x��ɐ�=�Nj>�5>ؓV���z�� )�UF�=}��>��վη�=g�Y>Up"?7Dy?�2?6T =b��>i�^>z��>�F�=�� >�T}>��>f?�5?!�#?d��>�=�n�o��=W=�`b��!���9�Q��ϻ��)���C�LU�<�B�=��<�d"<�(=1��<�=��s=9?��6?'��>�(�>�����i.��8e���>``�>b���Ȇ>T3>x*�>z��>���=*s_;m��n�+�����W��>��>R/z�cG���|�=5x>�=��?�<B?U_Ҿ
7ξ��=�*�>�Ư>cu�>���>�gA>�&>�ƴ�2�C�Կ �1���.X�=:lZ�C�3��"�#���[B8��Z	������<�4j>
�e>�h>�:J>�>��2>`�>�O>û=E�=Ua;�B/�W�%�'1��S��(z<�����;���4���x�P����E[���;N<��?�=?^=�3�<,�w+�bm#�j?�i?��7>>��>c�T�Ӏ�4_O�j�;�<����)?�n?�zc>g�5��?B>��ü"w>�-�>j�U>�_>(O۽b�ھ��e8p>E�"?���>�5">��O������y�OL"�Ͽ>��f<_���&�?�53?�Q�!yE�w1!���N��b�UQ-:@������r����*����nr��Q�H�?t>#��>���?!p ��a�=����������TEK��>Q�o�}�>��t�A�½�p��U�����:V��N(�>p�>�\M=�I�>�DW?j�p?]�T?��"?��Y?~��X�>C��<NT?!�(?��Y?�0?�N�>�|�����>u#�}����팾Q.=`����7�=�X��y��=L&���=',>$�?<��<@�g�=�_0=�n�<��N=�>�f=�&?�?d�����5���B<l>j�.��{,>���>=Dy����ł�6��=n��>��?�^�>�`�=c�Ͼ.#Ҿ����>>{�>��e?���>�>{9e=� �ȅ�̦�=)�>���=�!��J�	�V�"��4��A>tH>�l���<\>�х?�E?,SG?�r���/� �q�~��9���@=-��>'��>�K]�\��)O�c1��MN��+��1�=���t��=g�$>',>5�=��:�X>_U�=��;~�	=�(.='�r>R�>�:�>¡�>�x�=s����W����O��s?s�\�]<h�b�)�kɾϒD>H��>: O�$®���?%�Ӿk�n����ʦ.�&&7?{u�?��?6(?2=�>���G*�>�V�>���=�J��������̽��<��=�^=�~���V˾Y�\=WG?-%?�T<��K���'�V[=��ֿ�R��O�9s׾mg��btF�'�&�\��+�þ{��=ۼ����w���<-��=(���F�d���羖/���M��?w�?^d�>�����,�b�o�b4<���m�[0>X��m���w"���j:���\���*�|�.�A"ྍ^�=y6P�%	u���c��mU��������=ߧ�>��p+Ž�,��Z�=�dJ>J�	.������ݘ�A:��jSO?�F0?j�����Ⱦ��=WA)>�?�>���>���=]�Z�"Y4<� _>{$?�*?jP��6Ǔ�AɁ�[fU=/��?;��?�I?��;�R��D�eL�C?(b�>7? �G���$�e��� ?ucN?m�>6徵����8��t�>v�?S�O�b�J>�*�>u�>4��D�*�x��=�оi�.���>�Zν�J�������z�mIL>���>0��>E��Ns����>�v�2.V�Ɩf���6E"�ڒv>�Q�>>����>�&>�=S9�����
��ޛڽAw_?�լ?�?�2?����&��Sֽ�	��(26>n),>=�&:��)� y�>�>�;3������6��� ?��?�s�?T�S?�O��_���!�������=.��;��=BӮ���>��E=��h=�J<)k(>�e;>m1>��1>�D1>@��>yN>�y-&�-���(���O�!�9�~Z/�˒�����mAU�a� �G����־��W��� ��b����\��R��<�ϾB1�=5�>��W>m�2>��#=��>9���=V��EM�Z����-����Y�̾�=�*R����6�^E=��|}����<��C��?��<��5=���>
���^>c��>g�:=`�%>�cN>o�L>BK?@>n:>-�7>���>d;>���>׎5�xo������l�D�`�f*2>c�N?^TO�z�x�cN�c�������R�>�>s�>��;�ϲ���96��0�> Y>���ݾ��$��7�>��>$5�>q�}=6�&��2�WKK�렽q"�<��@>�)Q>��;� �D��jѼNg�>ۢ��Ɲ>�]->?M�t?�|&?�f�=��>��O>�^�>�i�=m�>Vdw>.t�>S?��:?5?Ό�>�h>#a��!>D�=Ysy�����r���R�����9���OZϼ)�|=�.�<�N�=�M	>��2<��=�Հ=��?�w-?z0�>�	�>S�_t��fZ�D� >7z�>ް���g?�b8>)�>��>\��>%\>?#��s��x���%!�>GFy>�*h���3>[�>u؅�ߌ?{g>?����J� ��Dj>�d>���=��(?^�:?�"�>}$��,����ymӿ#$�]�!�"5.��S�;�<���M��v�7_�-�6���GJ�<��\>��>+�p>�E>��>�<3>�U�>@DG>c��=\��=͂�;9�;*F��jM=L"�oG<D�P��q���$Ƽ=���5�PEI���>�6"��	ټG��>�&?򔽛is��;���G���gԾ�Z�>���>��>B��>�ѻ��L��{��/<��i�1?Թ�?I�>(H���tb>9�ɼ��>�nX>��=R��>�ͽ/�����j�|�m>V?8�"?�>�XD�*���◿��-�`X>�r���_̽�Ř?[�R?����b���#���L������=[��A@E�ּ��-��n}:�u��i"��W�����=���>_��?�v��(�=s5ž%-����l�Wf��U��=�\=[�>6�>�>I����tL������UA�1�"=i��>:xD��2�>�`?:r?h v?_'?��?���8Q�>����tX?��>� d>��!?SK!?u�l�d$>�F>��y��7�ix��}��=U��?>ݐ��E�<�޼(��:z>Z>%� �/��æ����>=?3=�T=���=�=�!?��%?����chg���*>ۨ=�P���>2	�>!�2❾ă4>��=�>֬*?n!�>��y=x�ھ��Q����=66�>5�?�l?_n>�;>���+w����m>#_>ǚ�=������j�5� ��>�>�>1��<]�B>Iӂ?�=,?8�K?$	�D�)���U��#�����,$w=��>�<^>��=�;���L�F���]N_�R,��֧�8��X�޼�9�=��R>KȽ�ۖ��s,>�&�����=�O�-�>�>���>���>�/�>��=j�,;�S�mq����$?��K�#P�8��|Ȁ���$=�4>��w�o3�X�=�篾����U���%9�M\?�p�?B��?�b?�	�v%��?�d�=d��>�|�<���f3k���S�j=8.��!XZ�����E�I�_=6=��>N�����^�$���XY̿�;���V�>�	�����h��-!�Bs*�at�v�>����%�=i�|>NC>󤏽�X����8�8����#?"L?9�>�S���t�HD�jo�==������@� �ﾜ���Ft��[o����`�þ��'��� �h��Ҋ�>a��v���(�o�TR�
1���>�? �G����/0����<��>H.~������k�J��}���\qo?K?���;�$��I��=��l?�i%?�u:>U�1��ꀾ��	>�4?N@;?���ye�n$_�a#v=a�?jP�?�R?����Ut���ܾ�>�=�/?��$?N/�>��f�;?��ş��L]?� N?���>D��e���(����>�M?�il�^��>��?Ȯ�>��q�t�<���=j	Ѿ9ܨ=jx���=i^3��ӹ}��=�u�= P_>�b>G�:0X��E?�VT��ˇ��0F��p���*=>	Y>��>����O�>,\>?�>w��)�����zhh��/_?Ӥ�?��p?��?�4��͏�v���G�<H��>�%�>Zc���=��C>%��>���������E8��]�>Zz�?��@�6V?���$�ҿ�᛿��0T��)>R��=-�>������>�t= �==nZ�;�>��>Q�\>��o>��W>��9>�>�?��*��<����E�0����`��k"N��c��y.h������%���o�������7�NCB��*	�+"]�>g��?�,>ॅ>C�>��>4b�>�j�=aV��2�A��/��";���G���{-�-�YΡ�i)d��T*���1������	�
��  ?�sv�
�<�>�`�aҘ>�V>���<���>�p|>9�>��>?=U=�#>��>N�>��={�p>��=L����~��~0���k��_D���@?;	>������7�т來�Fq{>��
?ׁZ>�&��p��(�u��c�>��Z��Ia����D�/�]%�>���>��=�=����f����צ=�2y>"l>ҿ��-���(�]l�=dA�>k�۾�� >�>>`!?�w?�.?�X�=�*�>��4>�Ï>F3�=D� >	:->B�>F?��>?�K2?�M�>ϔ�=��^�R��=$Ji=]�O��/���v�
7P��^�;�3<M}��i�_<	�=BF��mo"=�5�=[{�;52o<��;=���>��6?}��>.�>O�r�ɔ:�́]��h��R+>,�-���>�T�>#�>w��>���>��G>q�t�b˸�������>\d(>:3D���t��ǽ�g[>��=>; o?�T?X-E=���'x>VE>s�>���>5?���>�mE>�R=I���lӿt$���!���m���;�<�+�M����7��-����_��<��\>��>k�p>�E>�>�;3>WU�>KQG>��=x�=p��;�U;*F��pM=��fWG<u�P��v���ƼQ���U��[}I���>�:�JHټ��?�>?q��b�u="'����龶E��?؈�>lT?Y�?��{=����d���*�Ň4�7?�>��??f�>���_�=	"o���'�	>v�>Uf�>�v�<�_�)ݵ��BH>y�?�E?���>���]q���o�mw��"��>^�J=�<�C?[?"��_r�N"�7$@�P���I"=�й��Z�d7��ī!��/5�Ӵ������N�b�@צ=f��>�q�?�f�aQ�=_���ܘ�����-��\�)=0 �=�e�>Ծ4>��!��}���7�ѵȾ��6��c5=��>��$���%?��A?�:d?�C?�S�>mk?��I=�r�>�H�P?���>p��>�:?D��>u���@�<��<~�$��8u�⯃�j	�<�����K>֍T=�=4>׶�<*j=���=��4��so=��/�ب�=�x�;<�>V(+>�v�=���>�C*?��ݽ:�E<[�w>>�b�����&[�>q��>W�������-���O��:1�>�E?�0?_��e�C;����׵�=��?��S?�0G��G=Q��=�s%��O����=n�>N!ϼ�[��-�3�]zE��޴=EmS>V�=j>�Vz?�1?U�4?1޽���e�g����<�J���<��Y�>�
�>�[�<O��1�&��g�o�_��:�Y���E�?��<S>�`E>�W@>v��=�NB>�K=Hq����۽;P�=��[=�C�>{�>���>��=�H=�������?�	���s���.�퉖�_	;<�Cܼ�-[��-���=Α�%������כ|�g?�}�?�l�?�cJ?ҍ�T��ݒ(?�[>o�N>[	=(������l��=�&�=/�ս�W��Z��)7����>*?�+=U��5�M=��ٿ��.�a�>�p+��,��h�Q���9�gb;�8>GMþ2����GM����=�����Ƽ�d���Ǿ���qe?>�g?� v>���y|�0����콺����9��2���	����k&���|�߾ qƾ{.�<C���y�>i��"�a���m��k~�>�j��>�_?�׼i��=���e��>�?�,;=6��Xs��a��v�n���{?�@�?�WH�'�}����>G�?'�?ʲ�=|
ս�IH�*�3>g`h?�aL?t�<!HY�	�`�W��'%�?˟�?�n?�uV��!��	'�9oe���;?:?\�F?"��<����L���MX?;q�?��?	�%�Yᔿ��<�0�>�9g?��F�-,>���=8S>���>;���S%��O���E���G�>%���!پ���$��T�>�g�>S�K>J�K��/��S�>Pb�I�_�g�f�����4'󻐙�>�� >a˭���>�����>�������~��5\��H?�+�?gf�?�o?��0�D�t�sG����>�?x�>{\�4����=�
?���a��(���}�>��?/h�?�n??�~:���ؿ=ߛ��ϧ�+���Xx=�xs=�>�=�w"�{ɖ=�Ǝ�,n�=#��;��=���>G�e>��\>Z�J>�2>�@7>τ�Gu"�T���X����"V�^C��"�M����x�`�ES����t��oo�o�½��)���Z��6�-p�����p�/>�8�>�/>h��>��?p1�<���K@�c7������!��QA������$�����Y�Q߾���O:�O��|X�>Pjٽ(O=��>Ә�=�ӈ>OM>B�q>��>(�S>ن��+d>D�\>wRV>�lC>n#T>%%>SPB>M�=�c{�а|�3A�"g�P=i��2?b>I��Ԛ��~3��پ�����w�>�?99>(�+�2k���ҁ��l�>�0f�)B��:���r��#�>���>�l�=!��;Lm1�d���L�KMc=��|>!��=j�������"�r��=�k�>��پ���=X�_>�q%?�Gy?
�2?���=i:�>��f>=ŏ>�J�=(�+>��\>��>�?�4?�%?��>���=|�o�=1�=7��=}c[�`7��CWʽ��Z�ki����<Q鉽k=e1�=ɗ<�C6=bd5=����<��=��?��/?|*�>}�>�����ɶ9�Ҟ�=�lo=�R���>*?�>��?��?���>~|=}���8�ν(�c�A��>H>w�G�E����O��^�>� �>��s?I�S?X���?���5�>om�>��>��"?S*
?�51>[]<�N�qF�̰ϿF��P%������3�D?���}�z��vS���ڽ1���J�h=��5>�|�>I�q>!��=�>	�T>K��>���>��>&� >�y���^��U���<��X��n=`�[����= f>��E����N2V;�I���
 =�[\����>p &?�(?=c[�>:^-�R�%�ӹݾ�?l��=z�?r��>�,�X�Ȇ3���J�fX��[2?&�e?6��>FS��X>h�X�tW���='�N>�C�>x�>�?q>⯌��'>�H?A�W?+�>�����L�����]n�mѮ>�<�< �ۘ�?��B?�6�tCH�n���B�/�+��]�>���a���g^���4#����
����ľ,S0�}є=��>�|�?P}��!>�	��x3���im�Y�߾�����/�=D�'>sq=4��euʾ�i��۶���w��>/��>��=�@?6��>�C?��h?���>;?�Z>G0?|.��&4V?��?�?�<?ҟ>���d���T�^>��o_3�54u��Hn=&���CE�=t@=6خ��u��с<����kь>@��9p�����<�o=��i=���=>�7�;p?��?����p���aM>^␽G���!W�>B�>;�J�e�h�<��>܃0> 8?�J�>�q.>N�	�������>g��>k~:?(��>X6=Ũ������D����>O�_>�i�f�ľy��W�b벽�(�>o�G>ݮg>��O>ra|?r76?�L?f뽷l5��d��aؾ�����3�=88�>Z1>��>��Ҿ I�Y��ҧP��C���������-��)>�5g>�wO>�>�=��b=r-м㲾���=�=�'>J�>�6{>ϥ?��(>��T=+�x���LwS?Z"1�X>�����ľ��~>�/>�쏾gdٽ
�>4޾@k���픿j�9�܅?dc�?���?�6.?Dw>�ۡ��?2��>�_i>��Y�%Y����U��b>4��=Pp�#C�8����X�>���>���B��ʾ&��((ǿ����=����(��J���⾸�R�0
��1��02�������պ_W��¾�\��7�W�[?�c?�8I>[��<R���Ğ���c������R��t�+��Rmj��������V��������e��$�;J�83R>yW���p��t�,@��,ѽn�i>�?c�����l�):��=�z�=���� ���E��0�������4[?�S?� ����kM0��O>�"?���>=�>�ꕾ�ꎽ��>A9?��?�Ͻ���D<t��\=O��?���?�\?i\>�hK���`G��"?��L?8X>?3U>�����4��4C?��?~�?�킾�������*>z!?��g�j!>�@�>ۭw>��=ݻ��P=����4<r=Z�Q�6Y��Z9����"��c�>���>!>>@��k���T�>N�ھ�<:��E�8��D�g�:��<m�>z�*q�=�?(>h�=Q�9�d�����[�@�}?9?gm�?�#Z?�B?m������x~]�s�ؽ�n�>V>�>�k>���P@�>��?�oǾ U���׾{�&?���?u��?IR?�7_���ҿ![����帾�k�=O��<�=]�/�&P�<ݣj�|5��X��C0>U��>\$�>þ�>;9>��>�2>)���T*��즿rx�L�5��#�����R�A�B��Ͷ��������L�����Z=?��Q1����������7�	 ����>��?���>G� >�j�<��F�<Ͼ�<�x�=�����e���&�5G8���5�ָ���쾈P���|���w�OϨ����>�`m�h�=���>�Ʋ=��l>1��>X�C>�L�=@#�=�q=K6�=T#>�d>La;>�,�>�ر>tH{>b��=�愿�����9���R���;�C?�,]�<���T�3�r߾P���T�>Q�?02T>�R'�Y����x���>��D�O:a���˽M} �߉>Z��>�c�=ڻ���yy����5^�=f�>�>q���G��,�8b�=6��>�����=�>8�?�6�?h�
?���=,O�>�R>Je�>��=W�|>"9>��>+!?;?!?��?��>� �=G�����>��@>A�,�|���a�S�\��_=�s�uw+�P�>^��:�"�>f[>_�=1퍽⶗��2/�� �>�
J?-��>D�>��>.�$��!��\��\��>�01�&?�?�A�>?'?��?%��>G|>�ξn$��>�o>p�+��7k���Iu�=Ι�>�H?4�=?g�{>��-�n9>Q <B�Z>��>R�<?�?�V�>��<]/��:��f=��Xھ��o��d���4���~M��{����۵��G	b��C\='r�>���>A7�>���>s:>/�=ħ�>Y�[>q��=��>Ф�A��=��=4�=��#>�=�_$>�U=��ֽ�����cv��
��f <>Py�=�E�]?�'?��1�D��"�J�7������>�}
?��?@0?zS=�����-��=���=��"?�c?<&�>k.��U�=�XE��:����>֮�>�Si>����sL���O��ͽ(�>x�5?{�>2���W�gs�PQ'����>�Y��X½|��?[FJ?5zܾ�ڽ���%�	�F����X��3��@����{ ��d���_�ڐ �r�5�(���Μ�=h�>* �?~�O�=ő���!���4�P&k���=[z�<�r�>~N�=�bD��g��g�O澀+?��==A�>�tB>���>��? 1?��o?��
?f=?�ʽ�9
?��>hԳ>��>P)?>�?p-?�,?=(?��i�<�ڼ�ҽ�˛�*�����H=A�>�F>�f�=�g=&�>u��`��<��V�d\��&�>���=cG�=z�0>��w>8#�=��?�20?��=�!���>.j7�YX�>	� ?n~�>���>O����3��T0�>:�'??�Z?��&?�M�>�����Ͷ�R	Ⱦ����m��>�=?���>4ʰ=��0=��
��=;Z�>�A.�Cڱ��_/��F���Kd�ϡW�yxi>�LL>c	�>��>�ɀ?N\;?ˋS?ZL>>'?�������$�Y��E������>)ժ=�$a��B��n�����e��H�0$��������>�͙;��<nj>�=�e�=m�=���t=�Θ'>�x=Hh�>��?�?�a�=�+>�R��ۗ�wI?�]B��#��Ĺ��p���
�)$ >o��>^*=��?��7<tup�`ͥ�*c!����>��?Q��?Agj?�R�r�޽Ufa>�)>�_�<	�<�V+��n_<���GV>��=> �w��S��'�>=F>"��>6d��hϾ���)n,<"{���k�}錽)v��ے������&�����������b���tG�*�ld������	�K����8�X�!���?W�?@
�>ch��C���i�O�ΖB�����]Y��ͳ߾��=�ž��ƾ�i��1!�"�p���X���8��|�>����	������J&���g�^_�>��s?�	Q�y~��������>�m>���C%ھ~	���N���à=dvr?��X?k�	�r��U�N�=��]?��?�Ԡ>I������w{?T�2?C׀?��>�$����.᜽̳?-�?PY? ʽVш�nGP����hYS?~A?ڬ^>�Ӳ���|>�i!?e C?���=���Q���	���gm?N,v?�m�2�>@H?��>��>/dX�WVO�G����(�i��=TI��=�R��s�h�o;��/�>I�>W婾]6¾j��>���;�N���H�N���R��;�</s?"e�\�>W�h>g�>i�(�����Ɖ��f�תL?��?�S?SQ8?�}��:��<=��b��=�*�>@ì>��=�}���>dC�>zC�xtr�/��ȫ?�E�?0��?4Z?:�m������:��(�� ���&{>�6>X>®�4���J/�<�2>w�j:��<_��>�� >���>W�>��>�N>�u���o'�O����_��R��H9�L�'�� �=8�(���F��c����W�E���G���G�r�
F���.��B=>�>H�>?f�>�By>}>v(x�|)վ����{����,2������v(̾<�R��MW��Si��AM��Q��S���-�>����[I>
?���I+�=lD�>��=Vs�>7�>�v�<g�P>I�>�T�>�D�>R!>X�a�s·>�_t=h<��Sև�&pO�n�<��=�Q?֮O��(����.�ʾ�o��@�>�e?�
A>��,��?��*�g�'�>���lp����� ��G�>F��>*��=�}I�8��8���eнX�f=t�>;#D>�����a���w���=U4?27���;���X>5?պ�?��?o,��F?_��>-�>��>5��=Ds�>�>�V!?Y?J��> ��>*��>T-��z<4=���=��0��'=(A��'<���i=�X�>�A��r*>[qN<L�g��t"��7��`)-=�~��ȃ=��>Y�D?F3?���>d	���FE�6����=��>�W�>��$?�y�>��>N~�>�޷>�Ww>
ԋ>��3��� ��>�O*>�x�����߾ �>�?�$�?��Z?u���;�+�=d�罾��>9?�p?綬>��?�;|>s���gӿK���#��@�=�ؽ2T�$U>���h麻6о�?���w��m_=m}>�=
{�=1l:=�_)<�h�>�2>��=�
>����{����[=�ߺ�☼�s;=8�D�=7<x��>Ћ�=~<�=_7ٽ��j<,�A���}?r%?YO��ƽ�u`����/�����?���>
k�>G?��w=J���:����;���?
x?2-?��>��?�=�K���'r�u��>zp�>��1>[G��K[�>H��x���]�>`Z4?d��>�}���J�r�}����	��>��
��E�Ъ�?��P?kų�QԺ�ӃI��3A�9$�T�)>��V��e���]���F:��mU��������e쾉�Ľ���>���?��=ʻ`>�p�b���Pb����U����M��t�>a��=(	?����=�3�>���w�0�K���>J#S>���>Vs?�3?�i?^?J��>�6R��?��=v�?F�>�o�>�\?��#?1?q?w��^�Qɽk����Q����ҽ�{C=��>�o�=�\���=y y=G�>+�=M�>���=w����p=��C>��U>�"�=b�
?j$?�v��8�
���ռ�_��E�<db�=��U>Y�+��-X�v�ѻ�U>��>u�,?Q��>���=�Y޾�������u�=�a?��1?� �>�h1�.ޖ=HT���{��Y�=�LW>�~j������޾����������>3%�>^��=�>�g�?:�M?JfR?���=��3�/�t�H@�0��=
mɾ�>I��=.6ս��F�L�J����'�-�<��7"���M�$�m>"�>x<�=K@\>ZpĽ�1�=��>y6���=�<<��<��?��i�>�H�>�8?�~�>�4>Vۥ��/"�;RH?I�"�I�	�����ξ/,=����=���>��=�> �=%C}�񖥿����Q?�u�?�L�?���?h':��z߽&�m>��=͸�.-�=�9=�g�-����=��=Z��=�qj�W#��*��=�k]> ��>���p���XdʾI*>�\����D��ō�̓���Z���_��|ܾ�u3�[��=�Bɾ���xA>%��=X������[z���ھ������?Z�?:��>�$�=0�
�A��������|½���k�=�T��K=���"�a�Ǿ9��
ʾ��	���(�%�{��>v����i�����C�q���%>ѓ?շR?�
�=���DY��x�> �o>�P>9-��ǈ������@>�hz?j�?����=0�퇝<Ms�>v?�s�>�"=��\ƾ}��� >�.�>�#�>b��=!<��n���K*��4�?	Z�?��D?����U\�G6+�^>�q?[[d?l��=�ս&z��]��_�H?uv?�o>�l3��{���79�n^b?��?�������><6?-�>�%�_-��������* {>�V,>č��l��������0��D�= ��>�.K>1���s���T�>N�ھ�<:��E�8��D�g�:��<m�>z�*q�=�?(>h�=Q�9�d�����[�@�}?9?gm�?�#Z?�B?m������x~]�s�ؽ�n�>V>�>�k>���P@�>��?�oǾ U���׾{�&?���?u��?IR?�7_���ҿ![����帾�k�=O��<�=]�/�&P�<ݣj�|5��X��C0>U��>\$�>þ�>;9>��>�2>)���T*��즿rx�L�5��#�����R�A�B��Ͷ��������L�����Z=?��Q1����������7�	 ����>��?���>G� >�j�<��F�<Ͼ�<�x�=�����e���&�5G8���5�ָ���쾈P���|���w�OϨ����>�`m�h�=���>�Ʋ=��l>1��>X�C>�L�=@#�=�q=K6�=T#>�d>La;>�,�>�ر>tH{>b��=�愿�����9���R���;�C?�,]�<���T�3�r߾P���T�>Q�?02T>�R'�Y����x���>��D�O:a���˽M} �߉>Z��>�c�=ڻ���yy����5^�=f�>�>q���G��,�8b�=6��>�����=�>8�?�6�?h�
?���=,O�>�R>Je�>��=W�|>"9>��>+!?;?!?��?��>� �=G�����>��@>A�,�|���a�S�\��_=�s�uw+�P�>^��:�"�>f[>_�=1퍽⶗��2/�� �>�
J?-��>D�>��>.�$��!��\��\��>�01�&?�?�A�>?'?��?%��>G|>�ξn$��>�o>p�+��7k���Iu�=Ι�>�H?4�=?g�{>��-�n9>Q <B�Z>��>R�<?�?�V�>��<]/��:��f=��Xھ��o��d���4���~M��{����۵��G	b��C\='r�>���>A7�>���>s:>/�=ħ�>Y�[>q��=��>Ф�A��=��=4�=��#>�=�_$>�U=��ֽ�����cv��
��f <>Py�=�E�]?�'?��1�D��"�J�7������>�}
?��?@0?zS=�����-��=���=��"?�c?<&�>k.��U�=�XE��:����>֮�>�Si>����sL���O��ͽ(�>x�5?{�>2���W�gs�PQ'����>�Y��X½|��?[FJ?5zܾ�ڽ���%�	�F����X��3��@����{ ��d���_�ڐ �r�5�(���Μ�=h�>* �?~�O�=ő���!���4�P&k���=[z�<�r�>~N�=�bD��g��g�O澀+?��==A�>�tB>���>��? 1?��o?��
?f=?�ʽ�9
?��>hԳ>��>P)?>�?p-?�,?=(?��i�<�ڼ�ҽ�˛�*�����H=A�>�F>�f�=�g=&�>u��`��<��V�d\��&�>���=cG�=z�0>��w>8#�=��?�20?��=�!���>.j7�YX�>	� ?n~�>���>O����3��T0�>:�'??�Z?��&?�M�>�����Ͷ�R	Ⱦ����m��>�=?���>4ʰ=��0=��
��=;Z�>�A.�Cڱ��_/��F���Kd�ϡW�yxi>�LL>c	�>��>�ɀ?N\;?ˋS?ZL>>'?�������$�Y��E������>)ժ=�$a��B��n�����e��H�0$��������>�͙;��<nj>�=�e�=m�=���t=�Θ'>�x=Hh�>��?�?�a�=�+>�R��ۗ�wI?�]B��#��Ĺ��p���
�)$ >o��>^*=��?��7<tup�`ͥ�*c!����>��?Q��?Agj?�R�r�޽Ufa>�)>�_�<	�<�V+��n_<���GV>��=> �w��S��'�>=F>"��>6d��hϾ���)n,<"{���k�}錽)v��ے������&�����������b���tG�*�ld������	�K����8�X�!���?W�?@
�>ch��C���i�O�ΖB�����]Y��ͳ߾��=�ž��ƾ�i��1!�"�p���X���8��|�>����	������J&���g�^_�>��s?�	Q�y~��������>�m>���C%ھ~	���N���à=dvr?��X?k�	�r��U�N�=��]?��?�Ԡ>I������w{?T�2?C׀?��>�$����.᜽̳?-�?PY? ʽVш�nGP����hYS?~A?ڬ^>�Ӳ���|>�i!?e C?���=���Q���	���gm?N,v?�m�2�>@H?��>��>/dX�WVO�G����(�i��=TI��=�R��s�h�o;��/�>I�>W婾]6¾j��>���;�N���H�N���R��;�</s?"e�\�>W�h>g�>i�(�����Ɖ��f�תL?��?�S?SQ8?�}��:��<=��b��=�*�>@ì>��=�}���>dC�>zC�xtr�/��ȫ?�E�?0��?4Z?:�m������:��(�� ���&{>�6>X>®�4���J/�<�2>w�j:��<_��>�� >���>W�>��>�N>�u���o'�O����_��R��H9�L�'�� �=8�(���F��c����W�E���G���G�r�
F���.��B=>�>H�>?f�>�By>}>v(x�|)վ����{����,2������v(̾<�R��MW��Si��AM��Q��S���-�>����[I>
?���I+�=lD�>��=Vs�>7�>�v�<g�P>I�>�T�>�D�>R!>X�a�s·>�_t=h<��Sև�&pO�n�<��=�Q?֮O��(����.�ʾ�o��@�>�e?�
A>��,��?��*�g�'�>���lp����� ��G�>F��>*��=�}I�8��8���eнX�f=t�>;#D>�����a���w���=U4?27���;���X>5?պ�?��?o,��F?_��>-�>��>5��=Ds�>�>�V!?Y?J��> ��>*��>T-��z<4=���=��0��'=(A��'<���i=�X�>�A��r*>[qN<L�g��t"��7��`)-=�~��ȃ=��>Y�D?F3?���>d	���FE�6����=��>�W�>��$?�y�>��>N~�>�޷>�Ww>
ԋ>��3��� ��>�O*>�x�����߾ �>�?�$�?��Z?u���;�+�=d�罾��>9?�p?綬>��?�;|>s���gӿK���#��@�=�ؽ2T�$U>���h麻6о�?���w��m_=m}>�=
{�=1l:=�_)<�h�>�2>��=�
>����{����[=�ߺ�☼�s;=8�D�=7<x��>Ћ�=~<�=_7ٽ��j<,�A���}?r%?YO��ƽ�u`����/�����?���>
k�>G?��w=J���:����;���?
x?2-?��>��?�=�K���'r�u��>zp�>��1>[G��K[�>H��x���]�>`Z4?d��>�}���J�r�}����	��>��
��E�Ъ�?��P?kų�QԺ�ӃI��3A�9$�T�)>��V��e���]���F:��mU��������e쾉�Ľ���>���?��=ʻ`>�p�b���Pb����U����M��t�>a��=(	?����=�3�>���w�0�K���>J#S>���>Vs?�3?�i?^?J��>�6R��?��=v�?F�>�o�>�\?��#?1?q?w��^�Qɽk����Q����ҽ�{C=��>�o�=�\���=y y=G�>+�=M�>���=w����p=��C>��U>�"�=b�
?j$?�v��8�
���ռ�_��E�<db�=��U>Y�+��-X�v�ѻ�U>��>u�,?Q��>���=�Y޾�������u�=�a?��1?� �>�h1�.ޖ=HT���{��Y�=�LW>�~j������޾����������>3%�>^��=�>�g�?:�M?JfR?���=��3�/�t�H@�0��=
mɾ�>I��=.6ս��F�L�J����'�-�<��7"���M�$�m>"�>x<�=K@\>ZpĽ�1�=��>y6���=�<<��<��?��i�>�H�>�8?�~�>�4>Vۥ��/"�;RH?I�"�I�	�����ξ/,=����=���>��=�> �=%C}�񖥿����Q?�u�?�L�?���?h':��z߽&�m>��=͸�.-�=�9=�g�-����=��=Z��=�qj�W#��*��=�k]> ��>���p���XdʾI*>�\����D��ō�̓���Z���_��|ܾ�u3�[��=�Bɾ���xA>%��=X������[z���ھ������?Z�?:��>�$�=0�
�A��������|½���k�=�T��K=���"�a�Ǿ9��
ʾ��	���(�%�{��>v����i�����C�q���%>ѓ?շR?�
�=���DY��x�> �o>�P>9-��ǈ������@>�hz?j�?����=0�퇝<Ms�>v?�s�>�"=��\ƾ}��� >�.�>�#�>b��=!<��n���K*��4�?	Z�?��D?����U\�G6+�^>�q?[[d?l��=�ս&z��]��_�H?uv?�o>�l3��{���79�n^b?��?�������><6?-�>�%�_-��������* {>�V,>č��l��������0��D�= ��>�.K>1���s����>��� WN��oG�������;�<r�?IU󾿤>�Va>��
>��'��ό��ȉ�v0�0�K?�-�?�T?�E7?[��CN�ڕ��P��=G��>_ۦ>6�=�	�ȡ>���>��辙Qr�N��b?Dl�?\w�?�DY?��l���ؿ]ʩ��~ξ�]���z�<�S�=��h>ZC��!��AC<=�["�:��l>���>q6;>e(�>�_*>��>�[4>3W��f #�<)��!���x�@����Eپub��NݾN1���:�f�վ|Z���?=�>�F��=.N[�Q'�N�=�@e�p�W>��>���>�V�>�Ӹ=֏(=��� Q���/A�v?��!0�KH ��u��������B�A����@�������a6�5�&��
?r��<�/�=H��>4���5�>?�<�>qC�>5?!>��1�4��>#�>�p�>�9�>g%>���<��z>;҈=ℿU����q:��DS�Z��;�:C?��^��p���3�i�������>1P?l�S>.�'��锿�y�u��>rD��b�r�̽�!����>`T�>�~�=��лO|�s�x�Al�|��=�p�>��	>
8��� ��x�j��=Q��>��ʾ�G>U�>ۼ-??�c?�z�>.=��>�^>���>
�>�Ż�}�>G��>E�?��L?pv?�>��>��J��T�=?�j��?���, ='T{���L�E����̽ǟ��kT>���<r���Q�(<&&;��|-�V&\=���0D�>�[?x�?�`�>�0��9��.8�ET�=�q�>�(>J�?~7�>Q�>�S�>�?�S�>�R>����h,��v�>  G>(�M�!x���ձ���H� >.�t?ʥ6?�t��2�z���"=,��=�O�=-� ?��\?:��>�KV>?���
��6ؿ	|I��Q�q�������r>���C���y>a7����/p>Ϻ�>7��>���>�Z@>��T>�w>[[�>ോ>VZ�=�d�=�\<����,��`3�=v�ʽ���.�=ޏ�-���q޽8��)�1�z/=~��b��?�C?��N<\j0����|� �����.�>��?ld�>�>�E�>aG�ϰP��P/�m���>UZW?^t?K�v�$�=6Q�[�y=��>�Rn>E��>�ւ�Ѿ��þɨ��X�>Cu8?9t�> }m��D4���h�Pk��>�>��ǽ���'�? O?�!����о�A<���X�IEW���Y>:�A��w��Z����)�5�I�e�
���?������P��>X�?�&����RY������/N�2ig�(D<o[o>H�>�0>$ ����ﾬH4�v��1�ZM�=�_�>=��>JΣ>>��>�'>?EDy?�!'? {�>*�B�$m�>V���ë�>��?�>G6*?��?G�>C-?T�㽫�7��3���9�^3�����<O�T<�Z>��%>���=qK"���=����6=���=��=�~�=R���`
>��
>i^�=#�?��?�<�`��=��<�2󽵄�={�>>�)�>f���?YL<>���>�?�5?�?�_u>�d��d#���m��;=$��>�}E?z ?Rާ>+�>
��g��d���`�=������>B�[~��L�y���S>��>��<~2f>%	~?*�G?E)?��g>�x���������jf�����=�i>��0�o�\��I���6�e�����i��� ����=I<�=�~Q>*V�>���9%@�=k�<��>����,>:S,= a�>o��>@�>�ь>q��=�|������1H?{c�����������;�O0�w��=��\>ã����?J��)*w�龦�;[<����>WD�?$-�?��a?�E����P�P>h#A>?��=������6����������,>씚=l3���a��j�=��D>�#R>!%��i�Ӿ������#�J��%)�����kd��Vw��̪�Oho�Mz��[b�ߴ,��-����<⽢Bֽ�����0�������H@�?���?���>��=i�(����m%�Nr�cɣ<{�`�M�:�c��� ��
꾠M
���u�I�����M��m�>R�����7��Χt����=�`�>��x?�y�v񾽆9�q>$�=U�J<�ھ��������Z�>�k?[�G?��!�\vO��=)a>��[?�?��>��3� _��su�>:|$?E4?IB�<[NC��vg���;>t��?�Ǵ?�`7?����SN�?g��Ҿ�2??�U?�X7>1tD���ɪ���>�	?Fj�=�@u�sd�����X\f?��?�߮��k�>N!?і�>)�\��(��� U�epӾ,�&=���=nd��t�7��3.��������;P��>Y�>wfR�7(��)�ܽ����P��:IP�sU�����>����>�F���9?߃���'����a�����sM�Kˎ>[��?�q�?���>+��?p��)�]�:�g��$�<h�?�kA?}'0�
	�]h�>���>k,T����a{�4��>+��?!m�?R�>rN�:Gӿ
��������9��=D%�=��>>��޽Iʭ=��K=Ř�Y=�c�>]��>�o>�:x>D�T>ݛ<>��.>g�����#��ʤ�.ْ��[B�� ���wg��{	��y�����ȴ���󖨽���-Г�J�G�?���T>����ރ>��#?��>��>��=�����K�e���V�*��?�*�X���쾾�ܾA�i�v����Kd�牾y�޽2aξ��?4����{=
��=e`����<�?�=���=(2G>p�Q>w�=��=���!�!>A>Hӡ>h��>�ɂ>��G=���)`}���2��VM�?����c>?TV�o쏾��3��o�<���7�>� ?�bc>�"�9���WZq��h�>�9/��R�li���9�T�>b�>�*�=s��;��ּfe���i�� >*�><� >D1�0���w�Lp�=1��>K�Ծ9k>��M>�=3?�,k?�H-?+[�<l8�>�r>U �>��V=<�1>}�O>bm�>�^?�#3?��0?{��>��=�qT�Nz= �u=�aK��9���t��Q1�u��S�<s��lt=f�=B��<�+k=|ȴ=R:;n#C<;9,=�5�>�
?���>��>�T�=	M��#	%������ؾ������=�F�\�>[�H?�C'?�L?�'>�{�K��=�Ï>�ó>��J�V�#�=��=T��=enE�I��?�J@?��ݾPI"�=�>h���Q��>?P�C?���>Pu����v�1��bKȿ0����@�h��?��?���謽��M<����m�7�^�����a�<&W=���=Z��=��<�$v>��>B�=�.3>;V"��j5���@=�� =F�=Y:��~��=��O�:'+���J:���('-�����
�}���ٖ�ZE&?3��>����-�A�����澨�<��,?x�>�7�>�<J?n��>3'Ͼ<g�衁�aXE�/�>i��?�?o�L=?�T������as��[�>�?�br>�TC=Ik��뭾�8�>�M?!T?V�>r)Q�^�O�t:v�^��2?s�@=�������?oR?�2��yX���a��]B����+�T=}\�v�V �����?�2�F�!~���>�b0�=$��>���?�τ��x�=l ۾�ꚿ8ip��?��J?���7=���>�lb>�3��G|���C���J��:�<��>�V��{J?̆	?��>\$?QN*??W�>1o~�$�7?�8���(?��>��?��=[�H>~i�������l�=ȫǾ�?v�mɾɵ=�n���aY���b;¤�=3	�6�n���=Q�=�7J�'���ܘ=B����=��=�f>N:>�*�>*��>q@�������>k�Z�0ĳ�M&�=�"e>.68�I�Z�D ����W��n{>�,?��?:�>E��A�!�0��4>B�?HB?�5H>.=C�r� /ľ�;;��=��>��O�B����߾�+%�W]��Լ�>�)�>�,o�2�5>q�?��?�t?���#�����*�S��3�`>sD����>��>{�>zW�U]-���g�Y_�>7�U��A����0�>څ>B�=��>��=]k�=�^
>�b�'L��؆�ϒ��n�>��n>?��>p��=�g:Wd|��u��^<?�.8���}�J���&{S�r�
>��>�Bi��u���$F?ii��[�]G����ɾfA?e�?Aj�?��>�(���=����B�Ѽ���>���=g�B���v�����1f>Q9�=(��H���P>�N$?���>k����^%�!��ۼS�� п�V[�1(�=����Z��v~뾾�Qӽ�S��9��
[	�kBM�d���&�N��{���j��4I��J���������?T�?d@�><��<��+�h�/����"ּ@+����R=.��	}�]Q���$Ͼ�Hb����������He������>��׾���hS�e�:�@>̒�>$��>����O���W���d=��>闉>�q��ؼr�Ա���4��`?�m?<���ߡ�����wo(�K�'?��>�u�=�{B���w�]�@�S?G�y?:�>����ӝ�Y�����?���?�_?B*־hNh�?�d97�(!V?��?R��>T-	<�~<�N��I?��?P�?\�����5Wr�#��>��l?o1����>
'�>��'>��[�f��0��q��KU��ֽ$>���_�ԩg�1���(�d>���>�M>����=��p>Tr��kٝ�j�7�D�F��̏���,�g�6>#�#�?��=
O�|�%�9������N�j�<��j?�i�?��D?�[?���h��\�y>�e6�{$v>�?�$��Ž��>��>;�ھL�d����A�,?��?a�?�_?FV�3sѿ����+_�˅������ˁ=���>ˮ ���=��>�$�<}�<���=Mg>3�B>�R>��=G��=���=�܂��1��L���͉��@N���'����}��v1��A@���)��/����ݾq�ǽ�ʽ	׼?���z
�)~ļB1�  8>�1?M��>�ܰ>j�>����:�׽�Ⱦ�j�㱌����&��ݕ����ľ!*����
=��� �8��1���;����	?��������~W�>Jb�m�|>cN>������>`�m={��&"=o�m<[e�=�=�=�U>oz2>)�}>LpL=�_��SZ�ّ3��BI��ZC<��??�Z�"y����0��9㾉g�����>5�?D�]>)�#�����#gw�?�>��m���X�������oU�>���>嚽=�0;�l(�7p��u����=嶆>W�>�p��)��d��S�=��>CK߾�"9>E&>�j*?7k?CM?��=w�>�P�>aK>[;�<]ZI>hK.>�>}B?=�7?�6?�I?F�=I�S��A�=�7�=�	@������	��m��`�l�F=Ѽ�=(��;�Y;�kּ8�@�*5-��aY��И�������>�C?�_�>*�>ua=Ϥ����m��{νE��>�ӾZ!�>����X>�$?yu1?�c(?1�>�F��Է�a�>.��>s?B��N�&ָ>�a~=QZ�<N0}?��6?�~���D@�� f>�Y3=U�=�s?�?"ɑ>���'��%������*��1��󈾡E�Q#��{��X�=���=�0 ��*��ܢ����=��>� >fХ<&@�=�0=�H�>�5j>�,=
?2�F�c<��=�OŽ"��=T���Y��٬c�i�Q��A;��*E������aq�=�o��hJ���?7Q?���=�=�<�ӄ�o���F�<�R?N	�>a�>ޢ?�b�>g#���`��^��<u�xF�>PJq?��?�/=��<#��=�s�8>j�?��=�6<�:�=כ��P�>�#?.:@?�@t>��ž�]j�(G������V3?/7P=�X(��%�?$t>?%"�Dx��=[%���E��$��8=�$����	r���U�*���Ծ�žW¢��`,>���>���?G;��,>2�׾���;k��˾k���
���Y��>��+>��[�;�&��ܾ�
6�0c�⌎�=>#wI��EM?���>��?,�A?�5?	�!?�Q���d?�T��R?��>�J�>������=f�1��l���=E�6��罱�~�ʢ=>��E�=���=�H�=��=�!��T����<dNμg�L=�@=��^=���<}'<�4>�U>?�?���>u�����#=�U�>�@���M���>,T=<��=]�O���<X���5>:?�?e��>��j��,ɾ]֣=��?3�F?7ǟ=��>�� >���x��u~T>P9>yi�-�پ�����.ȾX0���>�֝>�8�<3>>�A�?�9"?c�L?w�	�����ܜ:���6��h>�Ӏ�4��>7�>��f=�ؾ�/�U�d�fhF��:N�yj?��m�{#>Ч>��=c	?>>��Ŭ=�n�=:�b=��i#>;�����>9��>�g ?�M*>��`=Z`h�i̾�~-?�h��Q�$�ja��w�l]�걞>=� ������X?�=ľJ��� ��A����A?J�?]$�?���>�'��@�>2��H4��/�.>���>V�Z==CG>�ݽD�q>C��>�>O˜����=}`G?�A?��������r��ZſG�/��pA�W(J���辁���ð���={��}4$�D���͉�xw��8�O{	�� �:.{�Xپh�Qs�?�|�?���>��=b��20�M(1�����c���P3�|.�/n���k��w0پ���y�ɾbӶ�z�V���/�>�f ����"����X>�A?Ԅ>�����=o�;��O���>X?�M��V�k����AZ�5f]?2j ?�4�ҭ�g��=��o�V7�>��>M��> ~������DϽ��?�8�?��ݽڰ���P���',��9�?�Գ?��T?��ھ�~t��nھ�[ �� ?���>��Q>��U�w(Y�U�d���_?�v�?�?'���$��R�e���>��`?�������>���>i�I=�q�=A��JgE�[�ܾ�둾b5>u}��c���f�� x�f�=>���>Kw�>�r���	�)�ܽ����P��:IP�sU�����>����>�F���9?߃���'����a�����sM�Kˎ>[��?�q�?���>+��?p��)�]�:�g��$�<h�?�kA?}'0�
	�]h�>���>k,T����a{�4��>+��?!m�?R�>rN�:Gӿ
��������9��=D%�=��>>��޽Iʭ=��K=Ř�Y=�c�>]��>�o>�:x>D�T>ݛ<>��.>g�����#��ʤ�.ْ��[B�� ���wg��{	��y�����ȴ���󖨽���-Г�J�G�?���T>����ރ>��#?��>��>��=�����K�e���V�*��?�*�X���쾾�ܾA�i�v����Kd�牾y�޽2aξ��?4����{=
��=e`����<�?�=���=(2G>p�Q>w�=��=���!�!>A>Hӡ>h��>�ɂ>��G=���)`}���2��VM�?����c>?TV�o쏾��3��o�<���7�>� ?�bc>�"�9���WZq��h�>�9/��R�li���9�T�>b�>�*�=s��;��ּfe���i�� >*�><� >D1�0���w�Lp�=1��>K�Ծ9k>��M>�=3?�,k?�H-?+[�<l8�>�r>U �>��V=<�1>}�O>bm�>�^?�#3?��0?{��>��=�qT�Nz= �u=�aK��9���t��Q1�u��S�<s��lt=f�=B��<�+k=|ȴ=R:;n#C<;9,=�5�>�
?���>��>�T�=	M��#	%������ؾ������=�F�\�>[�H?�C'?�L?�'>�{�K��=�Ï>�ó>��J�V�#�=��=T��=enE�I��?�J@?��ݾPI"�=�>h���Q��>?P�C?���>Pu����v�1��bKȿ0����@�h��?��?���謽��M<����m�7�^�����a�<&W=���=Z��=��<�$v>��>B�=�.3>;V"��j5���@=�� =F�=Y:��~��=��O�:'+���J:���('-�����
�}���ٖ�ZE&?3��>����-�A�����澨�<��,?x�>�7�>�<J?n��>3'Ͼ<g�衁�aXE�/�>i��?�?o�L=?�T������as��[�>�?�br>�TC=Ik��뭾�8�>�M?!T?V�>r)Q�^�O�t:v�^��2?s�@=�������?oR?�2��yX���a��]B����+�T=}\�v�V �����?�2�F�!~���>�b0�=$��>���?�τ��x�=l ۾�ꚿ8ip��?��J?���7=���>�lb>�3��G|���C���J��:�<��>�V��{J?̆	?��>\$?QN*??W�>1o~�$�7?�8���(?��>��?��=[�H>~i�������l�=ȫǾ�?v�mɾɵ=�n���aY���b;¤�=3	�6�n���=Q�=�7J�'���ܘ=B����=��=�f>N:>�*�>*��>q@�������>k�Z�0ĳ�M&�=�"e>.68�I�Z�D ����W��n{>�,?��?:�>E��A�!�0��4>B�?HB?�5H>.=C�r� /ľ�;;��=��>��O�B����߾�+%�W]��Լ�>�)�>�,o�2�5>q�?��?�t?���#�����*�S��3�`>sD����>��>{�>zW�U]-���g�Y_�>7�U��A����0�>څ>B�=��>��=]k�=�^
>�b�'L��؆�ϒ��n�>��n>?��>p��=�g:Wd|��u��^<?�.8���}�J���&{S�r�
>��>�Bi��u���$F?ii��[�]G����ɾfA?e�?Aj�?��>�(���=����B�Ѽ���>���=g�B���v�����1f>Q9�=(��H���P>�N$?���>k����^%�!��ۼS�� п�V[�1(�=����Z��v~뾾�Qӽ�S��9��
[	�kBM�d���&�N��{���j��4I��J���������?T�?d@�><��<��+�h�/����"ּ@+����R=.��	}�]Q���$Ͼ�Hb����������He������>��׾���hS�e�:�@>̒�>$��>����O���W���d=��>闉>�q��ؼr�Ա���4��`?�m?<���ߡ�����wo(�K�'?��>�u�=�{B���w�]�@�S?G�y?:�>����ӝ�Y�����?���?�_?B*־hNh�?�d97�(!V?��?R��>T-	<�~<�N��I?��?P�?\�����5Wr�#��>��l?o1����>
'�>��'>��[�f��0��q��KU��ֽ$>���_�ԩg�1���(�d>���>�M>����=� .4>.�ξ=��{J���J�����~=Cy�>�?)��5?�#�;�*\=�W�&B��X������L_?���?��3?V?x�'�����#����;T�?k�V?��ν�O����>�u�>J�^���U�����p�>��?� �?�pR?/d�ڿ�e��C;��y��'�=�(>3�L>�I���u=�=��^<�C"�KO >��>�&S>B�.>�>�>/Z=O���2(�6��������.��t�5n��F~�B����®ʾ��Ѿlf@��!���ؽ�n��~	�,gؽ$Dc��/
>?��m>"��>,>�a�=$d��P�ľ�� �?B��� �B��)�ɾ⢾�kY��n�F0��1�wڽ�対��>���=�0�;,k�>�ܽ㈮=��q>��>٬�>��&>	��=}M�=o��=m�%>"#!>�6Q>f=�o�>��=d?���#|�.���H��[�;v�6?��g�4E��{�2�������Tl�>��?��_>5�#��+��ϰl�<��>P�8��uE�{�޽3~��Z�>z&�>i��=�I�<1��Y?�������>���>%P�=�>R����6�����=L\�>�7;*z>.�>$�,?]h?��$?+,f=2��>�Zu>ڮX>���;�*>ۺL>$6�>0?�N*?S,?0��>�\�=��,�ޟ2=)U�=�P��v�<����8���v�=��=�[.=�vE=����&Z=��==�|�^=K�;9��>t2?��>��>��=:�3b���o��
K��B����>z��="�]>��>P�?# �>�V>�i�t����>��d>�6��m`�e��=��>ua��{8?b'?�l��\���R>Hޅ<Ҏ�=>2;?n�>�*�V׶�����ӿG$ʾ�J/�n����-d=��<�v��y���j�9�w����"�a��~H>�q>(Pr>�$>Z��=���1��>��=>Ak�>�&�<�H~�Xn��5�����=ʼ�t(>k���A;W����%z�+M��d��=֪޼�u=3�,>�L ?�?�O7>���<],!�q�d�jٟ��OQ?yB�>�$�>{@?�N<�N�_xp�C�n�}9�fO1?'Uo?�>>�h��B�{�X����=c?>��9>@��>�Ix>5h����7����>o)#?�??-�>Ux4�?yE��V��Z���E�>yV=7�ӽ���?�J?-a���e�����H�:�����·=���7Ɖ�����;����0�Z�����'�/c	>z��>�"�?t���{$>d�Ѿ�w���px�S�����y���<ܦ�>O�.>e9��刾�{����^ �A�=��z>��+�@o)?8O%?�3?�8?�>H?9��>��a�DU8?	���?8�>��?�t>Y��>�1����F�˾7���8��@�G9��R�*=��H���=Xs>و���O'=G�2=���=e��=[��l}�;%��ش=���:�[=`�d>+׾�s��>��>�.ؽ�>��o>�=P��$�@�8���<�k����3*���>g��>/�?�r�>9A�<�;��%Jξ\�ھ�җ>�P?��>�*�>��(�	T�<|����>}��=S>*������_��ڂ	�������>z��>��=��A>R�u?z?�ht?��/�������N��*>�I�S��>���>y��=xw���J�gc�Z�ډn��K#������r�>�q>��?>�>�D>4�G=b�
>�<������=o.�=�E�>nv�>i�?�}�=K��=-�z��w�E?�y���r����#�^H�<�I>��]��iƾ�<?�VQ��_��`���I��?<��?��?��?�b4�y�=	��=�G=��g>r�B>�z���2��ܽ�A<>#���螉��#��>�7?Y)8?���H5��B*���/>�̿�B�]�>��Ⱦ�t����Ӿ�F��N%�Ί���P����v�J�5P���Jv�Rf����R�L+��Kw|��(�?	�?��?T�^>��6��
#�I�;�J��B��ܾ[��=��� $��߄�����~��P��~���?��5��v�>�~¾����a\b���Nh3<�X>���>,`ؾ��=���&���.Ĉ>N�>&I]�v�f������T���p?ʰ"?jk˾�=���g4�@��<�w?^^�>-�=�3�ʋ����z=�V*?��l?~[�<`��Z0���s>���?Ȩ�?.W?�7����a�)��:�áI?r�?���>��\�`�0��t��;?S�?��?iy���r��j��M�7vw?[m;��>>ܽ�>R�->�Y���W�E������f@���A�o$徂�%��|���#�y>���>�)�=9v����Nh'>�sž�C���BQ�-�N�a��D��V��>}�U�V?	�)�-�����i��w�����tA=s�z?���?X?C.�?t�(�X�|�J�{��vɽ��,?1R?�D��o?���>˼=�,���;��m罼j-?Jr�?���?R`?Y�9��pܿq#��ȩ���ž_@�=1D�=A��>b:Խ�]=�eR=R�<w1���"�==
�>��y>�p�>u|9>�	;>7>�c���%�!��_���J�C��H��z�=�-���q`x�����ݭ�GV��56����r2��C�F�Ա �ˌ*��	����>�??{?�|_>�0	�:t�=���R�!���
��Q���� ��p��J��N�z����d=�U��Rx_�#�-�ʫ��_��>,�d���B>��>.���h �>��N>zj��?��J>�]B=<>��>Y�<�d�>2�==���#G�>��e=�񅿁�~�<�4�%I�#�;�>?�?^��T��.1�k������wo�>�C
?�W>0�&�`ޕ�!w�
��>[�`�t�X�R��Y&�ڗ�>���>A��=��;6F<�g�{��������=���>�I>|���䑾������=���>�#��p��=�{#>��)?v�h?�_?��=��>�w>�-~>�=��P>�2>�i>���>�*?{h3?���>ej�=�,��i�=E��=�V*�)�̽�\�3���}��MH���h��<&\=�P�;]J <|�d=�z_���J=��1=�@�>iV8?���>�"�>�@�=^�E�U$I�!���1�<���W�>k�>�2�>6X�>VC�>���>�*">�xp��S��q�>yf�=�I��g��L`<Xi >���=��9?��4?�Ӽ.�M�<h&=��j="2B>�D�>�*?� �>��=�ز���N˿�,��W(�����*<�����)>�<�<h�U����<�r�#+=�R�>z�>�H'>�=Z;��=���=���>��>�?�=Pۤ=�S'���ѽeJ�=|o=�	�\�a�����Ⱥt���=�����:���������=��?���>���=��ڽ��`kH�l���L.?�{�=C�?9�?���;e���|F��f��{���j?a#S??��	����U��p��Aѳ>*B�>�N=R(=M*�րu�:V�¦4?�%?�vE>҇i�i�i�Γ����Qg?�.�����j�?��O?������W�9����%��}>��ɼߕ���a5�ԏT��}�Z֞�R���/�=ս?=p�?�>�;�=H0�������X���_��b;�>�>��>eX>kF`��yվ%�aIоjVc�+@B>�_A>�	��NI?�;
?��>�%?�b?��>�U=yt:?~@����8?���>c-�>�U�2��>�p��:*��+�:�0�p~��4Ծט�=z}2�����	>�g�<T�=e�{<�=E%=>��*�<�U&=��=�=�š=� U>#m�=�?n3 ?�����98=Di�>*i�Y��=��̽��=J�
����}�f��=d��>���>RK�>\B�<Ѣ������"k�y�>r��>��?��=C�9�C������+�=���� �=� |�!Ҿ�N�}�����=�W�>�x�>G�=��C>�G�?L�?)�\?��D�"i�o5��-�q@>ʯD��۝>O+�>�޳=F�ԾAJ*���d���W�uVU�0;ؽ_ί�pȆ>�F�=�O�<BÛ>O>4۫=�2�=$���͆�Axn=�0=��>�l�>-�?�>�K�=I%꽷�Ͼ�'8?e��"7�
���D���:��C>�
k�0K�JT?/���o���͜��C�)
4?@3�?MG�?�1?pf�\#>h�[�#��<I2�>ư�=D�R�(���?���j>�_>B�=��پS�v>N�?!N�>�L��� ��L�v̮=W�ÿicH����;ǎǾ�E����Ծp4��,�ɽ�♾��޼��P�7���3�(����"6z�k߈�da>��H�?⩗?�z�> �K<����?+��W�����˾���<J/ھ�0v�����1��
�b��p���5���Z{�cf�>�\徰���?(�٘���[	=��>��f>wڱ��/�I>�i
a���>��>�1�-P�7�����I�7Ah?��?�E��{����;a��=�d? b�>���<�^�<�z���=�X?�G�?n��=<ɨ�����|�׽D�?>��?/S?p��"m��w��ϒK>�?�X�>�&>�R>,����A�V�l?5އ?6�:?������t�H���I>@�7?�������>&�>4��=$W��+�c�>)�;�e�D���>&I`�摀�[����͊<�4(>�
�>a�k>3�Ǿc�����>5k��)��j`��������p=-~:?���MP>9��>�;>��G�����Se�^�Q��a?���?Ċb?kr?O�$�
;e��Ӝ�Q��<7c6?�U?�@=>�r��G>FG�>�wӾ٦]��<Ѿ�M,?�?E��?�s?�|e�h�п�?��:���tʝ���1>�>�MT>&u�צ�=�6.=�a=�j<��8>A�>�z>��~>t,a>%Q>	�>>z����%�8ݤ��q���5=�##���Q�~��P�����Z���Q弾/����Rq��E���C�j��y�;�&r�[��>f�\>R�>���>E�>�}�=�F����:��x����Ѿާ4�F�Ͼ,�ξ�ߨ�U�ɽ6�W���Ľ�Ҹ��=��ɤ�0�?��ɽZ�4>�^>g|<�XJ>B�>J�
>�>>ޡ����=���;a�,>�&�>�̌>�+�=��>��"��g��5����0�ϋ��9=��F?��%�Mܡ���2�x�"��N��>mC?#qy>"�%�����/.i��r�>��6��K����ӕ���W�>aH�>��=��y��b��v���r��2�G>r�>!�>9�2������=[#�>'�;B��=Wkf>�D*?��s?�_.?��=5M�>q�T>�sc>/P�=$�>��A>�]�>J�?�o5?P,?���>G��=@bP�J8�=�i=�zJ������ƽ��/7/�cj�@[��KF=��\=5=R<$f;=i9*=�3����<:h=�6?�`A?�S�>�l�>�h�~DR��a�*CQ>+��>H%���?�?26�>%ο>;Q/>5\w<d����Ͼ�g��-�>b�R>6�l��%����>K�>��}>CD>?z�P?E.s�r* �C�>oه=U[�>G�?)�;?�>q���)����A�:Iп�Z�X��TnV��м(v��6h���K��S�<��ڽ�i߽�=�=�c>�f�>~�w>uTL>�/>Q->��>aR�>2N�=�)�=��,��}���ս��
=ơ{����<���A���Y�?�ñ��>�X��������[T���ԣ�]T�>UP,?+� >�F=�g)��㹾�M�ر�>�"�>0V�> �Y> �;i�*�J�L�ޒM��d<�J+?�j?c��>��N�o=�%���`�>��5>}�m>X_�>H�+�H�n�����I><�"?��)?�pD>�g��=~p�j������+>Ȫ;�|���k�?�Ui?���鿠��~�h�A�ZP	�ք[>5��=St��y햾��$�ՊE��T&�u%��y��j�=j$�>BI�?��F�����aھnO��f#��:kg��+M>h��?x�5>��A�����NW	�5�����1� >�s�>�l�=��>Ŀ?d%?��L?o
?()?p_Q�C?C|B>T��>�D�>i ?%��>g�>�v\>I�t>���q�����1֕�[��=Q�;-0	=��>'!<>��׼�tB�ֺ�=�=CÉ�b;�;�U�<��*;_聻uП=��$>`6>Ѝ?��?Y`���S���-����F�<�����>�eֽO�ܾ�z�=_c>���>I��>+�>K�-;��n#�R���W�>�N�>�U?gE?E�g=R��s��V�ľo@�>���>�҂�9�~�\���H������.��>�a,>�>��@>
�q?9J?�G?����#�1�L�	�!��sG�=���>�D�>*��=���'�@��v��]��%�||���A��%D��=��C=�k>S�;�I�=���=QBüD����=��=�M�>��>i��>
M>�	��;����2쾭�Z?�e�QV4����7Hm��>j�s>��>�R�a ?��ཨh��������n?]��?P�?@j?[6�`����v=/â=0��=/a�=J=1��}���'s>8�=]�Ǿ��վ@��>6`?��>�`���sX	�{BU=�п|�;���="��z�����!��侾㈾�i�MH�=���PB��,���0����=߱��q]F�����y�?��?�0j?	v�>;�l�u-�C�X0����;>7���\h&��^�GP�����Fþ�>̾�L-��d���"�94׾PՉ>����΄��{�v���C���D>�k*?&���ҟ�"������<�l:>��=i����c��4ӏ���%X?�Y3?
?޾���t�Bg�=`�?L��>��}>���:AI��?7>.�?�+?�޼ᆿ�m��@�˼eT�?�6�?_[?B���(b�D�0�v5�Q
(?AQ?&��>��S�'� �����>D�?YJ?��+��G��%�R5?�5h?*���"�>�Q�>Q�>�eþ�T��$ہ=u����X�G�]>����_�8�^�{>��yz�鈁>���>T��߄���>���(��*o��/��}P�_���+?d���<?V=>_�Ļl]w��p��R�o�8V��e�l?k�?��A?�p?~�J�M���������?��>6l�>��=AF�>�5�>�B��v�z��C��3X?z��?�d�?�'�?3/��Կf���F���#���n>�_>�b>�T��	 >���<h�i=�2=(>�u�>�a>��>H�u>!��>��T>�t��W�&����Qߘ�l!/�����~	��I�����L�������ٴ��k��I�m<SE켉p���&�����mX"=+�𽐟�>j�>�%�>��>��>3X>b7�"9 �w�M�n�� �O�E-޾�˰��mȾ�6�����o��΢4=.�潄���A?��=�>v>�F'���5>A?���>�>��>g��;%�=�C7�25b>K��>��>�$���>E.�������Ո�`["�-�S?�=a�K?_�������2�*m����S�>�T"?�t�>��'�9���}�^���>\����,�H�Ž��o�ỡ>���>��U=�}=T�*��þ�oν�+u>���>��>KS��žeR���>���>�}ʾ3X�=�I}>�0?���?�KC?��2<_&�>'�>҅<>���<�+M>�h�>'G�>1U
?�o?�?00�>���=�V���i>����s����j��,�~n��-�E�����I���6>t�=ׄ�=�e�=�t޼�~ؼ�ε=�^*=�*�>B?�X�>B��>E��}�a��1��=$>�L�>8]m=a?5�4?���>%�>l��>�A>w����վ�-��Q�>$X�=�X��`s�b�:z��=��>C�t?�%I?`�����y_!>!m:���>�l�>�B?�i�>��V>�Z>�g	�E�ѿ��7������|>C�>��B=#p���3�)���E<��h���+2>36t>�.x>A��>�}�>��M>X�?%�>5>��=;�>��<�o�P�������1�ܢf=�l�<����θ��n�����P���r�Ӝ�|��sͼ(�?P4&?�\t>�#U>�̐�E	پZ�-*~>�9�>��?HJ�>B�=�U)���K�, \�߅��IE?h`q?Ы>3<;�k/^=������=�8�=z�>�Vw>�r��v���흾[�>���>q�?�(>���5�\�y��2	���.>Xs1;]�a�ژ�?��'?������������LV�ZQ�����(�����H���,��-'���%���g��/�}=:��>��?�\�����=�qU��ᕿ�Ԅ���	���L=њƽ�V�>����2��u��l^5�߾�u�=���>e�?h7�=.z�>߸?[�5?��/?�yd>���>E0 ��7?o>o]?�|*?�H?���>�=�>�R�>W߹>��=p~�y���Q��Z����,�M�\>�w>�0�>�8�$Z�,+ͼL&K��8��=�l5;�_��K3�<���6�躿&>J?��?97�}'�=���!@���=���=�V>�E`=	<�WeA>']K>N��>Z?,��>ٿ�=S���x��������>�^?��T?"�??��=�&����p�۾{�=ޮ�>�x��/��,'�2}�X��+�>B��=#Ԡ=
Tl>��t?�Go?Y#?v#�������>��] ��n�=L�F>�i�>/�x>����J�&��x�/���@*f�%V �-P�������M<)�>���;>u�� D=~�_=��ƽ�%���>Ϛ�>�6�>Vҵ>YY�>���==����砾�l��X~_?c�����H�}���.����B=�>��>��w��0?��s�z�n�}w��5})�_?���?���?d�k?��5���z�Q��=d�-=��=��(>�lK>t0>z!4��!�>l��=a��TѾ�_�>i�?�_�>�@�<�$�[�=���!=�8��1�S�N�ս˝���l��]���t���������̭��y&��j5��8o�D���D�꒍��޾��?� ��`�?oi�?�7u>��������$�ib���(����ľ%L"�Pcx�K���n�����GϾ�5�6�-��L��L���>�젾�
��(v��h����=��>��-?��l���@R%����GO>�Ku>�wi�XU|��������IoO?��"?w���ɥ��)׏�õh�s��>��>;��=�_���x��|&=B#.?E?;�=�C���\��aB��Ŷ?���?�;S?�����Y�.1�)�ξ�\'?0P?O�>�ɽ�B����H�>=�g?@;?w��&�_�:`$�g��>��S?N�o�B�>���>�l?c,���ɾ�9�<��^v���-�>�K�6�ݽcx����<	��'�>�t�>����:y���ܣ=�'��M&�:�o���.�0#�����<���>����	�۽rH"=p�>U*x�eJ���}9��|�;<�?���?�e7?�J?BW?��f�x���+��$��=�>�>|�>yE��xp�>Ps�>���N�|�������5?�?�)�?-�N?��j��v���W��ok��衾ڄ3>��=��l>@B��gD#>�f=<�=��H=ԉ�=�u>/�m>��R>���>|>�f�>�Ӂ��"����t��B�^�F�@���������� �����.��:�����?��Z���rv��:��C���sQ�&(���>��l>�6�>۟�>���=��4;�<B��-�Aȱ�x�2����H���h�V�ݾ�$Ѿ3侫0��8?>ۃо��?y��=N��}�j> ��=��>�,�>Γp<��>k�>d~N>��=��<f>^�=��*>�>Z�>@A�<�a��E݁���5��F6��G�<BnD?\C�D�����5�0߾�J���ߏ>[�?�k>�'(�����}s�n��>C"��Q�#�����/�kӔ>�+�>�
�=���<�篽୆�ڷӽ���=y�>E2>	������H����=���>��ҾX��=fw>�O'?��t?14?�.�=���>�=\>׊�>���=p�I>YR>��>�?�7?s�1?���>9P�=U�\��=�ZE=�@�%�N��\���Z��=+�!�<���&O=�_}=-�'<�a=!,R=n���0�m;�
=q$?��*?ӛ�>m�>�Ӿ�IV��L0�\�	>:ߎ>�^J=���>@�?�d?I�>�OY>���=�<�@�¾\�)�n%�>0�$>"�@�P�^�_�a<�i�>�X>@�Q?��B?ڴ���A��=j�<L|�>�$?��2?���>�Z�=�������Ilӿ~$�A�!�#傽3C��Ј;X�<�
�M���74�-����/��<��\>N�>�p>�E>��>5=3>�R�>HG>�؄=u�=��;�;?�E���M=9��G<?�P�w����#Ƽ3�������I���>��4�E-ټ���>�?���<��=kҍ����)��#U�>��E>�@�>��>6D������s�Z�{Y�3[p�q1?	�^?�0?�z.��A�=�n��⡠;h%�>��^>�P�>&EA�v�@�?�����=�?��?B�>tPo��r�9�a�9����>���r����I�?�_?��Qsp����uD��|�4IʼU���|����>�'�G�+�ˢҾ����ʨ\�:{L>l�>=
�?�����U>_�ܾ�薿�1����>��==�x�=�z�>=�=�vu��M������{��;6 =m�A>�>�>C�>�/?K�?��:?r ?�[q>�R��n:?���X6U?�D?�^)?�?�+>��>=��>�A?=Xt�������)��/R�W��<�<z>��;>��	>;ܶ�l�	��S�=�.�<�<%�0�;^g��$g��u����=>�ޛ=��b>��!?�??)���;{����R������=d<>���>N�½�����M>�]>/|?�??r�>�Z������{B�DQ �M�d>� ?qA/?��>o�<j�8��(����q�=M�>��p��z��Q����ɾ�s����>,�m>]�=0��=(|n?�9?BA#?aս0E��XV��o�D3]��Q���>\�>�>z
 ���S������Q���"�=-���>�<��=�6]��ep>�yo=R�}>nQL>�9�P'�:�Hǹ� >?��>�D�>2�>�Z'>���9���b
��V?ںM�˪s���<�ԙ��ּ:C�>�X�>������?��#�Z3q�ر����??��?Y�?�'?�j8�V��==Vq=���y��=s�>u-�>h��=53���f�>�82>�����*�b�>�H?h;?9gd<�_�u�D��a>'˹�)J$��P���褾?��o[t�VؾZNɾt�Ծ��\=!��חϾ����&���	��I����8��^����J�uU?G|�?��\�B��=�
ľ���@�-�$>Mc�oY��8�xϥ�M���h���\�����#��a&�PC�$��>#�ھ�7��a������e>��>��-?��6�����0B�� c���?>��>���	CK��+��ż:�7�r?�?�XT�V����1����T���?��?�2="Ԇ��AϾ=�>�
2?�W?�XU>)E������|���:�?�$�?hHC?�����@O�^'�S�����!?��Y?�X�>�A�m����þ�6�>�E?ԇ4?u_U���Y�(����>7�?�q��T��>�^?b�>��]���˾����>���2&���Oc>Z�N�2��$�|������$����>��>����<깾����H(���þ��9���݂��cN��\3?y���q�>�M/>ioܽ�n_�`���0�P�BmS���a?��?�O?u�z?��*��.����wM�>@$?@¹>�~�>a�=B>��
�0d�!y����[?��?��?O|?����ٿ�s��C<�������f> �>���=����8I=4m=��=�5U���>{�>j�a>B�>��1>~|@>��)>A���#����������_��R-�)/�❚��(�j�G�zV�w��!�;������1r��C���X �樾�S>qHU>���>+�>@>D}R=R��b�@��V��2��j�<�$k��^Ꜿ�K��������־����6�z�9`���Ⱦ�%?�=�ɪ<<A.>���5Y�=VS�>�G<I=�=J��>X���t��=���=���=��+>��[>�˼��~>�֌=̈����}�E�0���8����<��??�f��}�� 3���律3��}��>0�?K�\>��+��k��u�u����>�^��id�Z�㽲�K����>��>�1�=�\<f_�*t���޽>��=Qׇ>Dm>k��&ȋ�ð���	=���>�k���~�=ݽ�>K�+?V�s?�1@?�*>
?}� >�Կ>9	P>qE�>:PA>��>$�>��1?xj9?V�?ֲ�=2����1>ʺ�=�Y���f�c�ҽ�^w�򹃽��1�������=$&�=���=8��="=�;P=_��=�4��	�?!�?���>��>_���Q+F��M� �T>��q>z_�=��>	�>���>��>��F>d=�槾�������)�>L��>��X��=���P>�6W>�la>>\s?��?ʆ3�ɾec9���L>J�>��!?8R?���>Kv�=(�������lӿQ$��!�}�N��ۈ;s�<���M�X�7$�-�������<��\>�>�p>E>=�>�;3>S�>�HG>�ׄ=�=C��;�;��E��M=�o6G<n�P�ڔ���Ƽ����6����I���>��+��*ټw��>�)?3|�=�墼%M�Lc��$�c�~>�@�>1ה>n��>ZuE>��jQ��&H�	b���?^{T?d�=��t����=�
��^�>�Fo>��>�~�>1�'��pq�H�پ�Z�>L��>��3?�i>(�=���g���Y�$��ܲ�>��<\���
��?j�~?<�$���K�g�Z�.��?�n>ϫY�w��+���+���:��N.�z}��z���O>N��>�}?wl�І����a�m�?����%=���>Ll�=��3?b�>�GO����],�ך������0�<S�U>-0�=;-?�h�>� ?��^?�i?�i?������)?�о>[?�
.?�?S?��>���<\�>&��>6�>*�>��㽚J��KMv=�»<v
�<�<>'��=s떼JG۽4��=g
�=�&���<]毻i��<=p�<������<��=�&?��
?�^�\Z�����w03���<��)>�X>?M>�ж�v�>��90n�>�}�>#��>=m=n�Ӿ�[�%������>��>�?Ϡ?wI�h~&<o���+u� H>��>�s=g�lX��H��W�.6�>�Qb>M�l>;6>�p?��E?5�=?v~�K�,�/f��5�4J���
<t7�>}r�>��^=/8��b�1��x�f�%������VoE�T�\��>%��>5��>�*�=��r>)�_�R�����M���T�l=��>���>�	?��>�����־�Ծ��t�J?qN#�n2���2�վΡ����G>^��>nx��;�?�쇾f?��P���Z+�HBB?���?ZK�?�|C?P��F%>�{=��H�_��.�B>@~�>��.<����8՚>�È=M���ދ%��Y�>/�?0h�>Ţ�<yD"���A����޿�Z��`�<Z���G�Ѿ@. �Ft��%9����.��=�꾾'N��$���u�4f/�4�Ҿ��ξ�����Ͼ�9}?�c?��>������Y-P����ɂ>����%=:U�������{侾��(�پ'�����������۰�>��꥝�𱏿7#���i>H]|>|$?Ξ��ب���0����kkr>3d�>y��V�`�gŗ�����TQ`?�?T��?\¾��8�=_����?�>BV>Vp���'��3ğ=��*?��e?O�>�ʌ�^옿c�����?���?SAI?����[e��RC����<?U%B? ��>�w������׾~Ջ>ǖb?u�S?��$�?l\�O}#���>e�v?$���3�>���>�u�>D�O����q��=�Ծ}OV�e�>�\�a�L=?=��y5Ծ̩ϽHn�>�Й>>ʑ������O�>uq���8���P��$��Ԡ���>�?J���ӻ<�]}>q���WF<�*����U�b�l�RB?�?�j%?��]?����'D��p����>"M?\��>��>�#��c�>;?����Y�'C徑�G?m��?zh�?X�E?�;d��)��`~�����c
��d���2�=���>3�/��	> v
>wM4>
�->[�(>b!.>
�=l~">\��=���=wo>�W��J� ����Xm��.�����H'��"VǾ����?�	�i* �w'|����)S`�����/Xؽ^񵾻
�d��==[˾	�>~��>i�>�Z�>�=R��>^�ݾ�K���컽�xO�����U�⾪���}��u���T拾1[���k=WA��Fn�>�}�<`NK>QO?>��Y���V>��?>�x�=�]D>K�2>���=Q>��.>��3>�2L>J�z>��=�Χ>�Ԗ�l��A߇��G�#���YI<6�I?�ɽ����?��{@������s��>��(?�b�>��#��A��gqd���>w�Z���$��̽c���^�>_��>x<�=���<7?�� �����|k>��>��
>)�s�Ͼ�Bнݤ6>��>�����>lJ�>%'(?��x?[?.#=�>�>Mjh>+a�=��>�S>$6�>��?��6?Y.?{D?�� >��=����=�z"=|Q�Ar�p�/��*=����l;�Z���]��	�3=���H��=p��=Ѣ�=I�=�$�<�_?�J)?^��>��>�aսc�Y�5`���v>R>]���+�>>�?��?�q�>���>�a�������% /����>���>�P�g����5��rX�>��Ľ��t?[z?�$=������lQ�H=�=>�?�^?�>\��>�����}�$2ǿH+���;SZ��˩Ž"�{��[��z#�_F-��v ��^��&>ĳ�=7�6=&��=��.=�(>�B>�I�>-P>�.�=y��<gA:=����F�K��=%����b�_�(�{ǚ��/a�����7ؼ[�f<��
<�ns���%����>u�/?��0>�F��g�ƽ�ž
��
�>��>���>[˩>��>:���sO��3��UU<m�6?��X?!��>����7�=ax�����>�>��=�r�>�nB������Ӿ't>YD�>�c*?\�B>��<�|��Ϟ���w9��t�>��<�u���?�Wb??��Ծ������D>�߽�I>���Ҭ���V�K���2�fz�m��������=uM?"�?;���\d�=��ܾ�꠿�h��=�/��3�=\�>dm?�j�>2�������5���վ�*L�s'=�6V>·��K�>w�?�o%?ڙb?-�?H+?ro8�"S�>hC>���>6�>��>̆�>7��>�"T>��>���8=tt��a��`��=�M�<�?�=��+>^��=����=���;&�<��<�6���=1�9=/t}=���=\��=S�=�,?�?}z�U
V�/�=����	���T�==��>��>�ᐾ$�G>�#�>?/�>��?�>L=>�w�1fξ}3�@�>G�>D�7?dq?=_=�п����_h��W~�>�Oz>5N�����3�+�����B�齽+�>��>r�y>e��=>�~?�S?��5?	C����&�J*<� �/�3md���s���c>kJ�>�}�=��x� ��nv�5N��l4���ν��M�9��:�=E�=�-s>$R�º�>)��rd �-߽(�}��[���#�>���>Z�?;
Q����ϾY�!�^�>?�����;�����`߼/>�_��7��>W��w$w>5Qp�Z䁿K۩�p���y�>��?,��?d�u?ڧ���;=D�����>8����X>��M>	-�����А�>X�>gx8�և,���꽽q�>+��=A)�=�"����R6-�g�ǿһQ�u>��eݯ��UH��޾f�]M�����ޟ��"F��dE<�&��Y��^T�s�|��%��򨾐�M��P^?�� ?v�T>ظ���B�������y����=�)����{�b+þ�Qվ������(�A�Ϫ��Ѿam�ٰ�/��>�WоM���9���X��/ZL>:�U>�7?A�0��a��q��~V�\IQ>u��>�&��"m�������&��Y?c�#?���jw���P��Kl�;�>���>IC�=������s���>t�(?\&Y?x)0>����$
������?N��?�b?z徉�Y��5��>��J,?��9?Xӫ>�pJ���;��μs>,ot?�Q^?eM���e�y����?��r?n n�7�>��>��>.g��F�侌��=}��_I���q>
�Q��2p������p��L}>�8�>��a�qa���>!';�z+m�U�d�7�6���ٻ���>���>b���>���>�)��d�� ���4����|>���?햹?B*?�d?4�6�i�C��C��8���1?��,?��>M�71�>Al?qX�L���ﾨ�=��?<��?2A�?��q��տv󑿌}��x<��Ah�=#ژ���E=��"�(EH=2a���!�<P�=��o>E��>
�>���>#�">��>�>�����#�O��b;���<�o�;��(��+���z��n��[���;OpJ�����yS��{���A�w��c��?�S�N�ܾ� ����/?�m���6?���}/>μ�������4l����=>����fH�"���þ�EL������2�=&о�h�>��A>�0P>�]�>��P���:>w�=i�>���>���>�0#�;��>v�=֎	>~��=\x)>��K>a�>0�=�����h��,�:�j�U��[�U�D?rzO����y�/���о	U��y��>?3
?�Q?>{�*�1F��
�r��T�>T����*p�	ո�d� �)�>w��>*��=�$+�Y���^�m���н��>-Ƈ>��>�@ݼ1#��4���5�=���>�8�����=�܌>|&?xo?:�7?Ό>�>��G>��k>�)>yck>�NO>�$�>��?Mh.?�d.?)N?��= u���7=
��=M���8��<1������vׯ��:�૽�l�=�O�=�(�<��=�3�=��_�H�"���'<P??U�H?r��>��>������E�!�Xy>;a�>�]o���?���>��>:�;?�la>�˽�6��Zx���پ���>�lf>P�U��sg��@���0 =ò>�[m?�|3?��k��㣽)�>\C�=�p�>v��>�?���>�Ǭ>v�>g���gӿ�	$���!�#ł������;��<��ZM��:9�j-�������<�D\>��>K{p>�D>�n>�q3> r�>� G>-�=���=��;PT;V&F� N=�`�T�H<�P�L����żs˗�1�����H�=�=�PI���׼�[?��?�{(�H�����f�9��T����>��?̡g>�&�>�Uf=5���.��Y;����6� ?D)_?$��>7�/�y:$=��<�ā��@�>�l�>j`�sd�����5P���>��?Q�?Ef�=3���EC�����-%��f>�=����?��4?�ô�����݁>�ߠJ��K'�|�廍gB��P�,Z��`|��6��o㾞��@�o��J���>=>�?濰�|vX>�ؾ�茿�;���m�������f��C��>�[�=d�k=��T��������D!��N�cCa>Ӗ�>���>�	�>	�D?��T?W�(?o��>`�
>�%?=�/�65�;��>?��)?��? 	7?н�w3>��=u�>s�)�T�s�_�=U4=A��=�C>��;>���1��=�N`=�����^Ґ<���<�{���g)=ZZ�=`q�=vG7�m?�^#?�8��=�-˽��<?�ܽJ��>�>���j/���u�>��>�V'?O�?��m<FW��Ϭ�PYʽ��۾X�Q��?t�/?�?_��=�U=�2 ����RԤ>P֪=�q>�\�K��ޖ�����֓>��<>@/���@j>�m�?��7?�?S���ô;��/��5�5��Z!�{���>�L�>�����{>�R	��?Z�3�_���>��$�қ=��E`>�y���=�W���M%��U>�g�>V�B>���hl�=��>�Wh>�r?i��>Xj�9�\ս(���qa$��.?�t>��B��)QY��<@����>f��>cd��l9�@kY?�Ӌ��.����I���j��R�>��?	��?��b?����K�9��W?7��>�/����1>i#��l�����o1�>q	��5�������g�y��e�=���>�<�fԾ�s¾�����C�I�O�p��<�����F����3������վ���:��< ��ա��K�q>�柾���f6K��� ��|Q�ƾ�c?9G+?�rC>�g�����վ��赨=E.��?��<�Wh�c����@��8�%���߾�g
��K�}I�"�}�;��>���ս��#�s�*�-�
����>�3?�����ӾI�	�h$>��>���=�۽�̲��f����H�x�U?j7?�=�Ғ��1��F>h�?s2�>t��=%�����<�{�>:�/?�+M?�5
<�a���Ƈ����=찱?C��?�f=?���c�/�����ht&���?���>Ĕ�>�$�F�;gꐽ�?f/7?���>��@���u����>3mW?/�U��;2>��>���>��ק~����������L�w>b@��#�#�
NQ��
q�'�=��>�q>ΓN��.���>�J�Q딿��\��W���=a�/?�?��3�a�?�5�>�E;:������V�l����Psw?$��?`?��O?��b�沣��:�>�Z.��
?fӢ>�!u>b:�q4?��8?z�BԾ#־��=��?2j�?��f?�CS���ڿuj��.J���(���>���=)�=����� �=,�=��U��������<�JR>��>�}0>W>EqS>Mg>*=��X�$�Y��a���c�2�������ь,������Q�d��
Nоٲ۾��D���S��4��r�<�lf޻��佮[0<e�!?�ސ���N?�)��s>����2����Ծ�
#���
����N�����Q��H�V�Y�r<�RyžA ?�M�<�g>�1�>h�ʽ׻f=���=��d>%�6>���>>�%>�K>pk���{��ک�]a�=� =�[3>���=�k�������,�I�n��L=��'?._�J���C�@�����A�о9.&>B��>�d>g%�Lf��UW]���>I{�i���1]%�\�V"%>�v?mp><=>��S���2��X�=��;>٪>>ә�=��=��:����V>� �>ϴ־<j�=Fpv>)�(?�v?ks6?�u�=��>�a>�|�>��=L>��P>�׈>��?!�9?�1?W*�>U�=[�`�'�=NE<=��=� |S��?���3�<&$�1ʉ<��1��#I=!�q=�&<�[=9?=��ļB�;���<���>��J?�>��?���,jN�:�/��o�>���>"���&�>���>]_/?��I?�f�>>"�⼭`��6�澳�>7�t>�g��OH�������=>$\�?�$?��������4x>��G��Ũ>�T�>˂?G�?�+�>��{>����ܼ����V�0���=�<<��E�%����q�1��r��u%�t$|��g�=U�->x��2d��ƛ�={!�>���>T�>q8>
�=���xe5뽹����)�m�</�T=X��={�='������?n�\�F�*�����=c�?ܴ?lN\�w���]q������������>Ϛ�>��>j ?��&>r���(D��8C��o�$��>
�S?)?
?�@3����=����{�����>�>�>���=2M*�	[Ͻ������=?^�>J9?Ś>o�3�TV��?t�����>�G�=�aR����?ְZ?$��'ま+��(M�����>���Tɽ�[��;�+���J����������}�h�=���>Q��?�Ӿ�� ?�[�O"����d�����vo�>�>�I.?F>~|�BLa�dm�В��/����vs��)?�ӡ<��?��T?�.?�0o?	?��_>%W�>��/?l˾F4�=��<???O�E?�5?o��N� >�ݘ=N\�<��/�2>��i��=l½B'>��>�N#>.����=�f���Qӽ��<�Cl=�v`��=�������<=��>�?�'?��$�j�s��>=ؾ�l"��9�>V��>�w��������=_P�=��>E�<?2B?V�>����[پ�/�G�4��?ę	?]�?;=W�!>���<�(���=Y�_>C�ݽ�[���	��	�Ծ�o�7�>�\><�޽��b>�b?k��>AZ6?u,U�>�ؾK&V�����s�>��=f?�\�>nRa>t�1>S�4���g�I�q��s�=�>��н�a<�D>v�E=��>�.=���=Q��=��4���}��><������>컘>:��>��2>��=�K�|����h?�(0��H�G�_�n���?[?�
-�R�8���D?�5���$����l��i�A?��?{	�?�
T?!��=5�T�0?��z>�^Ӽ�B�=�ξ�֑�I���x�=��������pG���t)��e>x��>k큽�%#����y<��Ŀ�&�F
=��!���{ 	�)��Zԯ�<��j@��3��:0?�QX��\�T��^�0繾4s۾��e֔���?� v?����~�̏� W��/�����<��J���Խ1ؾ�%��䥷��žݙ���c��gU�T�������>?xC�r#������/�"��|8���T>$�!?��ľ�츾u["�N,�;�·={����"_�������<=P?�~B?-���.�p���B�=�,�>�x�>0[v>�	���M��e
~>C}&?��&?)��U��r~��Y=��?���?��??~)P���A�}������	?D�?bg�>[��V�˾�}��_?b:? ��>�!�����o�y��>a[??0M�-`>���><1�>�`轧�����,��w��ܡ��w8>{� �> �)%g�(�=�J�=��>�y>�]����H��>��	1���X�p����G��H�=k�?(+���^>��B>`��=�Y��S������t���51?C�?�Q?�eC?�������(�p��'��> ��>�#>]Qp�OU�>�}�>�����P`�1پ��'?�?���?(>?)�b��7Կ���������Ͼ4k�=��=|��=Rq=�#s>$�X<���r<�;>�Cl>΂=)l�=	�;>�G!>��>?K��(����+��L�H�%�*�ae����{��"f��	�=��p񡾨#3��Ct�d[�*|��B�i�4=罺VžsE�:�$?@ú�!�?�8�x�	>����.����μ����3g���?��%��7��nҾ�l¾�Q1=ʉ<x�C���s?Y����R>H�j>*�ɽ7��>���=�>~(C>��>X!>B�J>WW<�@�>��<9�=.���_x>�����≿�={���v��O�<���>]F4?-0����=H�S�<$B���Q���>��N?7T�>)�L�z����G��� ?\t���w��"��<��=��?N�>�|뻷�k��K�= g��1^b�=z�>Ł>.��=�����i�	v罗��> �w��^�=p��=D.?�ik?V�?i��>��>�˽7~�>�@>���<F�~>-K�>�0'?ӲT?�xA?��>ss=� D�#�=R4>���uͺ=@�S�?��n'���>灠=��=���=�x߽%����޻�PI=��Y=f4����>�tQ?9��>.>9?#ʈ���6���\��Ծ}t�>�Z�7*r>�?�}�>�R?m(�>sm?0~�>!��,� ���>7�Y=K�W��SE��,��:�>K��>�U?
�?�a����S�����?��>q��>��?i?��=+�J�n��e>ӿϥ#�Ap!�v���(��{D�;j~=���H�d�9-�.�O���q��<�B[>�e�>��o>�C>��>=�2>�s�>�aF>�`�=o=�=��;ܶ;M�A�O�J=Q���]< N�3ʹ�j�¼"f���#���G��m@����=�Ѽ^?�-?)R���bռ�$���p������5�>R_�>剬>��?H�+>�z��2D��*�ۜJ�:"?��w?���>�Yo��β=N^�=2ʞ<Ҧ�>��>�V�=u���k��H�Ox�=�(	?��?�Ջ>W�_�:�d����� �%w>h=��{�:ݏ?�|O?h߾phb�|�,���7�Y�	�]R7>򝰼><��g;��@e&���4�1�����v-�3#=m��>�S�?�*��Cx>��Œ����^�M��m�=�_�=�H�>���>3<��K�O��RVؾ�C����WY�>*��=�D�>�@?>��>�Qm?�?��w>���7?��7Ϻ>l��>�G�>&5�>z�?��>u�>�lH=f�n��X����q�<|,f=$�$=�DM=��>_���
�=�
�=٨��b���H�<���=:��=�Z��&=�f�==7p>��
?�=?��\��1�=E� >k���x��W>V��>=.Ӿ;�)��[�=jx��%?DC'?���>��>�����:�4�¾S�D<��>�'?�x�>2?�E�L>k&����þ�5�=>�<>[:�<0��b����/�SH��=%��>�-?>Ͱ^>�st?w�>?�A?䧋�N�4�?�d��@�%�T���d=Y��>y��>%><���=���V��t=��r��2'�����>�K>>��m>���=��9��/-=���Z1>
=,�U�ؽ�r�=a��>�{?���>e̯>{>j����HK?di��Q��Tʙ�T�վ(�׼�">W>����>c��&W|�x>��#A2����>Dm�?�}�?�@b?�1<�/��h_>osG>p>���<�'�i�c���P�D�/>
�=�1�����e��
�Y>��o>2ѽR*þ�c྇�a�<Կ�<'�n�=[๾@���? )�������μ���={�L�.�M���o��=}7��Ⱦ�:Ծw�Ǿþl���Y�j?T�.?� ��β��v#����X�I� l�<��Ѿ���gH��'����-��\��غC��4���U ���=l�����>]D��-����J�:�/��#�>{��>c?S),�]=@��qP�Th��32=5�>A��cm��᜿��8��97?��?��:��7ҾKL��O!m>M?{�>�*�=�ѽ�w���.T��!?�hO?<^8�k���݉��췉=�|�?�f�?sL7?�ų�4�`�;�y���8�?��$?5��=
y�ޑ/<K/��Jy>��]?-Ǔ�s.�����+'���?H��?ɛ��˂?��)?��J>s�N���	�l�*о��z>)^�>U˽$!>fjƾ	 �&ٶ=6��t��>k��"��X�>�r�=f�:�B�GN�
7�< �W>���>U����b>\K�>�s=���� ���Wk�J�D?/��?�Vm?�K0?q0�����ټ(�1>]м>^��>"|<���%i>H*�>]&���c�|꾠�?��?0��?Iځ?��~��gۿ�����˾H����>�o�=N�>W����<�=�߫=�밻*N����=��>�zz>G�\>�>O.V>�]s>e��O�-�J^��v3���r;�8�?���%=��������r�����{�����j��34���)���1�v���U��dX;vTt>\۪>��>8Ӽ�:�=54� W��^s��ƥ���Ҿ^O{�$l��t���b쥾��A�N̗�z�u�gľ?�!?O%>���=I�|>��)>q�<�8	>I[�.B�=u�N>8>�&�����=���>z?�=%">!�>4�<>t��=Α��w������R�7ؽ�c(?�Bc��ξ�,�-�ž�:����>�?�X>m= �gi��T\���>��sΌ��F���Gƽm�>�}�>r�P>J��:x�,�� C���t�l-�=j:�>/��=w�W�ޞ��(��^�N>�9�>����~�>�y=�*B?�l{?	�?bm�=U��>�	�=�'=��*>I��=�a�>���>��>r]&?k?	�{>��b=�����=��=I��}U<��5��M�=��	� K����)���D��s�=�R�S,�=2�h<}�=�=P�ӽ��>R1S?։�>�]�>}�4�%j��(����=��>�0���(? Y�>�>L=p!&?���>`��>�8�>���Ҷ^��~�>�>$�e�l���#��_[=d^ؽ�'p?-dZ?G"�=0���x��<�	��f,�=5�`?�^?'Z�>�I�>P�=�� �i�Ϳ�fM�Y���~�=��>��v��y��a<	;���?ž�V��"�O>|Ո>���>7��=��$��#�<���=Q�>��0>��5>�m�=�0;��5��Vq��]B���=4>az�S�D=<5=֊뻹����M��$߳�������TD?2^?On_���H��Ѿ�_��K5��޿>�
�>��?r��>��V=�������51�A��n|?�cj?� ?�����L=@z�=J��ZL?�Z�>.�1>9�l��:;�����h@�����>�>�L8?1�l�O�O�Ut��,1>h�<C��߂?�h�?�B��������.�~���dS�=k2�u&�>F�;�mj��=����S9�����Q=�=�r�><{g?�����fK=�+�z��!�Q�w����=��>l��>�e+�V������CU����xC�;���|��>T��=(�M>��&?\�>#�X?�?%?��r>�/�<1�?�e�x>xO�>z��=�??X$?i�>]�>0�4��������]�=��=g෼H�>("E>Xz=s����>����r^�J��<R>�Qֽ�O�>��>�a+>^���g�>��3?�"">4ހ=�a�>�0<��X��j?��'?�ݾݘ���S>,���>L�K?u]?C�>���h��l���ب�3��>06?�d�>r�=*��=Op.��ׯ�����w��=�W�<��a=�������F�x�
�=�10��3�=}^><,�?�1?'E?}RX�`�4��xg�D���3���	���2?�L4?�:��� �+*b�$|���d4���B�rFѽ��=�z�4�:�q>{�p={��=Wݵ=��g=}Խ�A�=��&>*S>a�>q`?r;�>�2ڼ�Ԋ���~�[l9?�wN��#ƾ[�۾�ɽ��$�C�(�^v�>�l>A��>���}l�/���c����?!6�?���?/?�f���a̽��+>b0>v�S=H�=S40��ޓ�ڗ�=�>�v=ӷ쾆��Q�H��=�M>���4۾���x�=����(�J\���d���|/��M�R��(���M]�E��<�־qm���^Ͻ!O�ٷ���X��o8�����+����?� �?G�C���<)}Ӿ��S���.��k�޾@yR�2DX�Q�����������~.��<����"J��S�ھ��>���o����{�����Ք�Z/�>Z�	?������>�׾����.?��J��1�=*����{����B��?w?�#"����������d=�݌?5z<?~]�>=����TX�>�O?�A<?� B>�	���,�����=�9�?ʐ�?4w?�׾UBa�4��/y�֩7?��?�j�>��Q��7�>�ԋ>j>�q?�:�'�i�P�v�"���%�?��p?�ǌ��.�>�3?���>�o��{<,�V��"��Z��=e��=�䅽�%�=�٤�Gl�	�>'B�>��u=����䴾ˁ1?cQ����H���`5�'�%>״�>��>��\��k"?G�?���=�&C��닿�$���D}�?���?f�?�:
?)qܾ�����=t)>��(>)$����=��6>�Ԏ>�z?���@�V�s&��8�?_Y�?"��?�F?r-����Կ{����ƶ��r��X�>5!>o�>�t�����=�M�=�\��)�:���=�p�>�\C>U�>ǪX>��->�#b>J���a(�3/�����?B�����j��a}�`���@��Dڣ�����C����G����<��V����p�=7v�A[>՛?�>�O�>(]>��>�	��O�Ҿ�6{��I�C���Jپsi �:j����;�t�o4\�![���ⱽ~��6?�ֽ{>D��>��F<��<�V>z��=8ZI>�>��x>%m�>��.>C�@>o>�=���=�r=a�<��>脿͋��-�)���&�0@�=� �>;�=]s)��X��2h��x#=� �1�v�	?���>�*�i���������>�H��h#��	�=0��=
��t@?1�A���ֽ�V!9k� �����j��z���`��l������L�?�=n��>�k�����=��u>|;?�J|?[�?��=�>\�=v<>~�>I�>���>
W�>��?^g2?�C?��?��=�A��>��9��6��ڤ<�YֽC���.i���w�<�>����j=��=X��j=�z¼�o��ܢ�<d�I���>�?�S!?��>-4�f�?���ŻA�*�=����&?�h�>�6@?�3??;D�>z�>}諭֘���5�lݶ>=��>�k~��nI������{~>����\|�?@?0���hp�=F�࿎����>��>��(?gC>��>1�	���˿5�	���&���8�|�>� �=V=2=x&�=�����Dz�ʟ�>�Ӽ>���>݃�>\(&=V�	>R��>N��>b�=���=j�K>�B�;���;��=�E =�u�9l=�=8�l�ʼ̘�=􀍽����'
=P�ν4�
������	?��>;���e�R��`P߾'둾�[R>���>��>�ܐ>cx��D�éd�+�C���"����>��?%˃>�섾��� ��=�y����7?`o�>�>�B�y�m�~5ľ1����?P�C?9?w*�� �|��V��l���=糤=�����?��+?@�x�G|��H�0�>�g��~�D0��_��.<Q3���	�t�<��T��}��F��F���>!n�?g�����=��
�VX��~�|��'��Ͱ�<tQG>qc?X�\>a[g�O�X�����T���g`��}뽂�|>��=�S?��"?�� ?NO�?�GC?���>%>-#?Pܙ�H�\;̠�>�H1��e?7�M?�KQ> J>�G�<�>Ɏ��h��:AO�֮����>,��>�)߻�`�E	�< �{&�_	=�Rn=��Q>�Q
>2)>�L>|G�=�>���>i[S?G���8�v�P=$.��Ц��K?(��>豳�r��=d>-h�{�!?�b;?�w
?��v��J��Y�X���̾���=���>-p(?�?�>M?��I@�=H`����a�~�[>sJ�<��<+r�D'�<¯��r��@�>r��=�3>�=G>�,]?� =?`�z?�G�<:6��a��7)�]>NP�H�>T%�>���>u}c��.�����$Z����;�������) ��C>)�>�=�M�=���>���=ȟ����=�p۽l�>��N>�L ?芕�a.
�9�]���1p?m���A�˶����?���l>�a�>���=�.�R�-?�Z>�:�D∿Y���"?�&�?SA�?q��?�Ԣ���U4#?ȳ>��=�����Ѭ���F�5�v�>&�ֽ�����Ͼ�G�0	�9{��>��?=	��٦��`9=#����3�tE�xa��ࠏ�����⍞��3��[4�C�J�X�$���~�sg���:�yF�=w����z�X���A8��R��?)��?�9S�Be־�L�U�-��X��D�=��Խub����MT侫��Ӓ � �Y�M����	�sO6�r����>����h�C����S�u�t��G6?���>��3�K�!>�D�in��
>}"�b�@�g�}�]&o��	g�g;�?�{�?�R��N��hŽ~�O���z?;��>�+�>Y�E��%>�?��Z?�{?��"=�3��&J���ہ>���?�b�?P�<?�FR���:�e���Fƽ�?�7?���>>M��%"˾aK
�?Ȇ;?Z�>9�%큿�W���>?J?��I��5`>&
�>04�>�߽t����������m��D�'>]��<�餽�o7�z�/x�=1��>��e>��i�����r�>����s�	�k��"�N��=̱�=xL?Qࣾ�w�>crV>���>����܌�ĭ�����5B?��?9O^?-�y?=|g��(�tG�nΚ>�?���>
'�>��<5��>�F?�V�`��@�{��>�n�?BJ�?%7?L��l�ؿ:^���\��*��i�ٻW��<���>Q>z=��]=7ȡ<i�[����:4;>>bm>��s>0�>��D>�]L>���=
t��/�W����{���I>�������p��9۾�I{�Y`>���������@�Խ�X��q���pd�E�0�l�O�
���-=�(�>.�I>|}?LǕ=�f�="���%��Ŀ����H�>��H-�����2���P���Ƚ��F���=y���Ҿ�)�>����� o=�>�m0>
A>P5�>uq!>�j =`�=S��=�'u>@P@=��<%��=�	>�rջɑ�>u��\q�V�i��m�8��*<��]?KU��0����B��Z�3�ݾ:�|>#4?`��>��1����c�K�_��>��}=�Oҽ�+*��×��ڨ>H�>���=��=��~��R������
>v�>���=�E��i}��K��Ć�=��>�Oݾ���=��V>�)"?$�?R�5?©>���>��?>+��>�,�<�3>�R_>Q�>��?R�$?(?� �>��=��O�n��<~��=_�M���b���ĽK�B��A���
MA�Y�<�ő=u�<<�E��';}�\�P3�<j�<���>�[?m��>�J#>g����*!�*��'C����=f�����>Ϊ?�?
	�>�ʲ>���=' ������<�S5�>���=x�O�t����z;�M�>��>��P?�^?���=q�����>4ؼ�?�`�>,�O?[��>~��>��=��AͿ��2��y)�!�n�z��E =�� �����W�xս�t�<��S>���>��c>��%>:�>�F >A_�>t�R>Ws�="k�=�-�<�ᢻ=���a���'��==%�~��2м�1E��c�ǿx��ؽ�_ֽz��������?��!?��H=k�&<�5	��e��վ�)ٽ��`>aW>��1>66D�5^&�<'�sR��˳���?���?�U$?�`����=��S���:��=*�Z>fĀ=Z���dS>�D���=>O4?`,?��|>��B��f���s�;��"��>�=���6�?*�O?>Ծ⁾F��)�:�,�j�*�2�F���Ҿw�Ѿ�`-���>��C��}��;cC���>][�>��?�����S>3�U�pI���ƅ�u%��7j�|+�S{�>:�>����	�>%��Y�J�<&�r>���>p�-����>�Vg?\؈?��P?��=?l��?���J@?��\>=�y?��/?.�f?�u?�?H�>��>{�>��^ �
�{��,���G�����=��|>1j��d�<�Y�<G�;��>�w�K�f�
���!��=�f�����<y:'>�>�r?�?o�
=�I�<�9>��}1�9��=��4>�%?рB>[��0��<�&%>X($?�"?��>��^>�飾�@��>��֝�< �?IX?�?��Ž�gJ>^=վ����U	>�8�>��B��N6�����h.R���z>,�f>�>Z�A=V|?�W!?���>�!���}��`�b�L�Y�ٓ��J�u�h�> �=���>M��?41�].��;�l�h�D�=�;����I>]|%>���<���u�J=}�t>5�>r�q�������=���ץ?�8Z>�/?��>������]�G���g?�]T�j�v�m��.(>�½=B0����>�غ�fv�>���L*3�����ݝ�<�?r��?α�?yj?+r��P	��3�>5$d>2 >��<9���B-:�8���=@򝾓*�ݧ������>F�?�0�=2���H�@��=�=ٿ��!���<��~ؾ����K�	��]��$Z��w�׾R�ҽ��<m7���W�0�ٽ@ý�ԥ�.T ���澕S���<�?�c�?g��>�F<����`"�p���|G�,��i�J�8�-�l���Ǿ�������N1��~"�n' �}(����=�a)�U?~���{�:�*�-&����=��>�Q����������</=�=E�>-�<����R��X���b�a?�WV?�k�U�{Ȓ��=jJ
?�:�>M?�>�f����5=�>��,?C�?a�8�����0.s�ӊ=�`�?��?'�??�R�͎@�t��2����?��?��>�l����;Q(��~�?@�8?�	�>=��ޙ��uO����>�]Z?�AN��Sd>.!�>,�>p2�����b-�h������M7>����k���g�S�?����=�%�>Qcy>�Y��ŭ�L�?fiҾM9��3PE�$@#�ϼ�"�x���E?�'�Ib(��W�>m��>*b-�Ӄ�����$=��b0?�ɳ?=�?�?�+u��;i�V;}S����!�&��>2<��(�|Ҏ>�B?k��֌��h&��I�>?��?�K@�͇?������ٿ�)���^پ��о�Ԭ=m��/�E>kr���	>��=ٵ_=1X���f=Z,�>#�a>�)>o��>�D2>De
>�e��C�!�"���ޔ�;B@�]�+����E!ڽ��n�>�y7�Ƶ�J���]/�=�X�࿕��o����R���/<N�2�ˢ+>,��>�D�=���>d��>:��>R���Td������&'���(��j�z�Ծ�������n���h��?��m�$��'?���=��%��h'?�z���=���>��>�_"=}��>��F>��>kt�>�=�>�a6=��.>�>P=���>ާ>�ᒿ
�M����6����j?Q����W��cM^�Aʊ���ھV!>N�>���>��S�ѥ��p��?�"�X�Ͼa����=r��>ʉ�>�m>A����=U���zž����d>2�>�!�<7ž�H/���&>�l�>��`�Ȣ�>�7�>69?���?��Q?2�=��>�M>���>��=I�>ݴ�>		?�
/?�^?B�U?/�>���<�5_�X=v��0\*�������3�兽ִ���R��� >A��=�m={� �Z�r>Ǎ>(K���=�=9x�<y��>�{f?���>�r1=rWӾW�0��Z�'T����=�=#@>$�?]��>-]�>��e>�sb>ae��m���a>�0?;[=�ד�X�����=�q/>��*>4}�?�c>?��>S3��]4�=Y3��ۨ> ?鯀?7��>�T>�N�=�����˿*�%��oP��־ф��0=qF�;x�3�'���s*=;\�
=0*>\�>��>"7>�,e>-B=O��=�;�>v�Q>���=Z>.�s<E@�=�|��;�g<���� �Ũ���; �<k�<�ν��X� �;���
Ks��?y!?��<�A�L��׽����4�U��>9\�>���>W�>�Z����@�H�X��%<�-�Z;8;?ȯY?k��>��Ͼ%U�;��K=S>>9?�^�>5��>�\��dま1�)�~�W��>C�C?g�>e!��S�{��pq��=��Li>���=��g��Ӏ?���?�������$������y ���7	��Sf߾�W征�� �k������S+���,��>�O?R8�?:��l&�>�r�E����$�����c8}>���=�Ð=��>�A�*�Q,�&,̾ݐG�QDʾS2�>��(>}�<�7?j�-?��?�HL?�S:?�s>݄O>��>z[K?�E>�0L?:�"?�":?+�A>�@>���>�!n<=	���h�����<�Ȧ�<��=���=mx�='�<��c�E�O�Y׽�s���z<��E�N�D���
=��Ǽ�t�=��?h�8?�d�}{}=E���B�p�8�=�N�>j*�=`kK�c�&>�d>���>3�?��>��>����{� � �4�2;}�?4�R??g?�|�=Z
�>a���$���5��L?>��;���X�|���W��'�o��>��o>�7�=��>���?�@�>إ?��<{�� �������C?�����þ��>|���R�3�\�e��K�&���g�� ��-C�F��>N�'>?�?���s=0�F>��t>^d>:QZ���=�0g>����ٸ�>$ �>5*�>oG�=5�>������h�9�]?�;ż����  ����UF����ޙG>�|�=\fN?�X�X�n��H���P<�a�>@��?�J�?�[?�VH�~~2�1O>>�2�>���>Z�>dD���k=��*�2T6>��<��4�����������=��=YB]�V)��sڲ��P�=Fڴ�YJB�^	��Þ��/)���۾5���n��a�P�V!\��F;L��Y�l��.�����Ty��놾f����y����?<,�?�Ό>bo> �A. �*�*���[��>��F�H�↾K96��ԏ�	���.���6����,���\��d����>��<�!���6)��n��� H,=����L?���S�D��3<��*��0�H=�L�����p�J"��L�žKua?0�??Y���������3?���?���>���=d�E��2w���?Q�=?�J?d�Z�2������O��=d,�?���?��??�O�D�A�o�����-?�?c��>u����;���K?'�9?S��>���g��f=� �>��[?�>N��b>��>0S�>S��Ώ��9�%�!/��rH����9>[�� ���*h�)	>�" �=��>gfx>3]�� ��L�?fiҾM9��3PE�$@#�ϼ�"�x���E?�'�Ib(��W�>m��>*b-�Ӄ�����$=��b0?�ɳ?=�?�?�+u��;i�V;}S����!�&��>2<��(�|Ҏ>�B?k��֌��h&��I�>?��?�K@�͇?������ٿ�)���^پ��о�Ԭ=m��/�E>kr���	>��=ٵ_=1X���f=Z,�>#�a>�)>o��>�D2>De
>�e��C�!�"���ޔ�;B@�]�+����E!ڽ��n�>�y7�Ƶ�J���]/�=�X�࿕��o����R���/<N�2�ˢ+>,��>�D�=���>d��>:��>R���Td������&'���(��j�z�Ծ�������n���h��?��m�$��'?���=��%��h'?�z���=���>��>�_"=}��>��F>��>kt�>�=�>�a6=��.>�>P=���>ާ>�ᒿ
�M����6����j?Q����W��cM^�Aʊ���ھV!>N�>���>��S�ѥ��p��?�"�X�Ͼa����=r��>ʉ�>�m>A����=U���zž����d>2�>�!�<7ž�H/���&>�l�>��`�Ȣ�>�7�>69?���?��Q?2�=��>�M>���>��=I�>ݴ�>		?�
/?�^?B�U?/�>���<�5_�X=v��0\*�������3�兽ִ���R��� >A��=�m={� �Z�r>Ǎ>(K���=�=9x�<y��>�{f?���>�r1=rWӾW�0��Z�'T����=�=#@>$�?]��>-]�>��e>�sb>ae��m���a>�0?;[=�ד�X�����=�q/>��*>4}�?�c>?��>S3��]4�=Y3��ۨ> ?鯀?7��>�T>�N�=�����˿*�%��oP��־ф��0=qF�;x�3�'���s*=;\�
=0*>\�>��>"7>�,e>-B=O��=�;�>v�Q>���=Z>.�s<E@�=�|��;�g<���� �Ũ���; �<k�<�ν��X� �;���
Ks��?y!?��<�A�L��׽����4�U��>9\�>���>W�>�Z����@�H�X��%<�-�Z;8;?ȯY?k��>��Ͼ%U�;��K=S>>9?�^�>5��>�\��dま1�)�~�W��>C�C?g�>e!��S�{��pq��=��Li>���=��g��Ӏ?���?�������$������y ���7	��Sf߾�W征�� �k������S+���,��>�O?R8�?:��l&�>�r�E����$�����c8}>���=�Ð=��>�A�*�Q,�&,̾ݐG�QDʾS2�>��(>}�<�7?j�-?��?�HL?�S:?�s>݄O>��>z[K?�E>�0L?:�"?�":?+�A>�@>���>�!n<=	���h�����<�Ȧ�<��=���=mx�='�<��c�E�O�Y׽�s���z<��E�N�D���
=��Ǽ�t�=��?h�8?�d�}{}=E���B�p�8�=�N�>j*�=`kK�c�&>�d>���>3�?��>��>����{� � �4�2;}�?4�R??g?�|�=Z
�>a���$���5��L?>��;���X�|���W��'�o��>��o>�7�=��>���?�@�>إ?��<{�� �������C?�����þ��>|���R�3�\�e��K�&���g�� ��-C�F��>N�'>?�?���s=0�F>��t>^d>:QZ���=�0g>����ٸ�>$ �>5*�>oG�=5�>������h�9�]?�;ż����  ����UF����ޙG>�|�=\fN?�X�X�n��H���P<�a�>@��?�J�?�[?�VH�~~2�1O>>�2�>���>Z�>dD���k=��*�2T6>��<��4�����������=��=YB]�V)��sڲ��P�=Fڴ�YJB�^	��Þ��/)���۾5���n��a�P�V!\��F;L��Y�l��.�����Ty��놾f����y����?<,�?�Ό>bo> �A. �*�*���[��>��F�H�↾K96��ԏ�	���.���6����,���\��d����>��<�!���6)��n��� H,=����L?���S�D��3<��*��0�H=�L�����p�J"��L�žKua?0�??Y���������3?���?���>���=d�E��2w���?Q�=?�J?d�Z�2������O��=d,�?���?��??�O�D�A�o�����-?�?c��>u����;���K?'�9?S��>���g��f=� �>��[?�>N��b>��>0S�>S��Ώ��9�%�!/��rH����9>[�� ���*h�)	>�" �=��>gfx>3]�� ��I��>�'����`d�l�\��Ͼ����E�>�����J>^��=>�x>�;S��*���ѝ��G[�\tB?�h�?��A?g�d?&zR�r�O�K��=}��E�>�?C\>bF�����=s(�>O���hw������?���?�!�?�bY?b|��߿G������E�˾���=�ɓ=�m>|��<���=��j=8d�<$���8l>��>��>_j�>�.>Y>2d>I%��&z$����G���V�%�@���[�T����۾�,�ҋ澮���)䦾�1���Z�8��T<¡� ���s���1D�ë�=X� ?F�g>�`�>�L�>�]=��#�����p���ϑ�:$������;K��Zb�X�d���ھ[ޚ��|;�f�)��>�
�=
�;�|�>P3����>M�^>�V�>���=y'�=b]*>���>hh=�H>f��=��9>��=��>w+������0r��!M�rT�[[�; ~?�%C�ڝ����H�9�/�:ꤾ��>\RU?���>ě�����̭����h>�7>z@�<j53j��L>�`�>%5�<i��w:�&���Ѹ0���+>��>\==��h-��2w��ن�=�M�>ؾw=�=wk>��&?��w?ķ3?���=��>QMU>��>䓚=R(D>��E>�x�>щ?�U6?w+?L�>u��=KSg�=;=t{�=v�K�%?N�U֗���޲N�vv<��;�o6�<��n="��<�.+=�:=�U���;<lV�<&?�.?Yf�>?@�>mN��<�rE�u	:�_s0>p�#<Õ�>j��>W?���>�˷>1>�z���$ľT/¾[��>��,>;�W�G�r�N���>'��>�E?D�6?x���������<5�>���>�g�>�.?{S�>$�=�;�0����ֿ�	#�s�(���=�a�Ҽ��;�D ��ϼxu�<�'��*峽;`>=y^O><��>�~>��:>��3>\K>�&�>R{A>���=C �=��<��%�+Խ��׺I�L��}<�n��26�<v<��-��O���@�$�ܼ2�μ�����X?�J?�qý8w>U񌾙/���9ﾔyR<V�>!�>٫�>�Պ=���O9m�M�W����y�>��~?պ�>�Qj�f�5>Z�=:�����>��>,>W>	�z��`E��¾���>W��>���>V@e>��<�㐿�Г��;����>�������<�?:�>�}i�� ���E�$M�ȠD�7��>�ʐ��#���"��S%�֡F������/e��������?��s??������y��9d����i�t������>��>�9r>�fD=ԙ��� ���'��Ҿ`�h�F�0>e�?8�a��(Q?D\j?j�\?��,?��3?��d?���Y�?n��>��:??�?�XX?��B?Z��>�p�R��=��&>B�->�.�}�'�N��<f�l�
��<�m�=�a׼���;���'C�=�'=�X=�瑽}���f=�%�=2G;=nR>�} >P�?S�>`88�"]�W@Q�Jꬾl�o>�~�>_�=!�����ܾ�"þ���=gy�>�3?Ԭ�>G��g�(�q��b���%<�>�%?"�1?HL?�ɸ�4�>Ć!�8��݃��{O>@LF���ܾ)��`�Z�;��}�>�	!>O�����u>uQp?�15? {?P����	bc��/�H�޻�J9�y��>Ip�>
nF=���w�,��Iz�NTa�<z0���(�<3����;�>. =�y>B>>��>�1�=����˶<����H�H=�I�>F�>��?Cǃ>_�O<e��2���qS?��*��JO���(%����@����x�=o����>m�|�t���m�W:�QU>���?�H�?�e?�k���,���=t��=�&�>dW=�g�w�X�!>���>�)�=�4(�<á��>2�>Cw�>#�=���῾Z�'>:�̿je�Е�=���[�>�ƻ��[�&n��'�3�GE��A���8>;��/����-,���N��ϾE����	Y�?0��?�>��ƽc���tWݾ�_����z��	^F����lk=Ө�V����N����C����Q��U�>�ړr�����d�����b'���x�>�
���c�<�����L�=HȽRq����������G�޽!�]?q8U?��¾�:E�4}-��A�����=�;�>皃>T�=SO~��ߑ>�S?c/E?P)l��ڊ����Sn\���?_��?�V?�F��=��B-�1���� ?�?#�>�>�$������4?Pjl?M�?�� ��Ą��2�T�>�?OlF�_l>�E�>o�>���ψF��%�=���=�c=��O��R��;��A���V�=F�>�]�>k;�>um� �3�L�?fiҾM9��3PE�$@#�ϼ�"�x���E?�'�Ib(��W�>m��>*b-�Ӄ�����$=��b0?�ɳ?=�?�?�+u��;i�V;}S����!�&��>2<��(�|Ҏ>�B?k��֌��h&��I�>?��?�K@�͇?������ٿ�)���^پ��о�Ԭ=m��/�E>kr���	>��=ٵ_=1X���f=Z,�>#�a>�)>o��>�D2>De
>�e��C�!�"���ޔ�;B@�]�+����E!ڽ��n�>�y7�Ƶ�J���]/�=�X�࿕��o����R���/<N�2�ˢ+>,��>�D�=���>d��>:��>R���Td������&'���(��j�z�Ծ�������n���h��?��m�$��'?���=��%��h'?�z���=���>��>�_"=}��>��F>��>kt�>�=�>�a6=��.>�>P=���>ާ>�ᒿ
�M����6����j?Q����W��cM^�Aʊ���ھV!>N�>���>��S�ѥ��p��?�"�X�Ͼa����=r��>ʉ�>�m>A����=U���zž����d>2�>�!�<7ž�H/���&>�l�>��`�Ȣ�>�7�>69?���?��Q?2�=��>�M>���>��=I�>ݴ�>		?�
/?�^?B�U?/�>���<�5_�X=v��0\*�������3�兽ִ���R��� >A��=�m={� �Z�r>Ǎ>(K���=�=9x�<y��>�{f?���>�r1=rWӾW�0��Z�'T����=�=#@>$�?]��>-]�>��e>�sb>ae��m���a>�0?;[=�ד�X�����=�q/>��*>4}�?�c>?��>S3��]4�=Y3��ۨ> ?鯀?7��>�T>�N�=�����˿*�%��oP��־ф��0=qF�;x�3�'���s*=;\�
=0*>\�>��>"7>�,e>-B=O��=�;�>v�Q>���=Z>.�s<E@�=�|��;�g<���� �Ũ���; �<k�<�ν��X� �;���
Ks��?y!?��<�A�L��׽����4�U��>9\�>���>W�>�Z����@�H�X��%<�-�Z;8;?ȯY?k��>��Ͼ%U�;��K=S>>9?�^�>5��>�\��dま1�)�~�W��>C�C?g�>e!��S�{��pq��=��Li>���=��g��Ӏ?���?�������$������y ���7	��Sf߾�W征�� �k������S+���,��>�O?R8�?:��l&�>�r�E����$�����c8}>���=�Ð=��>�A�*�Q,�&,̾ݐG�QDʾS2�>��(>}�<�7?j�-?��?�HL?�S:?�s>݄O>��>z[K?�E>�0L?:�"?�":?+�A>�@>���>�!n<=	���h�����<�Ȧ�<��=���=mx�='�<��c�E�O�Y׽�s���z<��E�N�D���
=��Ǽ�t�=��?h�8?�d�}{}=E���B�p�8�=�N�>j*�=`kK�c�&>�d>���>3�?��>��>����{� � �4�2;}�?4�R??g?�|�=Z
�>a���$���5��L?>��;���X�|���W��'�o��>��o>�7�=��>���?�@�>إ?��<{�� �������C?�����þ��>|���R�3�\�e��K�&���g�� ��-C�F��>N�'>?�?���s=0�F>��t>^d>:QZ���=�0g>����ٸ�>$ �>5*�>oG�=5�>������h�9�]?�;ż����  ����UF����ޙG>�|�=\fN?�X�X�n��H���P<�a�>@��?�J�?�[?�VH�~~2�1O>>�2�>���>Z�>dD���k=��*�2T6>��<��4�����������=��=YB]�V)��sڲ��P�=Fڴ�YJB�^	��Þ��/)���۾5���n��a�P�V!\��F;L��Y�l��.�����Ty��놾f����y����?<,�?�Ό>bo> �A. �*�*���[��>��F�H�↾K96��ԏ�	���.���6����,���\��d����>��<�!���6)��n��� H,=����L?���S�D��3<��*��0�H=�L�����p�J"��L�žKua?0�??Y���������3?���?���>���=d�E��2w���?Q�=?�J?d�Z�2������O��=d,�?���?��??�O�D�A�o�����-?�?c��>u����;���K?'�9?S��>���g��f=� �>��[?�>N��b>��>0S�>S��Ώ��9�%�!/��rH����9>[�� ���*h�)	>�" �=��>gfx>3]�� ���Xj>�ݾs��!7e���/���ž��,>��U>�/?�:�=��->��F=�~A�����G`���O@<�Y8?�P�?^�D?΃a?�޾0��ư�~��$.?;�>Ou���������>�g.>*����i�5帾�d*?��?�O�?��R?1� ��ȿ�ј��Ҿ֐L���_>�g�;��>�����n9<۷�=�.E�����;*�N>�e�>@R�> <J>�=>��=�6z�h~$��f���y��%l'�u� �}�ae�6�1����ܸ���Ӿ�7���a��T�Cx��-<�֮e�����Kq�>X&?u��>\�>�v>l�=�a�"���Y��i���.2�������	������Y��}�%Z(��t��f|��N��V:�>h%=�|�m��>���=�So>�ν>��
>�$@>�r>�>��\���E=�=�7b>��>���=Rf�>TȚ=Y*��g��k&:��+�#�_=N?P�`��g��S���̾5l��sR>�W�>�N>��,�b����u�G�>c�мA�j�_������<�!�>���>�y=�S� ��<�(���
�a��=�m>�g*>���=�o_��&�E����>g����g=�Xe>VK ?��o?�K,?8�=��>#9�>�Q�>���=��K>�c<>K\j>µ
?�^9?D�0?SU�>�r�=�OI�6~�=jfV=�E��Է������T��Zf���D<"���"�=��u=d]T;���=NU�<�+�������=�L?���>��>M-?�u�& G��G<�Z�ɾ�b����=�kc>+�>��P?>�?��>׾�=����,+��T���>ڍ>�i��`��%��46)>&�?�h?� ?z?��̽�q~�5�;
�>+
?��?̾�=1��>k��=�H�^�Կ>�5ï��^>?����\������S�ǂ��J����^���}�=��Q>��7>��>@F>f)3=�ٳ><a�>3�=i(>���<�z+����T�&���Q=ݼ�=g�=�J�=����C*���"�������>��gO��n�̳	?	c?uϳ=R������ ^���Ǳ�(��>&��>�DZ?2A�>O�>���wKa���\�R�23�>3^?���>/ϔ�m��0�m�E��JL<�>��>�F>q���O^����>��?�6?�n�>e~�U�e��e�>u1��{>z��=���(�?'�M?�ྩ����D�{�i�-���=�m�qh��lѽ�T޾���w���b7��>#�����=0�?b(v?iZ��>ǝƾOÏ�?�p��,о�-��K>��	?�W?>X�z<ck��\���]��(x��0���,�>����<?��?|�J?�!:?XE�> �>S�C>bժ>����=P?@?b�=��C�E�a=��>���>�����Ҿ�N���P�%��=r�'=*m>��=�R��_Yp<��>6�Z�V=�@ ��p��>�ɼ�j����<	��=q�G="'?/
?'�s�x3=W��k=�н�>H�y=00=�s޼,�<��R=�Uj>B$�>)?N��=�Ѿu���ja���>���>m?[��>W���^�9/�/%��5�f>cg����<�����=
�����`6�JB�>���>�b>!�e>#�|?�oA?$_#?I� ��a,�qEs���)�c^�[Q���n�>+W�>�=�Rھoc3�1�m���W���0��t_��(F�%1=o*�=�)>�<>
�=J>�X2=ܯ���0�<��ټu�>��>-?ۢU>�YY=(���DQ����4?uv�����QF��
�V׹;X�o>���hO>_�>(D�����k.��pG���?l��?���?U�@?��=x�>>><���'��s�=�v>�،>� �����=��G>r�,�փ��SZ��r{5>̆?�?*�TD����j,�=nB��.#?��W��k\ľ�ع�Ӏ<��If�k�o��-��Fҽ���-�Hu�����Z1��R<�׾Z�ݾ~��R͓?��i?���>̹����0�á%�D˚�&s����W�`�;��<���.t�^s��e߾ ��&����$�o�оZ���O��>E#V���(���ݥ�ډ>[���� ?5�����i+�{�� �U>�J�>�Jx���j���T�ߢj?D"(?b���y ��ϔ>�O�>�?^ύ>�H�>�������c>�K?�N�?{��=ܟ��j���Oս��?���?Ms6?�hS��/>�o�۾���e?��>��>,�*�i;�H�ʾ���>��L?��?�t�J-��0Q��?��&?��$��3�>�l�>� ,=�rg�M-ڽӖ�=��0��·=�~:;te�<`�2��ܩ���f���=l��>TE�>mSо˭ �z�>(����
���d�",��Zj�<o=�N�>I>���S.>��>�
�;�H�穆���j��!E>Ib?�?�:?�?D�+�h����þ��Ƚ���>��>���<^0�����>�u�>����w�1(پd�%?)��?���?�&?i�&�Y̵��������R���u_�=� =-��=d��-ic>_u�=.��; ��E*�=3�\>��?>z��>Q c>+H>a�=�$��!4�"0�������k�������t��c����v�������z�ڶ�������=�ׄ������*��������>��}>|��>��>˾��͹>u���_G�@�<�/]��㾴���6��9"��������=8��=���*�<�G����?��L=�'�=���>,�ý���;���>F�ڽ{�_>�er>1�>��F=���=�+�<�ե=��#>��ٽa�>��u=O����f�	'����=����-�V?ܑ ��2������Ҿ�zɾ��=}�>��?>P/��ت��p���z�>��;�m�s%�=<`N�i~�=	#>� <>\&�6��<�;ڽ�P��X>�TC>��>�J�=kז=�Σ�q��&(�>��Ӿ���=ͷv>�'?��s?�6?�L�=�y�>B�d>u��>�з=)7J>(�O>u7�>��?��9?<2?���>	S�=+�\��+=)P=��=��T�������ǼRJ���q<i�'��(J=*�c==�;`�J=�y2= L��-c<��=���>C��>���>���>�g[��*=���^�{���Y*=t�h����>da�>.A)?�?ز>&#~=�����g������?�>`�p==|_�a�W�+r?��jf>�x�>A�m?je5?�V�D���@ݽI�#>S\�>ܢ�>�/?`l>���>�8��\�e|ѿBX%�� ��p}�G�3�r��;S:�LvM�|j;�w4�L~���<��Z>� �>�n>��F>��(>�=>Hk�>H�G>5X�=�ث=d�;�<e;1�O��M=e3ռ��;ݧ;�������Ƽҥ��x���kf�E>H��*���ۼ�?�_
?ٚ�=y��8*侮D0�����LX�>?bE?���>�~�>u� � �s��ti������^?4Ea?n$�>���;��<�茾�iǾ�y�>�S?*0]>gz�=e�Ƚh��[7�>��>��?$[�>�*��0�l��ۅ��!(��1 ?۶N=O��/w�?�V?�y�������,��d�����[h�ds�µ����q�3���±�K����^�Q��6>D�?��?qo?���=7D;9҉��偿���3j�=��m<'��><]b>�؇��m����S�ܾ{�V��� =��>��׾&�'?d� ?9�"?�f�?�Of>��>����"3<(��>�6?1��>Y�|>j��=�ei:ba=p^�>&�㽞Cоsfս��W�X�6>S����D>�>fZ�=W���9�=�4�<��%=�Z�MѼ�=���!C=���<V�=��=�	?���>Q��M�'>M|��qq�����\>���=�1p�.0l��lv=��>��>Զ?C:�>�==��ƾ����J�U�>$�?yE?pQ�>}傾����A��,���Ϙ>fA>��c�.µ��5�����H<q?(��>W�z>��^>�?l@?G�"?��D.�.ev��r(���߼�iͻNm�>w�>�њ=��۾!66��Sr�M\��/0��^�O�V�=+��=#q>�]L>�
�=s�>�?=�O����۽|	%;l/���t�>�6�>1�?@�Z>�=�N���N�Z� ?�G���\2�I��	�>��}>�!>}�=N�!?Y�vd��%﮿T'��.?^�?|��?,?2����?>ׇ9�g\E��6R>5�>A:�==�I��ڞ=�q�>�>��f����@�B�>Р�>JY�>!	����g��c�H��y���EF�+�B��Ծjݖ��߾VL���$��z��l����ޘ4���4����c��Xm5� D������R���$3�?)|?E�=}�˼X� ���b��0�5=`������>᜾�I-��!��ɭ�CК�2����#�_'�R��Б�>S����ڐ��Z~�M�m�>a��<�+?��)�����$��f��xH>�e�>RB
�r�}�����cQ
�� P?��,?��վi¾����v�NX�>?��>���=��׾��Ծ���F	N?��q?�H>{
�������P��Y�?a{�?ǷP?�M�Z�(������Ӿã�>C�K?�?����N:��Z��X��>�c?�U(?(Nὠ ��9m^�;�>B�:?ʵ ��[�>|I�=v��>��m<�혾�J>�y0���
�>x��Ϊh�	���-c���>��>^߮=��̾�1侮Xj>�ݾs��!7e���/���ž��,>��U>�/?�:�=��->��F=�~A�����G`���O@<�Y8?�P�?^�D?΃a?�޾0��ư�~��$.?;�>Ou���������>�g.>*����i�5帾�d*?��?�O�?��R?1� ��ȿ�ј��Ҿ֐L���_>�g�;��>�����n9<۷�=�.E�����;*�N>�e�>@R�> <J>�=>��=�6z�h~$��f���y��%l'�u� �}�ae�6�1����ܸ���Ӿ�7���a��T�Cx��-<�֮e�����Kq�>X&?u��>\�>�v>l�=�a�"���Y��i���.2�������	������Y��}�%Z(��t��f|��N��V:�>h%=�|�m��>���=�So>�ν>��
>�$@>�r>�>��\���E=�=�7b>��>���=Rf�>TȚ=Y*��g��k&:��+�#�_=N?P�`��g��S���̾5l��sR>�W�>�N>��,�b����u�G�>c�мA�j�_������<�!�>���>�y=�S� ��<�(���
�a��=�m>�g*>���=�o_��&�E����>g����g=�Xe>VK ?��o?�K,?8�=��>#9�>�Q�>���=��K>�c<>K\j>µ
?�^9?D�0?SU�>�r�=�OI�6~�=jfV=�E��Է������T��Zf���D<"���"�=��u=d]T;���=NU�<�+�������=�L?���>��>M-?�u�& G��G<�Z�ɾ�b����=�kc>+�>��P?>�?��>׾�=����,+��T���>ڍ>�i��`��%��46)>&�?�h?� ?z?��̽�q~�5�;
�>+
?��?̾�=1��>k��=�H�^�Կ>�5ï��^>?����\������S�ǂ��J����^���}�=��Q>��7>��>@F>f)3=�ٳ><a�>3�=i(>���<�z+����T�&���Q=ݼ�=g�=�J�=����C*���"�������>��gO��n�̳	?	c?uϳ=R������ ^���Ǳ�(��>&��>�DZ?2A�>O�>���wKa���\�R�23�>3^?���>/ϔ�m��0�m�E��JL<�>��>�F>q���O^����>��?�6?�n�>e~�U�e��e�>u1��{>z��=���(�?'�M?�ྩ����D�{�i�-���=�m�qh��lѽ�T޾���w���b7��>#�����=0�?b(v?iZ��>ǝƾOÏ�?�p��,о�-��K>��	?�W?>X�z<ck��\���]��(x��0���,�>����<?��?|�J?�!:?XE�> �>S�C>bժ>����=P?@?b�=��C�E�a=��>���>�����Ҿ�N���P�%��=r�'=*m>��=�R��_Yp<��>6�Z�V=�@ ��p��>�ɼ�j����<	��=q�G="'?/
?'�s�x3=W��k=�н�>H�y=00=�s޼,�<��R=�Uj>B$�>)?N��=�Ѿu���ja���>���>m?[��>W���^�9/�/%��5�f>cg����<�����=
�����`6�JB�>���>�b>!�e>#�|?�oA?$_#?I� ��a,�qEs���)�c^�[Q���n�>+W�>�=�Rھoc3�1�m���W���0��t_��(F�%1=o*�=�)>�<>
�=J>�X2=ܯ���0�<��ټu�>��>-?ۢU>�YY=(���DQ����4?uv�����QF��
�V׹;X�o>���hO>_�>(D�����k.��pG���?l��?���?U�@?��=x�>>><���'��s�=�v>�،>� �����=��G>r�,�փ��SZ��r{5>̆?�?*�TD����j,�=nB��.#?��W��k\ľ�ع�Ӏ<��If�k�o��-��Fҽ���-�Hu�����Z1��R<�׾Z�ݾ~��R͓?��i?���>̹����0�á%�D˚�&s����W�`�;��<���.t�^s��e߾ ��&����$�o�оZ���O��>E#V���(���ݥ�ډ>[���� ?5�����i+�{�� �U>�J�>�Jx���j���T�ߢj?D"(?b���y ��ϔ>�O�>�?^ύ>�H�>�������c>�K?�N�?{��=ܟ��j���Oս��?���?Ms6?�hS��/>�o�۾���e?��>��>,�*�i;�H�ʾ���>��L?��?�t�J-��0Q��?��&?��$��3�>�l�>� ,=�rg�M-ڽӖ�=��0��·=�~:;te�<`�2��ܩ���f���=l��>TE�>mSо˭ �z�>(����
���d�",��Zj�<o=�N�>I>���S.>��>�
�;�H�穆���j��!E>Ib?�?�:?�?D�+�h����þ��Ƚ���>��>���<^0�����>�u�>����w�1(پd�%?)��?���?�&?i�&�Y̵��������R���u_�=� =-��=d��-ic>_u�=.��; ��E*�=3�\>��?>z��>Q c>+H>a�=�$��!4�"0�������k�������t��c����v�������z�ڶ�������=�ׄ������*��������>��}>|��>��>˾��͹>u���_G�@�<�/]��㾴���6��9"��������=8��=���*�<�G����?��L=�'�=���>,�ý���;���>F�ڽ{�_>�er>1�>��F=���=�+�<�ե=��#>��ٽa�>��u=O����f�	'����=����-�V?ܑ ��2������Ҿ�zɾ��=}�>��?>P/��ت��p���z�>��;�m�s%�=<`N�i~�=	#>� <>\&�6��<�;ڽ�P��X>�TC>��>�J�=kז=�Σ�q��&(�>��Ӿ���=ͷv>�'?��s?�6?�L�=�y�>B�d>u��>�з=)7J>(�O>u7�>��?��9?<2?���>	S�=+�\��+=)P=��=��T�������ǼRJ���q<i�'��(J=*�c==�;`�J=�y2= L��-c<��=���>C��>���>���>�g[��*=���^�{���Y*=t�h����>da�>.A)?�?ز>&#~=�����g������?�>`�p==|_�a�W�+r?��jf>�x�>A�m?je5?�V�D���@ݽI�#>S\�>ܢ�>�/?`l>���>�8��\�e|ѿBX%�� ��p}�G�3�r��;S:�LvM�|j;�w4�L~���<��Z>� �>�n>��F>��(>�=>Hk�>H�G>5X�=�ث=d�;�<e;1�O��M=e3ռ��;ݧ;�������Ƽҥ��x���kf�E>H��*���ۼ�?�_
?ٚ�=y��8*侮D0�����LX�>?bE?���>�~�>u� � �s��ti������^?4Ea?n$�>���;��<�茾�iǾ�y�>�S?*0]>gz�=e�Ƚh��[7�>��>��?$[�>�*��0�l��ۅ��!(��1 ?۶N=O��/w�?�V?�y�������,��d�����[h�ds�µ����q�3���±�K����^�Q��6>D�?��?qo?���=7D;9҉��偿���3j�=��m<'��><]b>�؇��m����S�ܾ{�V��� =��>��׾&�'?d� ?9�"?�f�?�Of>��>����"3<(��>�6?1��>Y�|>j��=�ei:ba=p^�>&�㽞Cоsfս��W�X�6>S����D>�>fZ�=W���9�=�4�<��%=�Z�MѼ�=���!C=���<V�=��=�	?���>Q��M�'>M|��qq�����\>���=�1p�.0l��lv=��>��>Զ?C:�>�==��ƾ����J�U�>$�?yE?pQ�>}傾����A��,���Ϙ>fA>��c�.µ��5�����H<q?(��>W�z>��^>�?l@?G�"?��D.�.ev��r(���߼�iͻNm�>w�>�њ=��۾!66��Sr�M\��/0��^�O�V�=+��=#q>�]L>�
�=s�>�?=�O����۽|	%;l/���t�>�6�>1�?@�Z>�=�N���N�Z� ?�G���\2�I��	�>��}>�!>}�=N�!?Y�vd��%﮿T'��.?^�?|��?,?2����?>ׇ9�g\E��6R>5�>A:�==�I��ڞ=�q�>�>��f����@�B�>Р�>JY�>!	����g��c�H��y���EF�+�B��Ծjݖ��߾VL���$��z��l����ޘ4���4����c��Xm5� D������R���$3�?)|?E�=}�˼X� ���b��0�5=`������>᜾�I-��!��ɭ�CК�2����#�_'�R��Б�>S����ڐ��Z~�M�m�>a��<�+?��)�����$��f��xH>�e�>RB
�r�}�����cQ
�� P?��,?��վi¾����v�NX�>?��>���=��׾��Ծ���F	N?��q?�H>{
�������P��Y�?a{�?ǷP?�M�Z�(������Ӿã�>C�K?�?����N:��Z��X��>�c?�U(?(Nὠ ��9m^�;�>B�:?ʵ ��[�>|I�=v��>��m<�혾�J>�y0���
�>x��Ϊh�	���-c���>��>^߮=��̾�1侌��>��꾰nJ���G�l	�$�#����<f  ?Ik쾑�>��b>�K>��(������凿�@򽣮K?���?�8Q?";?�����w�x�ý�Ɛ=A �>!n�>S��=���A�>�W�>D��,�p�S.�W6?�c�?�a�?�\Y?��l�>Gӿ��"������	��=%�=��>>��޽�ɭ=��K=ʘ�hZ=�n�>��>o>:;x>w�T>Л<>��.>p�����#��ʤ�4ْ��[B�� ���wg��{	��y�����ȴ���O�������=Г�}�G�^���T>��־$b�>zk?M�n>��>Đ�������r�'ƾ��=�XJ��˾���+� ������������U3;�YﾋN���y���?]`Ӽ�ae<+�w>��;�?��Ć>�X�<�>|�<W�p=d}J>�'�><I�>_��>wr�>Myڼ?Y>a�y���\����-
4�Cr-��w�=ɓ ?��;�㶾S�4��/�u����i�>�pM?���>�j�KL��E�Y�`e(?��A������q�X:>�?�ķ>#�/>	�:�aF��LH�wi���6>�T?�>\/�@����K[�v��={�>�ʾ�(�o�B>��$?-e?��?�DK��?Q�>�H1>�<g=H�t>th>��
>�>sO0?��:?���>y�=�d���N!>�-�k����:�)@�i��������Ӂx=�9��=�Պ<LFZ=�0�=K���hD������>PZ?8�	?�>�?����S�O�L���� K���q�h�=w�>e��>pb�>w��>e�>v'�<u�v��꡾.R?�/1<Me�E=�j]���h>h�><ߍ?'I+?D:�>�[����3s>��f>¸�>�?���>r�x>��f��7	�*zҿ6!�h!�B����$�Dv��?�A��nI�$�.�,�.������<#DS>���>qBh>�6?>�>�~3>�r�>8�H>=�=���=.9V��l�;�?��SO=�q��T�<ݙZ��K(�Rfϼ�����Ջ5�Ԟ.�������R/?A�>��ƾ�v���ț=qY�ת����>&��>ԏ�>�g?n��>}��R�C�r��")��M?� �?��>)ui�=h=�[7��m���� ?0�;>A� ��j���S��������0�>�W?H�>�����E��򛙿E09��@?���='�-�-<�?\"O?�����F��X�n�����$����J����u�M��b���޾4� ���\��=���>6N�?��4���*>)�������}������qܽo�A����>u$l>v%������A=��,����n&<`��>��z���?��H?��>,-`?Ɠ�>��,>(��>��Z>@�>0�.?�F�>�|L<��׼'WX>�P�=?,�>�bξ�{��<�p�Z���a�J=~;����=�>%��<;`I=���=|<D�B�������EϹ=[<�"�;yG�=���ї=ȯ�>G��>���>������>:þ=3��g�����D��VИ�����z��$�{>{�?|3?\��>�=���<p�<��-�t,�>�
$?��>�-�>�����¸��v�,T�h�B>���=X㫽�/���F��\X�:��=�.?Z��=�#�z�I>�Ó?�?q ?�� =�9%���U�r,���T�$>c��>.�n>�Y	��@�)�*���|���=�u5j��沾Pλ�\�>��w>�M>�S>JI<��=�/��׽��8=��I<z�w��ud>T{�>�?�>�,w>�Lf�����S?�s�����R,��Z���K�<t'�>�>m>VF??R���{�u����_��ˮ>�e�?uu�?��^?N@Ǿ��=��$={s)�co��M��>�=�+>�[:=��B>�1�<'��>[����kv�G��=����y�5��}h��ѹ��/�?�ֿ��O�:��=A�)��=�^1�|.޾�
�����=օ����M᷾�o�>��4���U��Y��AM���C���?�T?b�^>��ǽ7�#�t

�(�_�ق���m+�s����Z�����S���`�6��o��CN��Ҿu�����>�H��	����y�֙��nh>��">s	?G�Y�b徯�(�u��O�>���>��/��;M�ˆ��l�<#R?��:?�3�(c&����>i�>�,�>M�>�gm>P㾈�׼t����\?�_�?�7m=f��yС���o��k�?̳�?zbQ?��E_�(�^� �߽���>*�E?휕>v��f]
�䤞�y�$?6k?�?���k�R�.4�M��>�dM?2v�U�"?}^>j��>V�վ)*_�{]�=\���n��dQ=n�����)���ž��S���!>�7>L�j>���Ͼ~��>?<�&��l�J���)�?�����d>�t�>����s?�JL>��W�=z8�	H����m��R�Ǽ�?��?�)�?eL�?�@�X\`�gj�p��> dD?��>C��>ā��L�>ap"?-�Zr���i���>��?z�?%N?��U�>Gӿ��!������	��=%�=��>>��޽�ɭ=��K=�ɘ�*Z=�n�>���>o>D;x>w�T>ϛ<>��.>r�����#��ʤ�4ْ��[B�� ���wg��{	��y�����ȴ���K�������<Г�y�G�^���T>�@�����=�H�>
Rg>���>��>R��>)���9�J��$�����v���<�
6���ԧ�E�<�e�C��+վ�.Q���վT�?��f=-����>��k�>�=�1�>���=E�>4�=�<�=���=X�:>���=�"�=�O�>�h��{��>.T�O����6z��;�6ü	/k>�dP?��#=y���	�?��vʾ�J�V��>�]N?_*�>p3�r󙿧�E�ԊP>��<y���vZL����Fr>F��>�&K�08>���;�H��̡=�u�=�.�>��>(۠=ud��r��$N>L�>��Ծ���=y�u>hw(?��v?>�4?=p�=m�>9^>{��>���=�G>��N>T8�>52?ӽ9?w1?1��>���=]�]���=D09=��=�e�`�[����Xἤ���E�<!�5�I�:=��|=r�;ܬU=��;=@󹼞�<�=��?��?���>=2?�!�`����6�8}�>��=5Uv��?;�?�2?�S?���>YJ�3Ǡ�V'T��떾E.?�&l��Q���Њ��J���w�=�?�Y?pa?� ȾD�־ixN>'��>-0?��?e�?����ӏ=���A��bҿ�{�d<������	���<Hj��]�6��0>!�B��o�<c�>r�u>xV>�C>�J(>��7>�4�>���>�k�=h��=2=����Ƽ ]z�g�<d����<{R���5=)���<�G�Ž��۽ʨs�JqA�𡷽��>��7?���=d܄�0rT<�M����/��D$>�?�%>Wu�>�5����ξL]� �z�e�
�O�>�B�?�5�>c�!� =��d<��m�N>��t>eW4<�}����)�n�x���>h5?�<?F�=�<��8o���w�yEؾ��>^]��� �RH�?<Bn?��L�����R�Εi�V�z\u>�v����I�yD8��e#�y�Ͼ�.�O��U�ܾ��;���>O�A?�K�x�<c��P�l�ܪ9�����O>*,�m�
>�NٽС������4�@G���Κ=��>�|)?�+ؽN,+?t��>V?i}x?��>��-?�W�T�1?o0����I>I$?�?��1?@��>�HA>8���<�
D>!Ws�᏾���;��ɽ]<�h�>?;6>���-">����<4��g�����=��n=A�=>ax��Q�=�F>
�?&��>�\󾛖w���>�`�� [>�>�i\>�9�yw��>d�>H�3?%M?�p�>i�лM��`e���T�cO	?`��>��?�J:?]J���4�O�*����wH#=���>�嚽�U���7�-�;��g��>h�>�� =n�>k�r?lsR?
?�l��hž="���l��H���N ���>�>��>֌�JZ��;j���=�L�Ҿϥr>��s�U���>E\?ܵ'>��G>���=��>r����H�=&�t=)��=w_�>S/�>�?T�=y>ھ�Gž�Y?��.A�-]���ٽr�>l>��z><]I�Т�>�5>m׈�!_��.� �i�
?��?*S�?�>?��þc-�� g>�5>h>0q��Z���J�A�����>�,h;��ݾ:����>���>���>��)�~ پ���đֽ�bҿA�#�x .>�3��>��$�����?R�ر;>��m����R	���h=�L����6��Ⱦn��sq�?�?�u�>�J�=(�X�A�+��A�����[���nT;>����C��<�5���b��Y�8��B��D�5�>��Hʛ>5�X��.���|��(�Aꓼ2?>*/?Eƾ|Ҵ�����k=�%>t�<5�˟��ڐ���p
��W?b�9?T�����<�,p>(�?���>��%>�[��6\�U�>J4?=�-?3�����::������j�?�	�?d�=?HT���YP����w>�Xղ>�q?�?��E��g �+ �œ?��N?��?�<�)y�Y�	���?"I:?� ��k�;>v��>%�>�Pƽ|����>P���}���]�>D�kK�g刼٬����=��X>^�b>�T��f�E�~��>?<�&��l�J���)�?�����d>�t�>����s?�JL>��W�=z8�	H����m��R�Ǽ�?��?�)�?eL�?�@�X\`�gj�p��> dD?��>C��>ā��L�>ap"?-�Zr���i���>��?z�?%N?��U�>Gӿ��!������	��=%�=��>>��޽�ɭ=��K=�ɘ�*Z=�n�>���>o>D;x>w�T>ϛ<>��.>r�����#��ʤ�4ْ��[B�� ���wg��{	��y�����ȴ���K�������<Г�y�G�^���T>�@�����=�H�>
Rg>���>��>R��>)���9�J��$�����v���<�
6���ԧ�E�<�e�C��+վ�.Q���վT�?��f=-����>��k�>�=�1�>���=E�>4�=�<�=���=X�:>���=�"�=�O�>�h��{��>.T�O����6z��;�6ü	/k>�dP?��#=y���	�?��vʾ�J�V��>�]N?_*�>p3�r󙿧�E�ԊP>��<y���vZL����Fr>F��>�&K�08>���;�H��̡=�u�=�.�>��>(۠=ud��r��$N>L�>��Ծ���=y�u>hw(?��v?>�4?=p�=m�>9^>{��>���=�G>��N>T8�>52?ӽ9?w1?1��>���=]�]���=D09=��=�e�`�[����Xἤ���E�<!�5�I�:=��|=r�;ܬU=��;=@󹼞�<�=��?��?���>=2?�!�`����6�8}�>��=5Uv��?;�?�2?�S?���>YJ�3Ǡ�V'T��떾E.?�&l��Q���Њ��J���w�=�?�Y?pa?� ȾD�־ixN>'��>-0?��?e�?����ӏ=���A��bҿ�{�d<������	���<Hj��]�6��0>!�B��o�<c�>r�u>xV>�C>�J(>��7>�4�>���>�k�=h��=2=����Ƽ ]z�g�<d����<{R���5=)���<�G�Ž��۽ʨs�JqA�𡷽��>��7?���=d܄�0rT<�M����/��D$>�?�%>Wu�>�5����ξL]� �z�e�
�O�>�B�?�5�>c�!� =��d<��m�N>��t>eW4<�}����)�n�x���>h5?�<?F�=�<��8o���w�yEؾ��>^]��� �RH�?<Bn?��L�����R�Εi�V�z\u>�v����I�yD8��e#�y�Ͼ�.�O��U�ܾ��;���>O�A?�K�x�<c��P�l�ܪ9�����O>*,�m�
>�NٽС������4�@G���Κ=��>�|)?�+ؽN,+?t��>V?i}x?��>��-?�W�T�1?o0����I>I$?�?��1?@��>�HA>8���<�
D>!Ws�᏾���;��ɽ]<�h�>?;6>���-">����<4��g�����=��n=A�=>ax��Q�=�F>
�?&��>�\󾛖w���>�`�� [>�>�i\>�9�yw��>d�>H�3?%M?�p�>i�лM��`e���T�cO	?`��>��?�J:?]J���4�O�*����wH#=���>�嚽�U���7�-�;��g��>h�>�� =n�>k�r?lsR?
?�l��hž="���l��H���N ���>�>��>֌�JZ��;j���=�L�Ҿϥr>��s�U���>E\?ܵ'>��G>���=��>r����H�=&�t=)��=w_�>S/�>�?T�=y>ھ�Gž�Y?��.A�-]���ٽr�>l>��z><]I�Т�>�5>m׈�!_��.� �i�
?��?*S�?�>?��þc-�� g>�5>h>0q��Z���J�A�����>�,h;��ݾ:����>���>���>��)�~ پ���đֽ�bҿA�#�x .>�3��>��$�����?R�ر;>��m����R	���h=�L����6��Ⱦn��sq�?�?�u�>�J�=(�X�A�+��A�����[���nT;>����C��<�5���b��Y�8��B��D�5�>��Hʛ>5�X��.���|��(�Aꓼ2?>*/?Eƾ|Ҵ�����k=�%>t�<5�˟��ڐ���p
��W?b�9?T�����<�,p>(�?���>��%>�[��6\�U�>J4?=�-?3�����::������j�?�	�?d�=?HT���YP����w>�Xղ>�q?�?��E��g �+ �œ?��N?��?�<�)y�Y�	���?"I:?� ��k�;>v��>%�>�Pƽ|����>P���}���]�>D�kK�g刼٬����=��X>^�b>�T��f�E�j�>7���;�PBl���@�=���ԑ>ݑ?�/��C�#?rp�>�!>�R����}ʄ�+���7��?��?�x?��|?��J�Na~�K��q�>��?^[�>)c�>����V�>��,?
�A��-���ؐ�N}?���?U��?��v?�];�yڿ	웿Q,���o��H�j>�=>j��=w�I�|��=T=>�
��<����=!�>l�`>Z��>�d>JdS>3�s>f܃�o�%��?��=��{-������)�gT�����D����"�ػɾ�)Ǿ���<+��E���fYԽ(�;��,~��e �='�\>�C>V�>�?�>��a>����#���i��uξ��H�k�+�%�侾����P�%&���������$�ٽڅپ���>)�=���<'G�> ��?,|>2�>�f.=g��>�eL>sڜ=œ�=v~�=�o4>y	>)~>@Bj>s��>�.�.z����NO�h���GA>^B?��󽖮���'f�~���-������>�M?��>������m"E����>,�>��/�H�N��^H�#�!>��>;�6��D=�#�'����>��<|s�>Z�������x����*��؄=G�>i*ϾɗԼ���=��!?�s?k-?X��=��Y>��>���>0�ȼ˧�=@?>l��>��?F�&?x�?���>Nڬ=̘���]%>OVJ=�!|�,P�<'.Y���Q������;?�=�G�<�e>���ˆ���m���)���= ���S	?�[4?��>�C�>S��bP�>冿��>YU�>� �t֏>�!�>�{E?���>��>H	E�̌���d�r��<�?q�^>N��>������=L�=���>�7f?m�?$�ݼ�"�(>c��>��*?��?8;c?P��>K8�>��5�q{�'�Կ�-��A���b;�G=R�'�]o��󡺽�"��A}���1���:<���>k��>�t�>kej>�>%>em>�\�>`(�>�%>���=D �K�M����;�?=�n�����ߺȹ=aJ�ʺ�P�J�	�'���E ���'k��?��?�
��K���D=��#��ؑ�����>���>���>���>z�;>����J�o�8�)Q�c�>
�v?���>?J���=6��K�q=7è>��a>=T�>�㿽G�:��.��a,�;�|�>M?��>�1��Ha���d�=����>���.��ۄ?#0?��K��v���w�[�H������I��{���d�y�L��oH���J�mRI�����F�����>2I�?����Q������;��T=��x���>�Q@>�C�>"R�>zC�_��!�>�"^��ط	��00>u�X?X˃��?Γ?v?��?��?6�/?K����K?X�\�LN�>�h#?�6?��??�4>Q�>㑷>O�=��>���eԇ���=aj�<'�=s�,>v��=�t��"`���>ی=�`����3�����'���<�=�$=���;֤=̦(?m?�|�
�ž%=I���F�=y�>�>?�����d�>�`�>^?�80?)��>�{7>��S���پӜ�3n�>�C�>�;?+�<?)�=1�>��1����5�0=al�>*D���ؾqx�?��ٯv���A>��>���=��F>G�t?�@?E��>�h���
��*����2���]4��;?~����Z�<��c����{|�i�n����]"�=�X��D�æ>-�>�4a=Y��=�n�>���w5~;n\�< ��<=�>P��>d�?/W׼����hZ��.�ξF�s?��H�{�`�����b��B��>�M�>�k�>�ٿ�4?��=�Ђ�~~���� ���1?���?@�?D:\?�;��Ký���>�;>>��>Y��U���D<,����>c�?=h4�G� ��V�>�)?�:5?��'�<�8�W�\��6�)���%t(��>Y>��޽KY۾/�޾����@
�Σܾۤ��wJ���$��!ʽ:M]�|o��#� ���׾���5L�Xz?�q?7��>r�*>]+S�m������伎�
����!4��$�	��Ɨ��U�{i��t#'���A��F#�M�;���>��Y��
��HJ{��W*�ɢ��'�=><�-?�žT鸾��vP=�z >@p�<S��x&����%���U?��9?���p;��my޽)!>�
?R��>�&>�����Y�⦒>S�2?v�,?���ʎ����閼]3�?���?V�??����=������ʩ����>��
?=��>�q���޾���v*?��5?� �>��q���r���?�|G?�ヾ��E>z:�>�>����P骾���=��۾��˼z��=;t��5=��8��0ؽB��=��|>Dj�>�%��J���~��>?<�&��l�J���)�?�����d>�t�>����s?�JL>��W�=z8�	H����m��R�Ǽ�?��?�)�?eL�?�@�X\`�gj�p��> dD?��>C��>ā��L�>ap"?-�Zr���i���>��?z�?%N?��U�>Gӿ��!������	��=%�=��>>��޽�ɭ=��K=�ɘ�*Z=�n�>���>o>D;x>w�T>ϛ<>��.>r�����#��ʤ�4ْ��[B�� ���wg��{	��y�����ȴ���K�������<Г�y�G�^���T>�@�����=�H�>
Rg>���>��>R��>)���9�J��$�����v���<�
6���ԧ�E�<�e�C��+վ�.Q���վT�?��f=-����>��k�>�=�1�>���=E�>4�=�<�=���=X�:>���=�"�=�O�>�h��{��>.T�O����6z��;�6ü	/k>�dP?��#=y���	�?��vʾ�J�V��>�]N?_*�>p3�r󙿧�E�ԊP>��<y���vZL����Fr>F��>�&K�08>���;�H��̡=�u�=�.�>��>(۠=ud��r��$N>L�>��Ծ���=y�u>hw(?��v?>�4?=p�=m�>9^>{��>���=�G>��N>T8�>52?ӽ9?w1?1��>���=]�]���=D09=��=�e�`�[����Xἤ���E�<!�5�I�:=��|=r�;ܬU=��;=@󹼞�<�=��?��?���>=2?�!�`����6�8}�>��=5Uv��?;�?�2?�S?���>YJ�3Ǡ�V'T��떾E.?�&l��Q���Њ��J���w�=�?�Y?pa?� ȾD�־ixN>'��>-0?��?e�?����ӏ=���A��bҿ�{�d<������	���<Hj��]�6��0>!�B��o�<c�>r�u>xV>�C>�J(>��7>�4�>���>�k�=h��=2=����Ƽ ]z�g�<d����<{R���5=)���<�G�Ž��۽ʨs�JqA�𡷽��>��7?���=d܄�0rT<�M����/��D$>�?�%>Wu�>�5����ξL]� �z�e�
�O�>�B�?�5�>c�!� =��d<��m�N>��t>eW4<�}����)�n�x���>h5?�<?F�=�<��8o���w�yEؾ��>^]��� �RH�?<Bn?��L�����R�Εi�V�z\u>�v����I�yD8��e#�y�Ͼ�.�O��U�ܾ��;���>O�A?�K�x�<c��P�l�ܪ9�����O>*,�m�
>�NٽС������4�@G���Κ=��>�|)?�+ؽN,+?t��>V?i}x?��>��-?�W�T�1?o0����I>I$?�?��1?@��>�HA>8���<�
D>!Ws�᏾���;��ɽ]<�h�>?;6>���-">����<4��g�����=��n=A�=>ax��Q�=�F>
�?&��>�\󾛖w���>�`�� [>�>�i\>�9�yw��>d�>H�3?%M?�p�>i�лM��`e���T�cO	?`��>��?�J:?]J���4�O�*����wH#=���>�嚽�U���7�-�;��g��>h�>�� =n�>k�r?lsR?
?�l��hž="���l��H���N ���>�>��>֌�JZ��;j���=�L�Ҿϥr>��s�U���>E\?ܵ'>��G>���=��>r����H�=&�t=)��=w_�>S/�>�?T�=y>ھ�Gž�Y?��.A�-]���ٽr�>l>��z><]I�Т�>�5>m׈�!_��.� �i�
?��?*S�?�>?��þc-�� g>�5>h>0q��Z���J�A�����>�,h;��ݾ:����>���>���>��)�~ پ���đֽ�bҿA�#�x .>�3��>��$�����?R�ر;>��m����R	���h=�L����6��Ⱦn��sq�?�?�u�>�J�=(�X�A�+��A�����[���nT;>����C��<�5���b��Y�8��B��D�5�>��Hʛ>5�X��.���|��(�Aꓼ2?>*/?Eƾ|Ҵ�����k=�%>t�<5�˟��ڐ���p
��W?b�9?T�����<�,p>(�?���>��%>�[��6\�U�>J4?=�-?3�����::������j�?�	�?d�=?HT���YP����w>�Xղ>�q?�?��E��g �+ �œ?��N?��?�<�)y�Y�	���?"I:?� ��k�;>v��>%�>�Pƽ|����>P���}���]�>D�kK�g刼٬����=��X>^�b>�T��f�E�~��>?<�&��l�J���)�?�����d>�t�>����s?�JL>��W�=z8�	H����m��R�Ǽ�?��?�)�?eL�?�@�X\`�gj�p��> dD?��>C��>ā��L�>ap"?-�Zr���i���>��?z�?%N?��U�>Gӿ��!������	��=%�=��>>��޽�ɭ=��K=�ɘ�*Z=�n�>���>o>D;x>w�T>ϛ<>��.>r�����#��ʤ�4ْ��[B�� ���wg��{	��y�����ȴ���K�������<Г�y�G�^���T>�@�����=�H�>
Rg>���>��>R��>)���9�J��$�����v���<�
6���ԧ�E�<�e�C��+վ�.Q���վT�?��f=-����>��k�>�=�1�>���=E�>4�=�<�=���=X�:>���=�"�=�O�>�h��{��>.T�O����6z��;�6ü	/k>�dP?��#=y���	�?��vʾ�J�V��>�]N?_*�>p3�r󙿧�E�ԊP>��<y���vZL����Fr>F��>�&K�08>���;�H��̡=�u�=�.�>��>(۠=ud��r��$N>L�>��Ծ���=y�u>hw(?��v?>�4?=p�=m�>9^>{��>���=�G>��N>T8�>52?ӽ9?w1?1��>���=]�]���=D09=��=�e�`�[����Xἤ���E�<!�5�I�:=��|=r�;ܬU=��;=@󹼞�<�=��?��?���>=2?�!�`����6�8}�>��=5Uv��?;�?�2?�S?���>YJ�3Ǡ�V'T��떾E.?�&l��Q���Њ��J���w�=�?�Y?pa?� ȾD�־ixN>'��>-0?��?e�?����ӏ=���A��bҿ�{�d<������	���<Hj��]�6��0>!�B��o�<c�>r�u>xV>�C>�J(>��7>�4�>���>�k�=h��=2=����Ƽ ]z�g�<d����<{R���5=)���<�G�Ž��۽ʨs�JqA�𡷽��>��7?���=d܄�0rT<�M����/��D$>�?�%>Wu�>�5����ξL]� �z�e�
�O�>�B�?�5�>c�!� =��d<��m�N>��t>eW4<�}����)�n�x���>h5?�<?F�=�<��8o���w�yEؾ��>^]��� �RH�?<Bn?��L�����R�Εi�V�z\u>�v����I�yD8��e#�y�Ͼ�.�O��U�ܾ��;���>O�A?�K�x�<c��P�l�ܪ9�����O>*,�m�
>�NٽС������4�@G���Κ=��>�|)?�+ؽN,+?t��>V?i}x?��>��-?�W�T�1?o0����I>I$?�?��1?@��>�HA>8���<�
D>!Ws�᏾���;��ɽ]<�h�>?;6>���-">����<4��g�����=��n=A�=>ax��Q�=�F>
�?&��>�\󾛖w���>�`�� [>�>�i\>�9�yw��>d�>H�3?%M?�p�>i�лM��`e���T�cO	?`��>��?�J:?]J���4�O�*����wH#=���>�嚽�U���7�-�;��g��>h�>�� =n�>k�r?lsR?
?�l��hž="���l��H���N ���>�>��>֌�JZ��;j���=�L�Ҿϥr>��s�U���>E\?ܵ'>��G>���=��>r����H�=&�t=)��=w_�>S/�>�?T�=y>ھ�Gž�Y?��.A�-]���ٽr�>l>��z><]I�Т�>�5>m׈�!_��.� �i�
?��?*S�?�>?��þc-�� g>�5>h>0q��Z���J�A�����>�,h;��ݾ:����>���>���>��)�~ پ���đֽ�bҿA�#�x .>�3��>��$�����?R�ر;>��m����R	���h=�L����6��Ⱦn��sq�?�?�u�>�J�=(�X�A�+��A�����[���nT;>����C��<�5���b��Y�8��B��D�5�>��Hʛ>5�X��.���|��(�Aꓼ2?>*/?Eƾ|Ҵ�����k=�%>t�<5�˟��ڐ���p
��W?b�9?T�����<�,p>(�?���>��%>�[��6\�U�>J4?=�-?3�����::������j�?�	�?d�=?HT���YP����w>�Xղ>�q?�?��E��g �+ �œ?��N?��?�<�)y�Y�	���?"I:?� ��k�;>v��>%�>�Pƽ|����>P���}���]�>D�kK�g刼٬����=��X>^�b>�T��f�E�&��>�G���N�֧H�U��������<��?�}�4>#i>^Y>F�(�����ʉ��3��L?���?��S?ah8?6c��Լ�F}��ށ�='��>߿�>���=�����>M�>Tb�{r����?SD�?���?�bZ?��m�=�ſ�r�����=�ƾYɯ=�9	>�h�>���<�8��HG=��&=[��=�7�=��>	an>k�O>���>�!|>l`��6���#�p������BnA�x
���.�ܣ�����O�a�^F�޼��c��]��$Z�F"��˂�q>���*��־L^����>�l><v�=�4A>س:>(B��'����Z0��#���%:�?���Z�éƾ�ݪ�����&9ҽL'=4"���?V��=�V��� ?������=���>%��=�~�>^�k8���>�R>��>���=���>��n�(*n>!�<�j��.���r�?�;���IK�=��>?�᥾�}Z�E�7�ttվ���R>v>@&��Z]7�W*��W)B�X�>��Л���ꣽ+:>�%�>��>p�<*<�eJ���<4�<������l�>�)>15�=���C�b�$�=O�?��M�k߬>�#�>L�1?�Ë?�1Q?G�>�>$>!=��^>>5A7>]�	?w�?B~e?�l?[j~?���>P?�={N�R�=S�="��Hwy�3����!�	X��´>!�N>쓌=Ư�;<��=�X��?Q>.jA���&�=�{?�RT?���>$��>%�j=˚>�s}\�pg}>B�S=iV?�>���>A��>\��>�\�>��L�EJ��C��ϣ>�_�>K@G��f��佗^��1�>�V?��.?&����r���QU>b�z��>�1?ol�>��>CL�>�YA�(����{��g�&�����n��>�	����a�]�H>�=�u�2t���u�@�u��h5>��>����dhd>�t>z�f;�	�>�r>R�=�X-=�I��	/��X&��x�::�������a%��i���6d>�n��3�����>�q=�&��,��=BV?
�??��]ヽ��R��9�F'����>0 ?a��>�}�>l`�=������F�
a"� ��Qc?�F{?���>5�)�<p�=������G�>�o�>� *>��I�Q�1�6Ѿ�;=r��>�O1?2˖>^K�9�T�+9n�%V��>�%�=�?L���?�Oy?�.���/<0\� '|�� ����>���>�m�$E��V�H�˨T��Qھ�$��y��=z>N^�>�:�?A�۴�=f���j��m˂�_+&��G>�1?)[�>ZH/>M�.>9�DY��>���*�ʼ�`�r�v>�s>r�>9=? h6?��W?oiJ?�1&?��e>�lB>�躽�H�>�*�>�ʼ>�/?3�#?.�?�?qƂ>kB��V�н�r��A=>�7�<o`�=�f>+a�=��=�ĥ��S>Z$=8g�	��<��=���=>x4>d�=	S�=I.�=��?�(?��ȼ!�=.���V�ýfK=
�	>��1>��4��	�J�(=_�x>�-?��9?B+�>%�^>N�о�����ď�_o	?1h>?ɠ�>�]�>�@�>
̷��Ñ�A��=@�d>�P���?��7� �@M��ʢC�y�><��>��=Wҿ>P��?u4?׈�>2\f>` W�#ў�h�@�:)>:�	��%�>j�+?9t8=��\
�9oK��sZ���¾�T���[��C�=�>G�G�ΐ�>�z�=%�z���f>l�	> ���mo����j��>�E|>17I?WO>���=��e������I?��o���l9��l�����~���:>tO�>��&<��?9.7��+w��*��2,�t��>�{�?���?�t?����e��-m>�t0>X]�=lի;	����O<MS��H>�֗�ꄾ��f�n}O=�$>V>����=���^��=ء�����}�����=��f�"���{��� >7�D>�t��\�W,����eV���L�:�d���%�x&��	G�ǋz?Y}f?��>�^=�,;1&۾�cs���=������D�v�оi4#�'G��I���;�� (��3���'��������>Nٽ|�������9����� �>��?e������R��������>�X�+;�u����0�����U?��<?�w��型�S�>��?��?L[�>�s��/����g<q�?A?f�=��s��Oc�����?�ұ?�H?��(Y�r�#�B-�=y��>"V$?oZ�=u�_k߽�6����M�� ?2$��L{c���;��b�t-�;�{�?>�x��t>��?�#�>����c���5�a-�����:�>\"9�>�㙾�H���=��>�MC>�� �V_b�I��>��n7H�u�J��?�O�F�k�˼Z�>D@��2U>��q>��0>�� ��)��U���s�8�,F?벬?g:T?�9?�D(��/z���A/=���>7h�>�;>��׽���>AS�>����9jd�(��|C?���?yF�?]�W?�*j���Կ{㑿{�׾-��غ���>��>��>̓�=$O ��߽^7>�(g>�N�>��=�R >�8M>��G>�z%>6�����ʬ��i����a�B� ��������'�����>�=�B����;�w�8��Po���@�R���_c~�&M�=�/��/+�E�>��>���=vo>Y�q>�t�<����?���d�L�/��H����C	���%pX��]��O��m��q+(���?h���);�8?@�򽞍~>�/?��E�U�e=�ޙ>f��=��U>ͬ�>}��>-��=���>��R>���=���;Ft��|��p�4�`�����>�qb?$�aC�$���#��N!�3%>��>����l���z�/��)��>1�����7#���>)G�>�?&�U�����b�Bz�Q�<�W��Գ>�c�=Lc>u:��YD��Lw>��?�����>o�?T�;?+E�?w�1?=r�=���=���>�>r�\>�&����z=SB�>��)?�6}?r
[?A�>|��=N�h�#�B>	s(=g���8=  ��X���4ݽ��=�y=��[>�.>�� >y2Ҽ�6�=��1>uw> !J>���>��[?�Ÿ>��F>U�\�5��n����8��>5��=�@h>y\�>C�(?��>5ה>2���!�]�j�� ؾ�.�>̗8>P�y�Mnw��$�<+W�>��>QE?�(?��#���˗�\�>u?>[C?�B0?��>���`�c���jӿ$��!��.���=�*؋;\r<��gM�����&�-��D��D��<�d\>)
�>�rp>��D>�>TD3>
=�>�G>���=�9�=��;E;�G��M=�����E<�&Q�����=<ż`�����NI��?�pw���ּR2?��?D�C���5��^^�+��������>xr�>̕�>���>�a�=n�w;S�X�C�.sE��;�>�dk?@��>�1�V��=��6�ح�����>���>­>�N�����9P��l<C��>c�?^.�>�@�)�V��dg�����c�>�롽��0����?�u\?m�;���$��� ��k�aJ���A>b�>u�ŽF�q9ܾi�[��
�d��a��g�>a��>���?�A�C�=W]��O2���{��3��߽�*�>�F?�ݩ>\�s�þ��
��v4�h��8�B;�X>Im�>e5�>��?�O?��k?��?�>_���8�?$��>�s>A��>)��>5�?'�?���>>�>54�=�ߕ�0$���Y��ݠ_���"�ڬ`���$>Z�!>�F���Y�=�>�ͩ<�4@����;&_�=,`>���=�`>ڏ=ی�=('?�WK?<����>N#�>/�b�K��o���g�>VI�C���2��3�>�&?Sv?�/?�=O�X�,�F�ࢣ�W�����>�'1?=��>�/.<��>�d���H���f>�J$�(���8���r+̼<S�>��>I�([y>EO�?�YP?�%?���"�7��t?�+�B>Gz;��{?g>�>��`=t�Ǿ��O�jMY���N�lhw�H�=
�ؽ:��=TKd�V=�c4�>ul>���=�w�=Vu+>����G�=hN=!_�>���>�	�>>�M>���=F�3�6�� P?9a�SD߾�N��ڤ�ذ5;��I>�yB>>1�t#?��ݼ��c����.�J����>���?)��?��e?�\�>'���U>K�g>�\>�Ơ:u^�#�ɼ�~��3��=ݻ�= �����u��<�6�>x�$>��������پ��Q�D�ٿ�b��(��i�g,��E�g;Q>���׽�����,|>�A=VY�@�����2����D���W�=;��?&x?7�>�l>I��C��<�����6Zھx
`>��뽿����.��ݾU;��:5��	��p��p�P>{$V��r��{R��;r+��4��w�>�=&?N@�4��m5���=5>��W��T��䍿�*��wu$���W?�g5?�پ�i������d�=T	?x!�>�qf>�g��{%�8b�>�X?��8?�==�󂿂{���)=YȮ?>E�? 1?�S���}����u������>3[D?'��>Ө�ݙ��FU�=5r��q�??���>W%�l=b�����1�=�q?�pD���E>�
?d�?)m��i;"o8�����6�']�>#���vѽ�y���k��!��,��=��>�N.�y��/��>�A�S�N�l�H����6��yW�<؆?��d6>�i>�@>	�(�����ω��)���L?�?*�S?�k8?�^��S��䮧�M��=���>1Ӭ>Ƭ�=���y�>h��>yf辙xr�6�E�?�J�?w��?!\Z?��m��<俬���
R���ؚ�K�=��ڬ>��<�քa��h%>��x�.�=�u�>��>��y>��i>#/�>�Dp>M�s=v/������Ֆ�T����}A�'�,���<���Nb��_�
���	��O���C�<Lqν����K�rg9����ޯ�ə>����>���>j>b��>K��>]��Ɛ��̀��� �%.���3��L�l�ܾ��þ��A<Y���� ��.̽Z� ���7?�q<tu'>J�?G�X���s>���>���.>�>��>���G�>���=�m4>���>xs�>�j�=�(≠*>(�����W_���&>�?8�$�n�����;��l ����M�X�f*�>2��=9D�
���`����>����G�۾�`���P<ғ�>�?E��=T��gB�<����þڌ�=�V< i������a�����S>m��>B�?Ʊ���c>aW�>��K?�>�?�Y%?��'>p��>5B�>NG�>�,�>��`>	�>8?YU6?q�m?�<Z?�?�#�<�u�]�<>�Z�=��k�Խ��	�5��c��N��QsR>���>x�<�7I>�>>=܋=b��<d5����佗c?>5?=�/?�^�>I��>DƔ�J��X����=C��>�>G��>�j>��>�?���>"��>Uo�=�;��M��([�>�+�>�J�t�|��~#�ßj�%<�>`{?=�d?P��=�NƾL���,ۇ=/g#>X?�P?C/?Q�>t������lӿ]$��!��킽,O���;��<�b�M����7;�-�����N��<��\>��>ԃp>.E>�>�;3>�R�>$HG>wӄ=��=�:�;ޚ;%�E�@�M=��#4G<i�P�����|Ƽ������� �I�-�>�7��7ټ��?�?�z��n�ٽ�.���Ͼ�A��YT?�D?l��>�o�>��6>�C�!-E��z�����|?W�w?��?���u�=撝��oF�u#?�>d=��Ľ��
�U6�$\=�
?|	?8=>��0���L�`i��̲�P��>1��=}�� K�?��n?�l�&�4<2�8�ʊU��������>q��>�d`��<j��&ܾ�m��>�yƿ��k>�>Q�>"6�?�������<�#��Ϭ�����_ھ��U<Ĝ�=���>~��>�w澜$%�aG.�*�X��-���"�=��>"�=���>�c?��?�d?�?\]?_��R?�]�=C:�>���> �?��?��?���>��>�-�=������w��<�s���=��>j�>�l�<��?=q�A=)Y=�4��@$�˨�<�O �a��<:�K=��=��>�?�?쿳�!�)>������ ���U=?�=q`>��=�퇾D��l��>�?V�!?/?Zs�=��׾����h��DS�@�?%t?]O�>9}�>Y��>�X%�7T�X�>G��>1Z��V���0��Pq����5�^�$?�K�>o��=�a�>���?�?�7�>��=-#:��������W$�>�Ӿ���>�y?��پY�X�7�C���e��r�h�����>��n���=Ξ�#���<>4�;�U�<>Z)B>1�Z�d;����W(ڽ#ށ>��>h�,?.��>�������H7�M�L?�ׅ�H��F����Ծ�.Ҽc_@>d�>�n)���?�$�тs�垿��0���>��?���?Ηd?b�"�-�彴�N>4o->M#�=}6�=z�彰]��Z��_>`}X������$�f���Y>�3@>ֽ̖󀳾g�n��߿ֿ#���~�=��+}���&�g*���#wվ�g\��Ǿ� M<JI�a�>�AQ=���G�����7���6�e�?.Gl?�>^��GM"�{��WNѾ7F�>N���S�۶���A����ٛ���s�ѣ�f���Q���M��>�>�.V������-'��N��!�R>j�0?��ξ	���܉���<� >p�;D��ɞ��yʛ�~�0Q?��6?ė�;��BϽ5f�=�?���>y�'>i9���νq��>��-?CO/?��y�ف��o����EL�?��?�^0?�3�o�P��� ����>7�)?re?�˸�����S�}�u�>ia?�0�>�1���~�~?8�$��>��,?��/L=>@�?y�>d�v��7Cٽ�,Ӿ���;LQ�>��N�����;�����zE�=�]�>���>y������T��>�v���N���H�����a����<�?Sl�u�>v�h>��>޾(����������,���L?�?v�S?kp8?]���i�
��>��=�i�>���>ͧ�=����N�>���>�Y辮�r���ݗ?�7�?���?�7Z?Him��$׿6���'�˾���U?=�>���>7���^7޽y�d����=���=�}5>r�>c�>���>l�}>0>�>UX���~#���PŊ���B�eI�G��j���{;�C���=��?傾XQ�=	��A81��~��%������|��%r<Q�?cx?�*�>U�a>��>2엽�[���	Ѿ@��]����
�6�;��}��,�^��x��h�Ca ����ן?)���I>��5?���=�}>��>��y>ʒ>��i>i�r��NV>x�=L\B>�3�>iQ+>��R>?�o>�Z#>M���<e���\8��3þ���I*Q?\���u��f$K�Q<���@)�u)>?,C��MR������ ��iM?�:�����MM�v}>[��>��>�	?>�\���=��ƾ�I@��Y�<0os>���>�[�=����8j@�u (��?��#�_EP>l�j>S�$?��?�$?ZE>�l�>���>@d�>;�>��>W_E>��>�a?{,J?�j?��Y?�Z=�[��7q�>�8>������=��-�����_r&��{�>8�,>��q�i��^��=���<n4�m�c�ٔq�K�#>"�?ķF?�"�>���>'�2�A^G�L�X��!�I;�>>�p�\#�>H�>W�&>�Y�>�S�>�@>��|��j��p����>�P�>4��P������=�t�<^~���i?��W?��5�n�ݦ[=5�>��=�� ?�._?e@�>��=�mý�(���߿���S���4|���=a�,>z���}þ������ӽ�v��m�<N9>�(�>���>L��>���>�;l>���>�;>n�>�� >�'=�t���� �9=��>R�~<����Oq��lռ������	�l!��4�,��#�=˘�=��?f�?�8�#��.ᴽ��̾h�����>��?�F�>��>��>�ھ|uW��#���<�?�O?�b�>ԯ�@"�=T㬽�)�V��>9H�>-tr>-½��S��EǾ�f�=ڇ�>g�?6��>#(@���K��_�$f�����>�����?����?!f?*�h��"e���H��P����v�>�]>� ���х�����iT����r4'�F*��:�>)�>Z;�?�!���.�=�������D~��a�����=��]<D�?Θ�>ʺ2�����Y�)�|�߾-򴾹����J.�!N>q��>:)?�2?P�K?տ&?�d2?��p�L{�>��>�;?x��>���>���>��>��>œ�>�M*>g�9=����񁾕�)<2~'=~��;���=@��=�5���GY=G�.>X&�=v��=@��=�hm=`z�<g[,=Ԙ=�œ=@D�=� ?��.?�!�K���J��Tþ�����k=ۜ�>au������g��W�>���>=?)?���>�F�5��2@ ����q4�%#?�Ge?f�?��/>�B�>����
��v%����z>��=R���h�7�L��������>�9�>;�0>��>�A�?� ?q�?�"���Z�k�����=���>.�?�I5>��=�G=�&���*�^sJ���m� V+�����l
�~��=�ӽ���"�>9�>H�=>��<��=�EPi�/w�,@�>�J?��?���=�ڷ=
���~��KJ?�����:�1Ġ�8m;r;"�:7>�H>ٽ��?�	���z�'��'�<�A��>���?��?WDd?a�G�;� ���[>��K>�>m�<O�4���H�w�/�5>6��=�p�X��}�P<|Y>�%o>+��ǾF�־>�1�/D�� �C���8<����$������x�o���O�nɽ�<��X�#���l�2����(w����Pڣ�p��Jj����?!�?�r'>\̑�ݙ6�?f�h��-+>�܈�Iu˽�`۾�~)���̾����o�þ�j&�lU�N�^�+�>�E�>�+�S/��bU��uE���ܑ�k��=�YO?2��2���R��
=*.�����`������ߘ��ɼ���+? �?/�ܾrAξ�7!�8�i>��?�>0'>8kԽk(a���s>��?�,g?��R�>�������>v�?}�?j�/?��O�s��)^��*���>MB!?�@@?e��񏬾�7��o� ��jc?vj�>"y�L��p/��66=K+?	�a�i�m>�b?B2�>p���&վEu>�|p��oj���8>�>#w<��
=��>�>>���>�z�>AȾ��
���9�>�e���N�h�H����N����<N�?��/�>m[i>�0>�)�'�������	� ��M?���?�NS?�q8?����*��cb��b��=��>�>kw�=��	�rÞ>u��>��義br��{�CK?1E�?���?��Z?��l�Q�׿PȞ� PϾ�뾄����=N�->� �C��=(H`>ȝ�SI�������>2�>��>�%V>(��=, �<�Ç�R�#��U���훿9`���a��=u��� �G�B����CþH"羺gν�:Ƽ�X>d�i���n��N���넾�?�<�)?�(?�	�>)g>X�V>����'��2����fD����@엾�����W������Ǿu̷�W����t9�¡�>(�=m��=�8"?�B�� �;��>��ý�F�>���>/�&<a�>�'�=�z{=�	�>��>B��>Փ,>�JL>����ʥ��k��G�_��[�Y?����}�x��@�_�s�c�>A�>A��X�;��r�������>�v;=��`������<?��>�ll>9���ا=�h�<�Ɇ���[���=$Q=´ <r��>��M�,��Z�?�
�׀�>��>*�d?蟏?��]?��F>b^�>��?j�4?/p?ґ�>��=^@�>#64?N�P?�p?�7?[> �w��cK>qj.=�,�wK�9t��ҷٽ� �<�LC>��=�� <xx�;b�">�L
= s�U[�#y%��}��4?��H?
�>��G>�]���9��F7��h�J�>�Ƌ>��>Ͳ|>�#�>)M-?�?zl�=r�������ӎ�>A�>��y������`�=�>r�F?ݟV?��H>�iP��	�=�@���-3>,�?�	V?�?;G>��;=����ǿB�R�MF:�Rڲ�m�4�*����
�⾫���m��������x�=vҽ�>��J>���=�#=׎�>�iz>PB>��+>���=��G��|���!y�<�ҽ36�P�Q��o��T�=���:0ý�Q�lq=�a�<�1�=�.?\|)?�S����A��� 岾&^�+*4?)�?�q�>�[�>G��>kƾF���|���0>�"?]˄?�w2?�����s=�N��-=6  ?�!�>$/�=�O=I�Y����� ��]*?�aL?@�=􆾲s�?t�[߾T 	?�:�<����Iٗ?���?A�A�r[#��D'�f�|��ܾ��ٽ�X�=̉���S{��v���5(�4$��1����>�>���>^o�?�b>��N��Ll���9����Ŋ�\��==n�=�S?Y��>��޽:�e��@��L�澰��=��=ۃ�>��>�~:?6_5?��l?��E?�8?O�&��Ո>N�>|9!?Ff
?2=�>��?��?+�>���>V6�>%(>�˽�}�����dV�ǉ�=,M�=���=�]R����=_&?<�屮��<B[A�ש�;��G<Ӕ7=��>8j>:S>_n?��C?wk�בӽ}ʽ�����q��H2;���>��=5p�Ċ��_O�>�G?�&?�͒>��N/��?v���N�TLA?�g�?���>
�>� ?�Q��I�#t�����>t�%�A�����u�N$���>��#>>�=���>�m�?��?��>�n��<i�����~�N�d|�>���m>�O�>�J =',��O��kx���\�*�	����^���d>��l�N�\�>��>��>��=ݗ
>U�=۞������O�>&?�IB?���> �l�,L���V��O?��g��>��M��KfӾ�J���7(>�;�>89ļ��?��ʽ�h��W��ִ>��g�>�"�?e�?�(h?�m#�c��;�d>;
�=�!X=�(�=�P�/����x<Ёt>�H=��n��LS��Z=���=v&;>�kF�`���Ћ�9��=Pk����C�p-�t���Y��J��y�<y����Gz	�[B��V肾`���jGT�Vw��rՙ�M����ٲ�~~���?��?�5<�' ��d\� �I�mH���: ?su������h)�+Ā���J%��J��)���{Y�1h��b�I���>^SX�|���Z}�^)�(����9>>9�.?�_ƾ���>����J=�`%>�l�<^���ߋ��{�����K�U?��8?����H��?�ݽ�{>z?i)�>�0$> U��J�'D�>#�3?<�.?{��k4��.���]�|��?d/�?�rC?l,���_?����3
���>o�?
�?[�K��j�Mg��(?�R?���>	��X������v?b_?tN\�,�,>��?���>-K��T��lS=�3���=���F�>��<[�a�=[����G��=���>W�w>��������=̓X�?Q⾆X>���������6[R;Ϭ>��R��F�=�P�=�����7��S��x8���4˽UlN?��?�K-?{�7?�<��+"�*�T����>���>�I�>�F�>9�1�k>:�>]D���!��+G����#?ׂ�?X��?�Z?k�P�#���q�卾�$o�N��=�F>�b_>�r���=7t$>�S�=�o<T�O>>4�>E\�>i�r>�v">�%>���=4���LZ$�J1��X挿��B��P��
 �u�w����<�s�,s*�A[�������f���~���ļ��e�R�D�^�����ǥ����>�U�>�~�>��>��=V"}��㾱j��/υ�8�)����T�(��nX�~� ���߽J�ؾX�����B{�11�>���=��=2ֻ>�À�)ѯ=��>���=���>7�>o6S>��= q=F?= g��g�������>.�����	����Y���WG��?F�??����Ӡ�#�V����u��=Q��>���>�Q>��k����C���>N��=�Q�����9���ra���z>k�=BÍ���=�I��B�T �?��>ʡ@>��=�A2��L��HF�;a$?�'l��8�5��=R$?���?2�?��=��>��t>Ű�>WLN>��y>�d�=���>J��>�J?|,R?>��>��n=J鉾7�=n>�>�b��<�����������v���@�=w8�=/��=�v�<�N;�(S������6=ݗ?=G?>��>Ѯ>l���,�j"V��}=��t>jN潭*�>�I�>�O�>Z'>H�\>MG�<z���K␾j���>!��>%<~�,���W�<͈>�_�=z��?$U?p�k��z=��,>=��<	�=d�?_�>?:4�>3��>HYH�j/���ٿ�$��J�򾖽�T���?=�%�lrw����<p,��pϽ���=���>~�>��[>��>-�&>7>�>)�>*R<��<=�?��JnǼ�I=�^�=f#��k�;])ȽO6���<=\��s=������mep�u�q�Ě&?ǋD?��&���T�-������\�߾^�?f�?��>��?^f�>��о^Vr�&�'���z�G��>%t{?�Q�>��̽��=I@�a<	��"�>=	?dn>M����-���;�O&�;��>� ?'��>�n<):H�K��'շ�� �>�0;��,��I�?C>?���]�̾g~�0�%��5�,��=bAν�����&�gh�yVB��t� �&�����7����>�:�?[�������f끿]������v�p=���;˜?>SO�>�T�Sh#���U���	�?�r�u3�>�s^?���=��>��-?� =?�Fq?��>?���>6��� ?���?�<�>��>_�>u��>�rQ=-%>�">~:O�O>�����7�=�ob�f�=���=ò:>$��=0 �q�>���=}쌾�p>FvR>W��=y�<�_ؽe�:=f�K=��?$�>
.�����<�|=@���)=~V=(>�4u��W���ZֽR=��?-�7?}G?9�3>����/��>%���>
�?Qk<?O�?ng1>*h���������kI>��=��w�bg�c������d^�=�g}=iϼ�Iy>tx^?P0?�<?_��=T���{���!��+�>����qr�>ny$?0�>�>��RS���|�_A��/�4�?�[�����G>P��>jk�<ɴ>-0�>�e�?n�]�μ���=�O���>@�>A��>��?=�:.>�|�����v>V?b&�5�<�.L��	������g�>d����B=s:?�������:���:y��%d?���?_�?.�A?=��vV�<n/���8�=�=>�[�wԾ�Il �¢&<0w�>����:�1n�6��=���>���>���=������+ν�ǿ�c��T��/���F ��Bþ��;�d�<iӦ��cp=p��x?�(��=WP�=F������5gھ<��OL�?'�?b�=���)�E�̛�8)��L��`pýj���p�'�s�Q�sm;���������p ��̾z|�>��F�50���
|��1���s�n�C>�&?P�Ͼ`~��%����I=(F8>�|=7D�D~��ri��*R#��S?J�3?�WھFeᾅ&ٽ,.H>�I?�0�>y=>q��������>�f,?�"?�����H���/��aڹ��ǽ?���?VH?�̠��D��'��n�z�+?  �>B%�>&���, ��=��?D�)?�+�>�+龐���L徽?��>?5_���r>�C�>(��>�F��������8)ؾ�=��ӽ�쇽�鱽�Q�������Y����>å�=SӞ�So��YI�>«��!�H�_\�(�=���	��D>�`�>3�0�ǃ/>f��;����;f5�xꗿ����@��gD?�أ?<?G�e?�v��m��x�&6y>6�>��1?
T>S�>�T:�>��?�5����������@?���?w��?�Շ?7�k�X�׿�&���W�������ǫ=�q>%��>��'�>O1>K�3�z�m� �>�x	?D��>�T�>�D>\�=�ɕ=#�����"��q��pW��V�)�&��V�{�ܪ�� �i;���Z�Ҿ��Ǿ�2н��l��2������|�v�^=����O��=Uò>f��>�-�>��>��>���4��V��C��=���j��ˢ���/��w%�D����������(���`��t�>�X->G��=�
?h�ܽ�T=��>�s;��XX���>���>���=_)�=?Ϊ=|�>�!>�w�=אm>���=����|�v�1��3���=�=?�����ᅾ���-�&绾/׃>��	?��U>�G$�����H��F��>3Oq�G�X������	��ѡ�>��>�{�=|�<	�\��D�`��@�=��q>���=��L�镈�,&���_=��?<�;�Y[>��?z}?��?`�μ�԰>�Z>7�>|c>��)>�a >ý>�q�>��i?�8a?�>NW�<���r�=��>2[2�%S(�������uT�S���6�ιI���\�=D� =��=�Ҵ=���S$ӽ�<?�7?��>:��>>���'l,���g�+6�>�+k>�Η��Ȩ>�z
?9��>�LQ>:o^>������`��ZI�$��>���>��s�0��X^f��$i>�N+>��`?�/O?�99>P��L�> �=1��=}}?�T3?�h�>*��>�-�=S��E��CG$�c+�ii����>�-|>}�ki>T�{>�ͳ��o�d��>O?v�?O��>
��=I��<<!�=1��>��/>�G�=��*>��=Nʽ7���1g�=�����ܽ��=)X%=��>�;��䓽�����|L�]������5�?@�2?�!��A�+ҩ���������5�>
?~u�>l�?_�>0ӧ���B���*�g�p����>�e?���>��"��>�=a�%�8�>ͥ�>�z>��t��[=�ѡ��}:=�Y&>��?��	?>	�m)�%A�r�.�>sLܼ�Y���C�?��"?b��Uީ���V�<�2(�.̤�D��j�fG��.*�+�F��
��#�������=
�?f�?j13�jゾ�쯾3מ�\�����U��}q��f�<��8>�f>>������a�������� �i>f?%k�=��E>�KW?��n?��?r$?���>S��1��>Y�,��ne>���>�,?��3?»�>p�>��|>�<�=�b��	�ҽ�~d��1=r����q�=PQ>�}o=�P�=�5�==��<Z��=�>���=��=��F��)��~�)=H��<%?>�?������ҏ�<!����=�=���=��b<���z����.�=���>%�-?nw�>�?�=�fƾ!��
���=͡?�� ??h?Rb>��=Nܾ�d����(<�U�>*�2�/0���ؾ�*ȾQ3f�C>���=E�/=���>Ձj?K�B?
4�>�3i�W(�X���1�1R>R��g>Q25?]�>�e����c����sᄿ�K?����>�f)�o#��F@>���>�)>>�,���OX>��:��2k��C�7<������8� >���>{�>	��=���=h���2��'�Q?K��kg�o�c'���>��v?G�z=�9���C=?G����榿��Ŀ�8쾕�.?S��?��?G�j?�Ki��"D�%%q>o��>mvi>�W=j;��0$����^�J>X��=�;'��#D�%�����?�>�>�����O����e�����L������=��LŠ��Qľ�^����5�����-��R׾��B�,�-�Ȱ�(�ѽ�;��k���'��ڜ�s��?�r�?�E>jjν�CS���;��O�_�;�0۾Pr@�xW�"�3���W����^\��:%���A�G�,��Ě�S��>�M�v����E|��&�������(>�'0?r_ž蹸�N���=/�%>��	<??󾤙������ga
��7W?99?�⾗��������>&�?o�>Y0>b��g�Ὓ��>t�4?)�+?�/м����
���D���х�?|��?X�??��8��>��
��'��?�-?���>��|�Cgƾ�ݽ�?g;9?�]�>\G�}�������@�>��[?2yJ�L�^>���>Z"�>��kk��B�ļ5y��:v[���@>3?�/)�<V`���2�$��=�ɞ>�y>�.Y�W������>�Go��W����|��� ?�ہ>{&?<�N�Խ�7�>�Z>l��S@��5暿�_}��?6y�?�f?��?��¾#���̵f=3�f>�Lѽt9鼕sM>3H0����>p�?�/Ӿu)����ᾕv�>�?9��?X�3?�$��+ҿ�ޢ�*Q����>�c~�>���>F�>b��Q�;>p���9��2|c=�
�=�>���>�p�>o��>UXP>�?�<Kt���i$����� ���r;�|m�����Bľ-���{���)�-�0Uоk����K����=����T�`��	��֔�=��>�3�>�5�>h�i>�S>[J��7���(������|#���� 
ξ�E������2��M���﯀�@�ս�
��d�>�>E�(>�?�j^=g�>ϱ�>F�<^�6��S�=��l>5Ȯ>۔�>�2�>vcW>.�n>ka<��~>TF�=e���V���@9��XM�1�;W�C?�rW�������3���ܾ�&���Ą>�/?iN>�i'��z��w��0�>�MI�4�e���ν������>���>�߸=��B@��}����vY�=�v�>>�+@�ة�������=z]�>A��	W:>+��>�D?%��?*�!?�ݳ>��>��]>>�����>{#�>n��>��&?o@C?O�$?��1>�4>yѲ����=���=$�L�׽�߽~������<���>p{���=*�5>m�=FdY>�s>�>���&1�UȼJ?��7?�"�>��>jYU���4�S�<��Ϣ���j>�i]>�[?}��>G��>M��>{y}>�{��y�.�+��*t��q�>�ܴ>|�g�����O��⁀>R�j>�*n?�N)?��@����x>�J=>�}�>>���>( �>&�/>��= ����ȿU�`����Q��i�&>�1]>/�-�CT��e����CG��Z*Y���.?��7?|,?���>ұ�>�}ݻL�>�6a>㖏��B�=��������_߽�L��J@w��8���n=�s�"�Y>�?&�~+��YM�=
�A�I�ռ
�<^�?��#?b���l��Q5���)�����_a?�bQ>���>�F?�7>T�!��VV���^��4�����>��H??�_��!u1=��>�:��>�?o?�<J�^�^��=W��d3A����>[1?=*�>�6=F�J��S�����*>J��<}���A�?GdB?X,���ھ'�k$�� ��ڧb>��"�F��N���<����S���;7�j��g�/��`�>�߬?�f���ް����@n���-��	�<��j>
�z>?���>NY�}���:���7�.FȾ,��%�!?G�>��>"$? nO?2�f?�&?�G�>T�-�*o�>l��>U� ?�*�>']�>��?;N�>KBo>=-n>��0�%��7����@w�^����=�a�=)�/>��>�T��ł�=�U>-��=t�����	�1S >l4�<_��=
�=�$->D��=��?��?9 �=#�=_e���&���w;�c�=�O>��(<g{�l�=��t>�0�>�a?Η�>q�\�	[�t��G�����Ͻ�?h`W?�`?�Q >�_C>^g �?${���>��a>�@�������m��yǾ�ɒ���>Ih�>�d>Xա>�0�?po?���>^]��Tr�:=���w�ɧ=���>��>��>��I>�����ﾇ�U���e��Qx� ��hz�ρ�� Q�([>w�F>�P�=e=�=Δ=}�E�k�,�4ڻ���=���>���>���>�>�$>��S�R�gF?�0��]�#���E7>��=4�> ?"�>F0?���>A�v�����ud"���?���?��?u�?B��Xν��>J(�=�G+>�:>!C3�l�i=��>Ì��Cy��O�<v��z��dx>9a�>��ֽ�m���uվ+2G�6��(�G��񽎰����f$��0���с���<ľsbr��ӾFs��p���5g0��׽t@���ʊ��د��iо�҅?6ň?�q�>�v�0� �,����⾆�>�\��`�;=��n�%r�<�پ��7��F%��>��Z�YIS�7���$�>�w?�O���I��\K]��[̽���>�?W����\�%z��'N$>��>�����0�����☿��˽͖�?�9N?�g��!�P���̾Ȣ!>z�F?�M@?�d�>�ož�k��w�>'�>-;C?Q>�'��|Rg����=hw�?C�?��[?|ؑ>��F�2o>�y��=}'.?=?ǎ�>��'>jžH����:?�u?E�}>���������rt>���?'�X��ql=r1�>���>w =�����=3N���ߎ�o��=6uҼ�y��`�����p2>V�>ꆃ>-�f�4W�3!l>K�˦\�=V��>�>㸾�m\>>��>4�d>aG�=n��<�A7�A>��K@z��A�<jl?���?.�#?���>`�.�K�/x��%#=��D>�#�>�>ż�i^�6�p>��a>66��Q��)�'���>��?-��?�g?޽@�sۧ�5������
����U^=l�=k��>ބ��>+�=�,�=��=c���M>d��>Q|>nO�>�rk>��B>`��=����������0����x���7��'ྡC:��z�0�p��&���پ�;��ؙ���Z�AGʻ�4�#��;�k,�M'���!=)��>���>���>u��=�!R>�[L���f���9n�^���׾��־��̾�(���0�����5��6��z��Ȃ�>��E=�0>��>z��C��<�ْ>)+���Q�='&�>վ>���=��=��D>�Ժ=��>�	�=������ �=oq��D`�n&����I�=��i?�W������ �����%�6̛>�j�>��V>K �_㎿�+��br>k2ͽ�uB�Ui�=�{�>N�>��'>���=��н�'4<�D�	!>>V��=�@����5#��ebl��f�\�*?pp��&ƽ�V�=	�#?M�?p+?{�=���>��>�S�>�^�>�=|>��>�p�>���>��3?5/L?m�>'!�=����=k�o>�,�e����=f��j�B�a����Bн]�<7WI<�����=hq�<��`=�x��!�� ?x�>?Ȩ>���>{O���3�_`���/<��F>���<4Dg>[�>�<?�1>���>8ɢ=K��h����S��̠?��>�pq��Z����=��=p�==ڌ\?2V?V]`>p��(k�=Bqh���4>�{?U�B?��>�p�>2�������iӿ�$�?�!��ւ��\��"�;��<� 'N��w�%g-������:�<�r\>'�>�p> E>�b>��2>�c�>�"G>��=1��=uS�;�;#�F��GL=�[�`�H<HnQ�M�����ļ͗��ϋ�C�I�l�?�B��7׼�1?ґH?/"	��I�� q׽өҾRj��v�>���>$�+?���>az>�����T��a ���r�JD�>��q?�
?e|���L6>�c���� 
�>$n�>��>�n��A}�\�+���/>���>�k?<�?���/�
$��ɾ�b�>)������ Յ?_�D?<��Bs��#'�y1,�%�B�
����z�/y򽋐J���#�
H�j�����n��n��=}U?dV�?Q���nF�r*���� H�����<W�>R/��A�>��>a7���C�����g辘������>nn?�P�=b��=�`?��c?���?3?Ψ�>(�����2?c(�%]?���>�
-?sn[?��>���=`,�=H\�G����z����x����=�ʽ�h뼪�g>�`L>)�=S�=�	6>�(z=S콠� >�fK>�qx����<���Cq�<|���?�c?�M��=�Y=e�-��.<��o:�.>O1���K�w�=��^>���>��"?���>��=Ƴ���оX[��\�<�0+?�F?�A?� B��A�<�� �
�J�]ֽ��=DKӽa�v�8 ���]��S�Ľ08=>�r>d�>��n=Ëv?��?C��>䡶�����������!�i=8'��T<o ?��>VV��^h�0J��%#����+����>��G��N8b>^'�>;<�6�=.#�>�tR��0�8�>���Qҩ�n��>-x.>�I�>�>��>N��,��F�?��%��cg��c�~�I��M��F?Q�Ƚ��ѽWh�>�w��b˚��(��zj��;�Z?<~�?]ֻ?+zQ?Ǉ��1��>Х�>q>0�=m�_�:�=����=A�=���=/w&��䞾lv����>{�>"��%���,�Rև�Wv��R�\��� �����]����}��V�P׋�4�ƾ����	������櫾(L �e๼���������d��?��b?	�C>V�Q=�+�pC����U���NҴ�����h��z ���}���־���[��2�J�Q�����[i�>��O�����bj|�J�&����;/>��/?CpȾ����>[��ex=c�%>���<�������ɚ���'�V?�9?��侞������>�Z?gL�>A�'>?�1�윎> �4?.?��Ӽ%�����N�̼@~�?-f�?�tE?�|*�6�@�������	?jl?H��>�(����ž�Ƚ59?�[6?f�>����̉��O��y��>�V?1�]�ָ>>���>���>|�Խ=畾���˜����[��=¼�u#��5d���<�2��=��>�Cn>��x�밾��>��˾��R�QmZ�Rh��Y�G��>K3�>��9�0��=;d�>�N�τA����eE�xf?C��?~�>��W?d�󾓱]�sp���>���>BT�>���>���7n}>~jA?�+��&Ր�S���?4��?L��?�"�?۵���a̿����+qM�|	����=<=��>�Y�;�G>Z5�=M���U{=�Њ>��?>r�>�>�>���=)�=v{�kR���� �����A�p.�����a��n�⾳�^�է3�38Ⱦ�Y��/罏���M�h:Q�]��K�lz<O5��SV=C��>���>*G?�q>c'C>��="$�xg����y�<� ��{>��x"���ͽ9GK���n�I��8��	�9�>��=a>��?$�x���<�
�>o�k��&�=^�a>0��>��>�>�`�=��=�n=���=5{>���=k���ꀿ(:�Q��E�;��C?*�]�y���as3���߾�ϩ��g�>�}?~�S>�B'�$���� y��f�>��G�J]b��̽|v����>Ն�>�ռ= r׻+1�a
w����	ߺ=���>5e>��x��@��������=n>�>C�̾��=�1v>&�4?<$�?2�,?��=Q��>��>�c�>m��=i�}>e^�>��>��?]�)?}/?�m�>�H�=�������<���=��.��Oi�W�׽�jf��������<��6>�(>#�C=�HW=�Q=�r�j���W��=� ?w�=?<��>�*�>3�q���%���R��'<��n>��=
_2>��>��?��>o�>�;s���B'��9yO�WJ�>��>ĕm�2:��X����>�#�=g�f?��~?���>���=(��>���=7O�>�j?�%?���>2�>��<"/���ۿ��!v�;綽Ƙ����=�t� �ռ2�=������Lن=i`�>�c�>�]�>'e(>Ⱥ�=��>B��>��9>�=��~=㹼����<��V;P��=��A�g��=�"4�Gx�cZ~��#������ ���A�)��F�)u?cO$?(�����+�iSH�z�;�Ħ���>���>�Q?�E�>�p�=��#�8��	���+����>>?]?��>�L�D�=�Y���3Ž�`�>�m�>C;%>*%�C���՝���V=0�->v!?教>��2�Jbb��]�X� �C>SԽ��׽��?��F?.��"̙���o�7"������m�/^<��WZ�_50���<���@8�L�Ѿ�O>!p?���?�'��0�k�;
ھ&ӊ��}����S�=����X�>C9/>�)��#Ѿ��:��t��BX�PՂ=/W?3�?>�!�>�s?~F�>̢X?�E?���>�S�m�?n!>���>���>%P?WS<?�|�>��U=bm>rMT=���h�����t=ѳ�=�3i>{Վ>�=>�`�����V�^���>/J=��<�=�>k�<�A%��;��*>�U`=)?�'?�����Ҵ�7�5�i����䩺���=�0�> *˽��R����=3�>���>մ?룵>�0|�p������/c��р�<�C&?�s7?i2�>
�x=���=����U��t=���=+�N�f��{���	|��F,���>�s>�J�U�O>�a?�5?ġ�>Am�<aL������ʾCv��%����!��>8}�>,�侁y2�N�k��bs��+V����>\Q����c�X>�Ƙ>l��;2~���:�>Z!�;A�c5>�N��e��Ð>�Ϻ>��>'_^=Ux�=㪗�1(��]qK?�3��w�u��oڽ���_'<��s�>��>CNZ�X� ?޷T>ځ�%���q*�;G�>���?��?�4�? TȾq�@�ߐw>RS�>H��>��=T��[�Q�z�(<���>��_<����Y��3��秆>bɪ>ڲ��o��r���mǿYRc��٨��jS���y���1N����Ⱦc]1���g�ؾ�K����F��[e��Vݼ�Y��ۧ��4þx���3W�?6��?�/x>s���ʲy��$�6���vt�����uͽ�(�����}�"���!�r\<�w]�3}>���/���7��a�>oY����ƽ|�)�6$���K?> �.?�bƾ_������e=̣%>A�<��:�������,=�@lW?c�9?�뾓���V���>٥??��>	�&>TX��h�%�>��3?w-?��N���+��̝��#_�?���?Z�O?rUq=3;�sG1�k� ��8#?��>�N�>u�`=�h�]�>z�D?X�R?�� ?�k¾}�m���� ��>PSi?VEN���=KS�>��>�o	����j̽��-��r*=3����� ��/�&y���쮾���:N�>��=�����2�����>�������5D��4?�oH��e_R����>����>l�>GD<��"��K���Hy��s��B?���?�Z?d?<d!�=�7�gl�`�!��.J>u�?�>4>m�>y�?�g�>\i��$�h��Ğ��D?���?��?�r)?ؤG��=տ����Hk�������9R>��7=��H>{�Ѧ�=>&>E:�=%ǻ�`y=�0�>�>{Q>{z>��>N�/>���������蕿1�@��=����X|���*��Z<�T!�pq���=���G*��̽]%Ľ�
�=n���[V�%AǾ=� >Ȣ#?E6�>ud>'N�>0�>%�`5�5=l�ʟ"�
F����q?�e��>`ԾA���Wܾ���ZԞ=EA���0?yI$�	��=��>�K2>��>���=�n>��==@��=旀>6��=�_=��>,M=Ő>�G�>m9�>J�=�����Z��)�/����O�&�2�Z?>�"�[㞾�"�ٺ;K���傅>�y?�a>["-�񖔿�ʁ����>��W�=XH�g���;Ki�>��>�<�=V����<������v��=���>d�.>�=�ǁ�^��F;&j�>>߾έg>w6%>�zH?f͈?�9?�<=Q`> ӌ>��+>�S>�͛>+6�>�>gk�>}�#?�E?��>墥=B��m�*>���<_������0�þ�ي�ҟ;�v��T0��:I�3��<�S���='�ʳU>>�>��>}�!>���>E=?��x>Hd�>��M�G:�qt��� =u�#>�Ӿ�'�>�B�>}ɺ>,{�>�>�>Ѓ�� U�{a�롮>��P>*8�w$��M�${�>��;>�4u?�#?�\��x]��E���g�=���>���>��M?Mc�>b��C�t�^	�Nǿ�(��7����l������;^���Pe9�F�=���e���mė���h>�\G>BE>��>�]�=	�]>�F�>�4g>�]�<,O<���Τ==L�����;����f�� '=��м^Ҽُ��3+:�GP��*��:W#�%���ڙ�>(?X���C=� �!������$#?��>��>A��>�<�s��ua�x�T�T�N���?���?n�-?
K��>����­>d�>�6=roH>��ͼǽ?��ڽu�>�?^�>���=������G���K#��7�>���4j�j��?F�P?-�����%�����4�!QE��4<�Ԉ�����6Ԃ�XY*�B�F���޾�L�1����C>n
?׃?r����ͼ4��������١�Uw<=�B<{�?Z�.>|\c�	򉾟H޾7�=����= �Y>~��>�<<��?n�=?5D&?�Jq?(?��?��F��?��>#�.?S��>>c�><�>x\?~�c>Qә>&�%�e�=QA�"ꄾh�=���=���>��>#*>̚$�ј<s3��Y�=�8=~�`9��<=����k�=�zr=���=i�1>*�?"�$?��/�EX+�;=�Gk���=�	>��>�t�=���h�>�g7>���>��=?7%�>:�3=ㆬ�3�z���|�>�z�>�J=?�?��Η>���=�x�:�F>t�v>����Ñ��p���VO��E]I���>|I>9
�>UD>�\�??�Pm?hw�<�r�iu��V
�V�=K�j�?ʎ�>k�N;j���G��Ԗ�UHJ����3�="f��#�<$i�=�K�=;�O=Æ=��<��;s�T=- ��p�<(����K>�>�=?���=�����O1��Q?��ҾgR!�E	��C���ƽ�Eh>�{>BHn>h�.?�3=�jv�=������?I��? w�?ƭ0?H��=Ld=ݲѼ븤�B��=�j>sA�=�[">���
��>�w�L�<��Q5�I=��?�F�>��ֽ`u���q��	O�=ּ�6(1�d琽yܾ��e��䉾yľ��U�	.��X�Z�V��94���S���0\��H�W�0�1�����3x��L��?	��?�>O��=ܫ
�R�;���"v>K���Q����)-�nc���ܹ��Q��^���j��1O��0��2��;�>��߾#����w�RI� k=�ҽ>5�?����������;1}=��>̚�>_��l�g�y䉿v޵���k?��%?���Ѿ��*<��[>Br?�B�>sq<�I
�������K>^`m?-҃?�� >�2��M���$���m�?P��?��_?�g���@�����<��40?�ZI?Pڲ=ǌȾ���*����i?w�?G9?^m߾W�d�����v?��
?,/Z�͔�>�C�>#�Y>~|W����}���m�d�x%d>\!���
<�-����þ��7�쩟>��>�%��5�Ԣ>R��IiѾx!��p��uY��;����H�>������>8�����Խ'{��V�� v��z��(uA?�ڤ?~�f?P�j?��,�<�C!��{=�u�>f�?�p�>��>���>v�>^�Ͼ&yk�ȤG��Z3?��?	��?��?�b���ۿ����b2��|9��× >�`>�F>��U��=]1���=Ƌ�<%%>���>u��>��>�Ne>���=�p�>#т�iU ��v���l��C#1��"�"�/���{��5�����˯�����O� ��r�<(#ԼF����&���6=���ᡞ=Y�"?.�>(�����X= ��=E}��:4�H�W����U5��Ež���
�����
���%k���=�K�M?�񕼀�p>]E�>/w��k�=j�31]>�z>=�j|>�*D>���=@V����">|?>@��>>��>	��>.�=I�u�埅���:���I���=J�`?�����i��\����˾�򙾂ʇ>��>%�8>�5�%ۙ�DI��j��>Ȣ���?��o���9~=�!c>g��>l�=r�F��uG=J�m��MZ�]��=q�>b�3>&5�=�����7���暽H�>�T����=���<�#?TYn?�0?���	>d�S>�d>sM>2jX>�m�>�9a>�
?�<6?��@?*�>3��=4�-���+>�`��h���"v�Y�ͽIH#���	���>�p>���?�=�Z:=� >�G�=t>>�	�=�v�=���=	�>�l0?$B$>e͜>|���+K��Y�}����
�;��ȾTǁ>���>S;�>*F�>�|?�a>�=ؽ����v8�u��>�C>���w��K7N����>�w}>��?�[?���=J����ۼ�Y�=y~>�/�>�9?rN�>�W4�p�Դ�.ҿ4M�YD������������\�����[R�<���½$���=B�X>a|>y�l>�}>��8>3�l>���>��M>k~�=�|l=-!��ȅT<�Xh�v��=D�/�x�<F�F��62<�k#�C������]�U��n��Gb���?�*?v	���;@�=���?o*�"?69�>�/?ؤ>ـ>�S6���p��wY�QR�%�-?�^?eS?��o��2>��6�>>W�>r����>�=�Q���ʼ��?xד>|�?��=�=�
���e݊����ɿ>�O���[��=�?f�R?�<
�f&U�y	!���B�O�%�/�c=��C�B܇��e��b6���G�������:���Z>@��>�G�?�H[����=�`��v,����������g=%7+>E��>+'>C�'�Z"�����6{��P��>릥>o�ѽ/

?k
E?
 ?P0X?:!?��>�� >}�;?���p?�Bm<Z"�>vУ>Yk>Zc�=v�{>� ;�,u��h(�z�Ӌ��o�=���=�<�>��=ã2��]�;���_=��9�d=�w�=T�V=?a���
�B�}=�>�_?�=?�c����������Ԛ�����t~=vV=\�*�޽�^�<N�L>"��>"h-?^��>L�:���9V�o���0Ą>>q�?��?����f^�昮�a��!��>���>Z �����N
��(5����<?λ>�FC>�s�>UPJ>)P�?���>�!�?���=hT_��|�c/> ����
?;�q>�+B���*�IW9�\���XyI������&��=�3¼�1>�0>�K���=�Kg>)-���=���⍏=Eɧ�ȹE>VA�>�p�>TW=��P<��!���N?������'������N���[�=[�%>�>yE�=��O?eҶ���H�Aj��������>vC�?�y�?�?3���UC�=���8�Jsa=T�=/�?>�(��E���@ ?R^>��ҽ���������>�Ө�8f5��n����iwf�:�ſ��=�g8=ɾʪ̾�,��'����*��☾�T�X� �5~��g�����\��˹�����?�Ǿ����-���ϐ?`ʙ?��>
�+���C��M�����l�1>`}��e`�
�73��f�ɾ�S߾'eо�4��JY�/n� D�I��>���Kw���e�� �[:>y��>��>*҈�B1_�{�0�<���>�V�>~|L��Z��z��G:���W?E�?V�־(�z�zJD>=��>g��>a��=�������Z��=Bn?uB�?,�3>�隿���i���:!�?Q�?�y`?������R�w��	&���6?<�^?,�9�В���ʾ�m�D �?~�?�k1?�v�v�M�&�۾Z?z.	?������?�3�>��>ap���I��2m�.�g�ܽ@�^=��=;p��T��>����s�=~f�>Əe>aU��a��_i�>�ܾ����}"��� ��	��9j�j��>$�D�"�>o�:� �y`%��y��A2���s1�X�U?��?o$W?�w�?�9�$eH�8ղ�!ߋ�0��=e?l��>�	�=#<�>"�=
ϾoW���5�R?���?��?��?F�N�qӿ���噶�%��Ӓ�=>�=�p=>Q����=:H=��v���I��+>G�>��n>��x>��S>�<>��.>{x��h�#�����@���a�A�`��&v�QSg�K	��jz�=������>��'���u��m��PuF�ͯ�D�9�2����x�=�?��>ag`=w@>�hQ>܎>����N$����پ[P"�q�o�񾊁�>O㾗���۾G���4#=����?5���=�=-��>d믽���=�:H=޹P>��c=1.~>8~�=v>@
<;��=7~�<a2M>�+V>��>zۃ=�R��Z4��Sd$���G�ma=ðY?�)��+_�Ȓ���׾94���>]�? SZ>��'���U�h����>-"��q���7�]=%ͭ>�:�>f�=�f=�]4�g#����𽆭[>���>S�o>�<�����P��H<(��>Eо���=��>�l?��?73?j	�=f0�>��3>�>�x2>.�>GE�>(>�d�>�;?lE?���>��=
�H�(��=18f:4r7�ݎ�!6�\G������fl�����#=X���ZS�=�J�=�->��=A�=��=�I�>f16?%Ӧ>��>dvԽRJ���D�z�A����=���࿢>��>�϶>ͷ?���>�	s>���<�>l�?O_�@�>-Zy>U�f�s����F>��=��>�H?��?�W����
=�j�:�1�>	?��4?'>ڽ�+�v�D���ſ��	�Z+��szD<iS=5MW������>fQ0��֠=����R=vA>��>��>M��<�O�<�X}>Y��>�~>��=��= �1��`��XԻgp=RՌ�	Ӎ�N,ٽ��L�c��#���]��1���/��$�+h��B�?��,?�ǽ��S>�� ���Nܾ٨?:x�>�	?C��>���=�T���X���E��̉�Tv�>�,?d�>����Ј�=��ʼ~�V��π>�2>���>1�����MW}��-�>'ƪ>���>�w8>4��[G���������M�=�B	��Cc��|�?�<;?�4��+���0�;"��>�4�z,���LȾ1=���X�d�#� �n]���D>��?��?�*��f��]����R�2,K��!ļ�h>S�?w�]>lg��ڣ�� �x����RI<k{�>�?�m7��`?��<?Wi?P �?3p/?٨�>p$����v?:�>]Ł?��C>k��>�Nv>�X�>���>l��=M�"��\9�i��^��� ���2�=d '>Ў�>4+=�C���l�=�p%�<>q���?=D?�=��<�Ȉ=B�=9P�=�6>��?7z1?B�s������>U�ƾ��F�tP>T�>-��F
=���&>�t�=ػ�>�i;?�\?V��=��c�1Ƽ�=�3�Ms>f��>�| ?l�>H��=�C����;��3p�n\>�Zz=H��8�S�6�/�i���V�꼴��>��>5�:>6#n>��y?�&8?տ?³x����<XW��Už.[�ʽ�=���>1,�>�J��F�%'@���~���E��)����.h�����P<>�	>V|> q*>x�=R4��W볽Ϗ��r��<gV=>B�>Uh�>#L?j�6>��j��>��B�ܾ��@?�`n���6G���L��%��������>��߽��>~)���T`��2���Z�^�>p�?L��?�O?����qC�<��=÷��ܮO>��۽;L�K)�=���;�H�>+�[>����S��y���½>�Ɠ>>$#�Wy�����`$�X軿�K�wB ��=���=���2��p��������8��;Ϸ�O�¾v>����C�R?��I��������S�P �?v��?�ʊ>���:sB���������I�>� ���N�z���슾�>��U���%�ľB��#|2���G�@/���>����X��������k(�)��=!�>�F0?rɴ�����-���	� �>)��>2�*�JyJ�/�s�������?q!?�S��4%��)ɻ���>f�?M�>�j=���߾*��R�>�F�?-!�?�+>��)ך�o ��g�?{}�?3g[?���4�[�Fk�; �W}X?P+o?�,7�E����7�"�M�?��?��8?�-���S��g����M?H��>����*E�>Q��>>�8>I����
>�l���O���国8
��碑��!˾�*C���={ά>�R�>ʡw�*�ɾy�>�F�ž<�׾�!��<��_ս�,�>�11��O�>�sl<Fӟ��]�]~��G/l��s�;5�9?��?]L?�c?j�,��I)�K���K���w�=��>o@i>L>Pg�>k��>�'�C�n��sq���I?m9�?ZM�?K"?3�U�D�ͿW����a��M͞��E > �=��>�E޽>N��<=ڎ��
>�|�>>Bp>��x>��s>D:>:�>c���$� J�����H�C��G���!�}OU����h����X���N��[��.Ur��t�z�)K��������&U�>#�(?:`�>�?_���=�20>��S�p���w�r�׾�/�����#����%
���ܾ��������M�=�	ܾc��>��<�]�=&D�>IgK�*>��E67>4�>z�>&�B>YF�=��t=��>���>���>�*�>T"}>��=�܂��}��?�x�G�"q=�=?�Z,�wK~�
e6�������F�>?�	?Je>��%����q�n���>���yǀ�d��M�;g,�>E��>��=�<I�=�>�}���ϽO�=lI�>w>�8�Sg��H�f��=�|�>�|Ͼ>�=��]>�� ?,�w?��'?t}�=�/�>$�i>{�*>:M>�g�>A��>�'A>���>�oB?�+?W��>�
>e��~k>ϣ�el��d52�d�"�������<���*����K>z��]�O��u�=v�h>$�,><>���=��>n4?���>V4�>r9��4L��`R�5\1�Jֆ=Ù��ܣ>�e�>�F�>�
�>��?zH�>���=��\�8�C����>�>�e_��s�+��=>�5�=+^F?E,?M5���ؗ��M6=��=0<�>��?�=?��E>�׳=��=�
� �ڿ&�)��[���ɼ@�<�U�t9n�e�\>�#A��>I� �,����C�>���>���>�M�>�Z��y��;�v�>`��=E�>@�=�=m��=�ѼWv��iq���=� �<���;�ؽ$m��mͽ���|ఽ�qλ�h~���?\�?�D=:��9tF����������(?à.?�,?�z?���=�\�7�:��?�:�.����>P7c?|x�>o�t<!"C��n'���>�8[>~��> �ֺE�������L�>9��>�?��n>#�;���j��
��e���.0>���<����y��?[�_?`	�,K����4�q���&�=�@彡�q�����L0.�5�>�(����E5�jG:><%?���?����N=2T��\���^���vv��"�=M>��>��6>��X�Я��0_�A~����E9>>�Y<9|?���>��5?�W?��?]?��M=�>&?s���[?I�G>�!�>�f�>��H>i�Y=�D�=���<��5>�p�hg�����W@��G�=v>��<��=(�>��l�TX?=Yd���>��="���Aٻ=��:>/��=�8>7�>�D%?��2�0�D��~�>�Ӿǁ���ژ<~$���j���Q��]#=n]�=�<�>�aj?E� ?�J_>*�'���,����/s�>���>l�2?M��>k?�=���c�ͨ�7��>��(>�P��/׾/m�a��{MԽ���>�� >dX��{�r>uw?e3?Xl ?��d��'�qR�1� ����=ܺ�>!.�>S�	��a�#� �G
k���g� T2�=-�)ƈ�ɶ�=��>X�^>� >��>�fb>��(�!�v�[��;/=v&�S�>#ݷ>{��>+�W>��=�s��,�Ӿ�:?BR��p���%ɀ�į��@��\ q>B'�=�;�* ??ñ��U�⎿��
�?%��?�%�?��P?�F{�a:�=\�=����&���s��<���,>64G�Ǘ�>p�Ž޺��_闾^�=�n�>��
?�F�=�O�����^>̜����/��y�=3���2`۾�1��C����b���S���\��I �����O:���w�`�5����[�׾iB"�y�޾�T�? �?�ě>h�6<�NT0�`���`>��K��# ��8�@Q��<l���پ�Rʾ����tJ�bR�|�(���>_��D���H�`�*���W�=g!�>Ҥ?z�}<��/&�J�޼�{c>�A�>O�Q�ϟZ�_v���f(�h�q?��%?��UW���sҖ>�y?��K>Њ� ]���Ӹ����>��k?���?,B�>�!��dc���!�N1�?��?ܙ_?�V�US���?�j�2��O?�}/?�iw>�����R־(N�=g��?�6q?�v3?�Hݾ��m����9�>%&+>3�ʾ/�>���>�8�>b��}�]��h2�����`��\}=]R���Q���w������h��=WSp>UJS>;)j�s���|�>[۾& �nO�`�4��)���=��>b�����>�BT�%[�4�E珿�7e��4�0�Y? ��?Q�Y?R�w?�� ��.N�isɾ�'��oů>�<?
r>�>;	?2�>������J�}�ؾ�@?��? ��?F�!?HV\�r[ÿ�����Ll��uѾ�=v0b=p��=����I�=G�>>�n>��=��=���>U�=�L>�>Ci>�O>�`}����v���.��$�[��78�����叾(���z���M�PO~�cLӾ�9ϽGd_�ᚋ�o�[�[j罸��<*���AF>y��><��>�*�>�ی>�o(>\��P�"�.���Ǿ�����ɾӾ� ����� d�sn����D�<=�����9?(����%>�>ױC��[>z	i>�s�>��ؼ!Q>�bU=���>��=>�*>X�+>܀>�=�`�>:,�=��4���|,���l��p<��]?N���~���X#��s��蝔�ͩ�>��?�rS>B3�=Γ��{��4�> ���1�O�[4��C�c<�w�>BԷ>�J�=1�O�e�3�o��*�9����=�^>˽">ũ�<������J�Z����>v����@>�B�<�W?�\�??�z�=nU>�.> {n�s�7>g'�>
��>�kj>x2?��:?c6;?5�> &�=�����u>�=ބ��t�ֽx����޽�(I��ҽ^u�,����u��~'� �<4K$>:�>QDK>�}X=:J?�:?���>���>Joc�ens�G�,���s>:�>�C�=t�+?{x1?�)l>�ָ>�1�>��ｹ���"ɾ��[�YR�>�>>a
[����$"����>�W�>�U�?��+?�<������'> ��>�&?� ?J\P?Z�{>�M�<W���p��0 ��2N徖:0�xQ=[�H��i��gF��K=Q��=�Ρ���9s��=��=�T��=�Y7>Gk�=1�>�>s-����>PN=�>��;����!u��Qν �I��悔u�$=�k���=�J����<�ٷ�/V����?�,?)�=�u=�����ԾJG�p�?�i�>>o�>�r�>���?D�L�l��zs��q~��f?;�^?��>�pY�}��=o�c�m_v>cz>B'>[��>���X��I��( �>B��>��>)_>?/ �䪀������1E��H�>@+켊P�z�?��?=ϕ�f�4j!�;K�z�&��=�l�3*��=���`<���`��6��)��/���->�?Z'z?�q�+��<{`��,s���I�p.e����=�Ė> �>`��>��|�����
��-��2;0�[�b>ڦ�>��=4?p�?��8?�Ղ?	?�i�>�D�<��B?�7�=2A?j:�>�<?�}�>��?�r'>�s�={�
��(-�2�9��s�M�0�(�:�LV>�3>3H=��M��#�=�����=-�˽�e�;��%>ȍ����=P�>��>�w�>��?t9?�O�";��r��=.$�9�<�H>>w��=�A:��^�#<�Q>Ն�>� (?�>�yS<K�V	,����ԃ�>6��>C?��>�, �������ξ������=���=YH���uz����}�����޽�F�>��!>h��iY>�?�??�Q?%��=�(�I�[�*���I-=�
 <�>]4@>w�ļ���%�4�C�v�@[�.�S�#^��2�h|=}X�=㏇>��l>Pb���V>b �������`��e�b>5~�ՠ�>1�> �>,/h=�N��^��a钾e-K?���ka�C�4R�M21>a�q>
&+>1�=r�>E���ق�a�����S� ?�s�?�^�?Ѧ6?K�񼪼�<�r�=�ʪ��)�=�;�>X3���f����=~�;>�ֽ��C�.�w��=\7�>�Us>i�������k���H޼���n�H�����l�W�w�����(G����o�i���B_c���Ǿ�}��E����5�t
���U��r������m���|�?���?���>�8b�A��[���̽�=�=1�����W������9��^ʾj��9��3R�Ï(�ȣ �`ײ�/��>h맾�~��nPr��!%����<���>�v#?�ɞ��d�� (�۵�����>j��>'H�am�Lv��{�н%�h?I�$?$�پ�z�����_�1>���>��>��>V������W>U�m?-��?�>r嚿Fy��fzV�o�?�Ѯ?�S?��� g�R������ީ�>-g?��g>���Z��΅R��mf?�F�?h�8?�/��U�F�d��}?I�E?�/|�N,�>�ȿ>zsX>7S�z��8�j��LվT:=@�&>_�<�D=����~�����.���>e-�>s�=�;�̾#�>��澵�K��OF�:� ��x,�o{d<�X ?�|���K>���>P�>�9(�dx��C���k���[G?O
�?�O?>�.?�����Pԇ�ua�=��>f��>�)�=<rؽ3��>{W�>���0\m�$w��?���?���?��]?��b��㪿X���D���)����>5�=Y�a>�8��LQ=A�:>��=Ḱ�Л>i�~>�W>�*�>W�C>�UP>$�$>���j��ㄿ�O���13��#�y�-�A���;b�>�m�y���傄��N����=��e�8<�Ծ�����`��8۾t�=[�>vX�>vo�>��=>fҎ>H�*�vg޾$l���R���������$��yҾ/����Œ���5�]a�(h�����--�>1��;TB@=�b ?��=Չd=���>�V>�=�>�7#>�K>`4�>3_v>DNt>�k>D��=��)>Va�:.���T������`� ����=��?�Ҿ��/���H������H���߼�n?ga��C�Z�|�(Z���i�>���SR�!t��L�];H��># �> �*=����ׂ=�h���m>�U�c<��=d�;�%�f����uE����:�Q�>�;���f=��>�%?<In?��=?���=e�>k��=��=!Rd�J>�o=�F�>Z�J?{�a?ڗe?�3@?m�=�$��/��;xս�𢽺��<��>L#����=�u�9>f�8�[�9�y���뼉L�=��>�y1>!X�=-�,<}�?s4?���>_��>������Gg�˿��h-7>�����i�>�F?�8?�?Z�>"�5>1� �^�Ҿ|��?
�>B��=a8i��S%�7�P= .>?=�>Y[`?�C?����������>�s=�=�?��K?��>�_?��	 ��!пD�/���$�����=��@>�N�G�=�x>a���H����^�>"'�>w�>2Y>�z�=V�3>��>�ut����=A->85̽�[B=k}�����\*6���=�����=�}��3�=�P5��g4���Ͻ��ϼЙ<�*?�0?6M��xu�VE8�ts���������>~'?쪺>�>�W��!پ�qT��NS��l�<^#!?��w?&-?!��,|D>�<u�&&>�
�>���=�(�=0*�=��@��Q�a����t?��>��*�8oV���U�����>��
=5�.�B�?h�X?�!žbD���=�L�S�����=g���%0a�7s����-��PF���������,�<r!�>?�?]��[��<r��<�$�����Fsm<ǯ�kf�>|�>��#> ){��a��6��;���۽9�=�s >P��>A]?��_?�!u?��?�n�>n3�E>�>AO�q��>���>�I?9&�>XU"?�̌>a�>�^>��a=u^�/^v��ɛ:p|�=Ft>�wL>l��>"AǼwjͽ�p�<�P>�G��[/�s�6��h�=���<��=S�>���>�?�"?�&ʽ�e踾�+;����I�<��>�t>�����_��$�;ͮv>��>"-?8��>&:�=�ϻ��ھw�����=�V?�38?R��>A<�v>z0ܾ)Z��Tu�=-%?>Nd��"֐��t������ؾ�X��>�A�>XJ�=�ۆ><��?[r?fD�>s�&�%G־�q�g�1���� >JLA>�i�>��>�f�<��X�~�|�j5�c7c���D0C�yܤ=��=��=��9=��O>�o�<�j�<���������>s���>�>v?�S�> Η>�z��D����q�S+K?X���8�ר�����e�<N9X>s7>x}���� ?<�U�b�����D<����>lN�?Y��?�lo?/Rҽc7�1)V>iU>>���=LE|<�z(�b�ü�����l2>�4>��n��{���V�;%�>G�`>[�"�����ھE��nH��ũg��b4=i����J��<
�|U������̾OSn=�׆�!pg��;�tz>S��dD^�r;�����Rھ��Q?�~)?N��ή6�LU2��?_����hv�>μ�����mw��%W0=W�ξE�����Y.�\�8�}^#�λ �I�>�`{���$Cw���)���p��1->l9?���~T��V����s,=V�?����N������ث`���'?��?K����~��"==.�>'�?jk�>��c�te}��>7=j?�)?��;?���T��GDw�o�=��?~0�?��??��O��A��!�Oz���??�?�E�>@� �̾<��
?w�9?�3�>�L�Z���/����>�L[?K�N�vb>�T�>㰗>��@(��wA'�v����e����:>+fŻ�����f�9>��x�=Q۠>\�x>H+\��֭�_,�>��龅�N�F�H���v���͗<�?׏�>w�i>4#>��(�l���������L?K��?ȮS?�S8?|������DZ��x�=p�>뭬>�H�=�8��>��>ņ辞	r�����Z?@�?e��?�EZ?�Pm�h�����������T؆�,*>�p�=�:h>�-н��>L��<���<B�:=���=���>b1L>�Fe>]w8>2&k>�<K>d�������Γ����'�[���A�Ĭ�������V���&�b�ν{���a.=�}��M�`�����瀾�\�vȾ�z>Ռ?J�>��g>��z=��>N74�����[���p���#����v���3�¾*�������h��9#Y���J�-��9�?��=>��?>����<:,?\:�bc�>�!��"�C>���=�$�=z7>3��>؋�>_8>��=ұ��g��J.������=���=p5�?�k�����*�o�OX��ٮH��K�>@�7?�d����#��I����a�>ɑ��0髽9B���9<�3�>�4�>E�U=�#���va>n�g�����ԥ<�SY=t�<x򽽥��i�����>9w&?�:½9b�a_=`�5?LЋ?]yI?�w>�:?�����0>�Ҿ���>�3>�&�=NJM?��k?� o?� ?���=Zyc�h�>u�G>�6Y<f&"<1����O�>&���{=��1�Z =m�+>�2h>d!>k��>��=Z"�:�C=��?��)?��>��
?C�H��T��5�Lfk��I<>E��B��>���>`?~=�>���>o��>��<�o���d����>��t>x�m�����ˏ��r�>�>�7p?��k?ҫ��E������+��A}>�X�>i-?:�?��>=>���2�ֿ�<���_��u9<��e=�7��͚�2�<� ?�7���7��c6>�2�>�kf>��;>wy>��6>|��>3�> ��=���=M> �-L� ۬��iu<q)7���=5�8���6=JFA��Ԩ��5���h�^�_���S���=���$?�<)?)"�\�(�QOY�1�ž�����>�>
?Z�>���>ƫ~�ھ�m`�%@�<�	��<?.�s?-�?����=� ����O��>>_�>-R>�"�<��	T��9�A��=L>{�?s�>�nP��E��S�9�����>��˽��p�%�?,�U?��оs�E����פ\�o��L|3>��M�����kX���j�:������L��Y��'{�=;@�>WԿ?�|c����<3ѽ�򏿇���'D����A	�2$?��>��z=�0��{�?�vO&�,����u����/>!��=w�a>4�?s�J?�[?��?�p?*G��P)�>M��=F�?��>y??�/?DϞ>���=N��=�@�r8�|g��\3=F�=S,ټ��i>�8�>�ҕ�i��p�g>^P��Ӽ�,�=�8�<��f�G2D>.��=�V>�)I>��?F�"?��۽3}Q�9��j���;
=�I�=OJ>p�����l�"\>P	?�-?�5�>U��=�Ӿ���V� �PM�=�? 3?�e�>*��;�=�"��C��M*�=t i>�#g����3��#����j��7>;�>ͼ>B�=Sm?�:n?K?���=��5��*��+DV���<�Ry8>/V?a��>�K�>(���{��@���D���/��y�<�5e�����<�[�u>iSB>$�0=�� >X�?>��;��Z��=r{"=`B%>T�t>��?�V>�6>=Ј&��ʾ*K?����,�
����ξb�	���>�?>���>H?a��hz}������Z>�Y��>�\�?7��?C:e?S�5�V�� �]>�K>�>��q<��1�����+�h�	96>���=��x��盾-�<��\>�n>h)ƽPǾ�ܾ�E��s��;x���߽n���D��23������Q��O�Y��}���;즽鴾�(	='���R�@�,��������X?`?�N-<U���Kb���,�
���(>A���"=��F�>�.����þl,�r��a�
��C;�8��:�>IU���4�}��.�*=��n�<>�i1?��f�����"�K�3=T��=_�<0�得��������D�o�J?��*?�~۾�|;lѦ�ʜ3>�
?�}�>��=���5\彙ɰ>�#?��4?�������������u���?�E�?�/@?jP�A�,�)���	?%?m��>���W�ɾz��8	?19?@�> ��鄿]$����>D\?��K���a>���>00�>A���ד��D+�K��U�}�#y:>�D/�M+�Crb���:���=��>�z>!]�����|V�>��žZ>B�Y�P�����;�ʥ���?�D�{q>$$>��>�0�ȏ��d*���#p���.?Y[�?͹O?DV?���-v��v����>1��>p��>��=�񠽏i�>�d�>�ާa�Yپ]�?h��?��?cZ1?�Mi�Gۿ֨��AT��6�޾C&�=B��=^9?>M��g�<��~�t�<Uͽ㌥=�)p>�y>�>�:>>O�m>PL6>�����%�De��E����\��b�7��JZB�S�䆾�I�w���1���ڶ��}.���d�/t;����=�����N�N>���>>>7�G>Y?>�`I>Z�>��r��T1N��~x��F%���վ�dȾB��k�پo,���˾4�a��}ɽU��'��>	y�=��EL�>
>H��u�>�%�=�Ӌ>��7>J��>���>G�k>�>{�.>�>��=���>�87>2��(}��S8���ؾ1=/�h?h���&=ھ&e��儾�,!�#ֱ>wB?y%�=F4������㑿G�>�]�<�����/��\��c�>A	?�NU>��>�uY��;�挾>w>QG>���=�С�����T#����=@��>��.�������g>G
?�Hb?T�e?��>Z�>}��>���>�6�b@�=!��d��>�?�17?%]?e&?5ik=}����fY=�y>���:�x��"Y����d꽐�=�K9=+�U>�CֽK�q<r.�=�:�k�Z��л�k~�m��>Q�F?T��>���>_��"�7�H��+���~>;�ν��>���>0O9?�GQ>L��>9�>`��=���%uξޤ�>�9�>����Yċ�iN��Jۡ>z�z>�uf?�?%K�=)3���̜��P����C�>�p8?�b!?�1�>�;=*��#rӿ��#���!�#x��X'�r��;�=�)�J�"�:Oj-�����?�<B\>3�> ap><�D>ǣ>�K3>�S�>t_G>�x�=�$�=��;��:�wH��\G=�X��;<��Q�,���Iϼ{8��2튽�vI��3>�E��
��?f2*?��&��z�1�T�پ������>��?�>�F�>�G{���ľ5sZ�d�K�^j�~�?p�g?��	?�}H����=r�1�����&�>
@�>gc>%�½��!��F�K����cP>F�>b*�>{�󽣞6��E��P��?��>�q+<�Ĵ��;�?�P?���/~��p$��`�<����=�ͽ�ӽ.騾���A���+�����h����9���>0V�?@�����u���x��W���܌�w�ﾳ'��ML�����>&�>����_�y�����F圾s�*�<r>���=8�>�/?��U?� J?`�>�C�>��K�h�>���=?�>dD�>[�%?0b�>��?�9�>|�~>c"B=�1��G���~N�{�<A��=B�>*�4���>y�U>(c-�ܢj��B�=�b��%">�X�<�,=%͛<�?=tv�=2N�=|u?��.?QsE���1�y�<���:���=�P
>Gw�>}+-�Q椾R�_�E|�>�}�>��(?rG?�؄>l�p���������v֯<�??�R3?���>���=�uE>k���2þ��>=��=����-����mY]�+�]�e��>���>p��=��*>�?:�p?��>�߇���۾��x���k�8����>���>�Ǒ>K�>���E�^�������L��B�`=8��Ny=/O>rD>2�>�9
>�l=���=J��;-b��!h>�1��G��>1ի>��>�zc>�f�>�Ք�xz���<J?隒�L��
��o�ƾ�S��j>�?>��Ž%y?���Հ�p�����9���>��?-��?��f?�u%�%M�7:N>�`^>S�>��<ݸ(�Cke�����<>���=4�v������!m�Ehc>�w>����{LȾ_�ݾ�&*�n�ƿ���.p�>}�<@���B�H��%��ɼ�U�!���r���&�}��>��ɾ<�>!����C���H���!���L���o?he`?V��=C�������#��־� �="Uz�/����O��C��=\H���O��"�Į}�����(�������>j�)��ņ�r��Z^��@W>R�L?��5�w�2�A�f��J�=�ڏ�eY�����
5��4y���S]��)?�?纾"�v��R<Y �>�-�>K>,L���־SL�q!�>[� ?�?�a��q���HR�D	�?˲�?�>?�&��A�[���H�� �>���>��>9砾}N��T-I��r?�?�9d>VF�������)����>�Y?��u��tZ>�?.?�>w�<�R��{�ѻ��2�нUҕ>썵=P�(�z�k�ۘ5�� �=���>�=�>�i��$���p�>ʕ۾n@L��'D�{0
��6�xS�<m��>����->�+c>V�>R'/���������G!�}�??ߥ�?��F?�P#?���/�о�)����=p�>�6�>�7=
V ��N�>`�
?$�y_l�v����?R�?�?�W?�Qd�]-ѿ~c��%���ξƾ��>�a�=0}}>�X��;�=d�=q㼖-��� �=F��>��>�KJ>I*B>�n`>�\R>������(���Ɋ�%9�f�-�Ʃ+�����!��V����
ܖ�o��Kn=���e���"���x������+پ�u>Ӓ>*ϕ>���>�q�>�>�4�խǾ)��Ӝ<�H����kv.�Çq��{��Y�*�xjʾN)��"9�V�Ͷ�>�-�={�>$��>G=��d=$�?�ʔ�|�#>�'>��>��>_&�=�n�>Aqc>�A�>��=.�>2�S�����h��ka��j���\�<=�{�?�'���a��1e����*�4�9�>��?�����?�����~������>M�;E9�j���"oo�	{�>%�>A?�=4�);��&��۾��>�;'>c� >>���O�;)H#���ƾz�>o��>4Wɾ �=��b>�NQ?��?-Wj?���=	��>��>DQ?%�P�s:f>���03 �y�?fh?�)e?��>?�ʴ=�I�����<��ټ����;���x���T�=�^�=�>����5[<��D���}��R�;�h=���;��(;�H�U�?ځ0?n�>"?��E����ŹT�ѹ���,f>�6$��/�>oj�>��<?��>���>nK�>I�,=����O2�l�>���>��U�ᒿR�l���O>�]u>t�?IM?�r�������#�'��=�I\>e�>9U?,� ?Q��>ݲ�=�b���ӿf�#��� �!����?�;��=���B����;�-�l	�Wo�<�TY>���>M�o>�C>50>IG1>"/�>tB>-e�=N]�=�j�;¶;��A�GO=20��+�;�Cb�R3��:�����Iz��b�<���H��2 �G]弫	'?�Z9?D5��D�V�O#��`�������$?F�?c�H=^��>�z�㼛�� ;�E�M��'�=��?X�u?�0?���rY�=�	���=�q�>.��>�k�>�]�=ѩ��Ī�I;]�@�*>I�?FD�>�$���w�+lI������]>u=�n�����?��V?k������\�
lI�+��Ă����/���}ȧ�^��ģ �������.��3�G��j�>Ѽ?G5�bA<ĺ��m����ד�]�ƾ�Fd=���=���>���<q��	�&t�����ّ����/�p��>*�>��>L?�.??�5w?�/?�c	?��5��?dD4����>n��>��?,h�>j�?ob�>�F�>IL]>N4�=�3	�6򴾀��<�#�=Ŝ>���=�9>֖(�]ݡ�V�����=�4=+b������=�<��X<"3>T>��?��E?Ab�|ҕ��3 ��,=3��=l'�>!v�>����d���h�ƾgݢ>m�y>�t-?�)�>"��>��ýv��9��oA�}M,?�.1?��>x4>ѽ>u4�V���M�>���>��T<K���8����:)��Q��> FK>�n>��>���?�@I?~�7?n�u�˽پ&���u��f9��T�>���>6V�>)ٱ>;��>����B��e�o��2��sؼ�sͼ��|��[	���>(�0>	4�=����&a���]z�ğC=V��=�ޮ=�-#?6K>�:z>)�>p$�=�M�=�t%��-J? 6��[�i9��>4о����1>y�B>�����? �
�G:~��餿��<����>P�?F��?�d?��>�C���t\>�,U>�>��I<u�:�y=�Gv��Z5>`�=n9z�a���oϴ;�^>�|>nӽF�ɾ3���FX�A���?s���>9�`�w|k�	�@� m򾂉��+k����>6|����>ug��UU>�@���\�7��'y����'�Ɂe?�L(?MNr= �z<T_���@�>3�þ�e���w���k>n޾�!��2�l��!�.�UJ0�GM��ì>+�X�������*[5��F��FtA>�9?��Ǿ�S��W�:��(�=.ސ=���<�����n���ӛ��T�M�??8*?�P;���� �9�9�>���>��>;�=c7��J������>��.?�I,?�� ��	���a���0��ބ�?�2�?�@?j�B�m�E��l
�P�-�α�>��	?io�>o����ξ�y&��{?g�.?��>�*��e��� ����>�S?0_�Lk>v��>]o�>��ҽ�{��_Q�:Ǟ���-��\>@&=!���Z��j���=�4�>�N�>�\U��Ӧ���>�־�UQ�f�M���\�|����<�X?�߾փ�=>�->	.2��0���ʁ�#/罐K>?���?FC;?�<A?�:Ͼ�������	�;���>�/�>��J>^L۽�I{>U�>5���Vu�����g?@/�?¸�?57X?X�e��,ɿ����N���M����5�=U��=2+>%i��}�3=8[�;�Me<r�\<mg2>gĈ>��;>��\>s�<>�R>.  > ���d��Ֆ�Iy��Wi?��C$�Y��H����|��ϭ�ْ��W���+���m���'��Eݽ ے�+z��*K�r/��F�>�հ>�C�>E�>�c\>Ol�>�Q-�Z����K��&�@�ۮ�>W���!/��i���@��բ����W��.���C�{
��'�>�T!>Xkp>k�L?��>�<�<A�>��<>�̗>�L�<���=㲯=���>��>wx�>��>�$�=�>�>z"�=�f��(|���~�t�����?>|J�?|!~�n����x���ǽ�o`�6�=*��>�a�>���4h���֎�t��>l�#���*�_)��S�=���>PM>�/(=����L��������f��;�=1M�>nF�=��z�6z���e��?=�N�>��#� ����Z�>i�/?�!�?	#c?�0潳�?'��>Є�>���^�>#ܜ;=��>��?��I?'\_?1�1?���=�}����=C�>^X�J{��	�͐��_zl��7�=�����)>�{���=b'��%b���s����>\V?�Z=?ԝ�>���>؂d�����NG�e>��q��>���ǘ�>�`>�2?%�>�Z?�SL>��=��|��-��v�>"�>�O�QO������>��>KN?��y?�9Z�BZ�!�\�B$f=�CG>(YP>��P?��>n�_>z��=6���ҿ=�&����d����5���<��5�W]��W�;�)������
=%X>6��>�us>�;>�; >��0>d��>��1>p8�=��=��ʻ�����R���Z=+�8�w�<UV��.q<�y߼�0��y��fp*��K�v�U���I�F??�~?g)�﹌��@g�����=骾��>�Z�>���>���>�z�=z��1�T�%�@�CPB����>Bhh?X��>e�8��#�=\�3�3�'���>��>q�>K�^���������3�<�#�>�g?�a�>{�%jZ�t�n�t�	� v�>]�=xk�Q��?�X?vѾ�%�WQ��ϿC����^<@���T\˽�)������I�r�!��K��ʋ���
>�;�>c�?9��
�;<e�ㄒ��<��>����g=0�r�Ab?�\%>�H�=$����"�<���a������f >j1>���>��?X�:?�h�?�?e��>�L��k?�8�='?�O�>��?���>��?>�>mG�>��n>�~�=A*׽ ����	�<�W�=@��=���=�^j>ׁ�<�{�����=��:)��<˺ݽ$R<��,>Č=��8>�8T>tX><�?�T%?��Խ_���ĸ<d���ȽK�0>��>PPѽ.�T�W�T�H2�>��>��'?h׷>���<A���
Ͼ����<wx�>��6?�8?d��=�4>��ݾ11u�o�����>��"=AJ�Ƿ��ś�c ����>�(�>� >j1�>,��?�*j?t_<�������}��d$��`t���>�ue>�ri>���=�l�����v��i-'�O�Z�������aj�=�;�=��(<S�=1�=6Y�7x=w�;��=��ݼU�$���>1��>��?���=��=
�+1ݾ�I?4����j��]���Ѿk���>��B>���E=?{?���}��z���@<�C��>���?Y�?��c?�`>������[>�T>��>��[<�8�X
�������1>�D�=�pw�\&���];R[>�s>�qȽ�^ɾwm�<�X��߿�AT�-�>�c�2�u��"(�S_��E��˕���Ⱦsxؾ��>�r����>�0 ��'���C�r�����jB?�:?�����T��X�%�LR4��,���%x>�����<�^ɾ�	�<���:3���`8���������F�/@�7L�>m�1��:��;y~���,���f�>>z4?!ܾEž��>�T�Q=�3�=i�<������bF����^��-2?�.?�iȾ� ��<v���XE>�/?���>?�
�9����ĽR��>X2$?%@?�� ������W���b:�j�?r��?!�??W�O�c�A�$�^C�4�?�f?��>+	�� �̾������
?�9?�u�>��}r��O<��[�>nA[?�N��Zb>�R�>�×>n��[��p�%��ʓ��+��!9>�F��!`��Mg�3?��{�=n�>��x>L�[�.-���A>�_�����A����Jҗ����=�Ά>�B��'>
H�<o�<]���膿������<oÃ?���?�?��j?_t,� d+���Y�v ���/?��?���=�]���M�>��>fm��	�J����hV?���?�<�?l$?��3�Fط���|��\9��[+���/>U�=	Mm>�ҵ�g�~=��5=������=<>�X>�y.>m&>*�d>dp>`�<����7���� ���6���F��"������(E��b��1?�;�辘"��TS��K��5����:����������,��V�;W�?f��==�>�8=�s>>݋�~���ee����nA����A��I Ѿn碾�Z0���%�a\=����=M���L?��E�"R=]~�>������=���=��=���=ߕ�=%e�<��e>� >�E�>���>��>z�����
>���=�l���ʎ� ���mＱ�>T|2?��뽧q-��()�ĝ��򡾲B>�Z?R��7%yR�+`���x&�	8�>�aĽ�=��o����s�>�*p>CR>����m���q�*�K�`w\����=:tU�p6D���=� �5{?��-?�J"���ҽ�<�>f7?f�\?�0U?|�%��J�=��?�)>4G$���?�N%?��?��?[P?ӱ?��?=փ=%=v�>�>K�>S��P
>��=�4�=}�6�A���iY>��>F9��wv>��=�6����R����>�b	?׺C?㰕>�?	��O�sH��y�=t��>r���*2?�o�>��?/�>.��>p,5>�h��3��U�8�T��>�	�>E�l�Lqe�f�8=f�6=�C�>۸m?�7W?U.�~n���ŭ>�)"=�w>Z��>�*?���>A"�>��=���?HӿX�#���!��\��R���;=�=�aR�੢���.�������<&9[>rn�>/Yo>3�D>� >,P3>�M�>l-G>Rs�=�֤=輲;���:6VG��`N=.��� A<IEO���»͉ȼ"|��U܊��!H�U=�,}�ؼ�&�>�7?*�F=RN��}�F�!���.��V�>k�?���<���>ڬ�>+���v$��P�.U���>[d�?T!?E/��=����n ��ȫ>SN>	i5=XG�<�)>�+ֽq3>��)?�d
?jJ,>z�Ӿ
#x���k�V�!��4�>s�=U�����?{�I?2I-�H<Y��h'�x� u�"⯽��������I�Ͼ����]��徵�徬:�z� >�p�>(�?��L���x>L��d��un�����օ��S$��x�>P�Ƽ2�C�TJ��)���B�T��=�V>�Z�>Cj=k��>�� ?�$?\�P??��>@�����?���0�>���>�w?���>��>��	>�>�*<�Jʽ�O��s���=��ֽ�Q�=kq�=A�l=z�9���=�ظ=S8�;~�;���C��=e'�=�P=�U�=��>4yH=�H?\?��\��o�d�&��俽�>c2M>x��>���>���6��=`{�>5�?l�=?k
�>�-��։�O��l����>�{�>�ސ>+{�>~��<����k���I߽����y)>�b�ɫѾ����¾�,���[W>��F>�kP="�I>��q?��$?�?�K����e���+�М�>l����&?�@?qYE>����lW��+n�1Q��J=�+#�=��׽�����{�=�v?p�U=T�Q=��A>+E=Q����I=�/>^w����>t�x>B4"?�	i>`!=����B-�E	O?;9���X�n]r��>���X>-��>S�'�WѾ�d@?�ǉ=�Z��~��2�۾k?�R�?�(�?JG?��ľ�=�y�=ٓŽ\��=�i�>-CD�	���=��B>�X�>!�F=���~��="I5?�o�>�b���:��-G��c���Z˿��E� �2�˫����n�@��󄌾$�b�bk���`뽵#���K�+����q���]�MR��gvh�dFT������Sm?�U?Z>d2���Y��������#.��о����B��!�j�Q��!�վtξ�t���4��I�W�˾#x�>��X�)����}��(�ꐂ��n@>�v/?'�ľ����h�:�[=��>���<���G���B����"���U?{8?;徘S��X�ͽ�q
>X�
?G+�>ie">���a�>�>��/?�+*?�Y���
;��Mջ~�?*h�?o�@?~vu��F4�n��B9��?g�?�_�>;��BϚ�s�"����>��I?#��>����Vl�|�����>3]?��V�z�>g�>A^o>%�F������b��p��V%���=2������}��G��>�=�r�><_>�i��✾T�>Y	�	����(������%�[PX>��>�-����=�>��нnM�и�����u��=�� ?�6�?H�6?'vl?Ps���QL���۾NW���>FL�>TO�>��\�Qw�>�ڋ>k0/��tr��p־֚�?e��?!}�?	E,?e�c�O,̿��������>�D��=2u >���>��d���:���>f+a=���A�>�̐>��>�)>���=K5�=��T=���&�^a���]V�r�&�t{�Q���AqR��5��Ƚo)��t��CB��䏱��^,� �<N�C��������t��@>i�;?tj�>
�>��<�Sy>@����E ��1о��ξ����� ��:ھ �*����wм�1،����-{��ɾt�?f�=�B�=���=ټ}��pf�>nT�>,L�>̠�>��6>���=���=C�>�;�=;�>.��=��>���=Ç�/����F�tfѽ=�j=q&I?<r^� �v�
<�W���ƅl�>'�>f�?�B>��%�46��eB�� �>޿���?������<����>���>�r�=r��=�ڽ��S�6Y0��B=k�&>��{=|Χ�_����@6��&��l��>F2��D$=ɯ>>!�(?JEt?ES?0]�=X��>aG;>�ޘ>�)>>�nD>��Q>C��>�� ?��=?��?A��>B��=�����g=T���4���T���sν���:���<�|T���꽺D6�xBF=�H=�� =,S�=~Dۼ��<��+=A��>RK5?��>%��>S
޾��0�h�C�JrT=00�>�S�=�FF?�?A?v`�>�ܣ>v'�=.O<@��~��}�>�&�>AM�;8e�dDn�5>@m>�}?гJ?��T�Ų��4��Q�>���>�k�>Ӿ"?���>��>�>���㿚��T>�#���
�3>)���7A�RX�>?.n�;?h��}�>��>2�=���>�B=(T�;�J>�#�>l�>� =ۣ#=�
x��A=wK��t4\��j�=����d_ ��6�=���=S��M�$=y�ռ������=&��=a�>F?_w��������o��� �<�.��>���>���R~5>�N	>w[�r�d�)����4�Go?�N�?x��>O4�>� <zFB��|�=���>�-{>����O>y��/����B��_?���>\�����Ľ:�S��Y����S��>1�^��i߽�J�?��Z?>ǯ�tNƾ����VfY�� �`�	�����������4�!�U�P�����b�н��A=k�?�<v?�lr�M�>��־b���<�i�ᾭ�d��EZ>���>����j���t���1��e���=���>s��>9Џ=K*�>&&�>���>��w?��J?)��=fs[���Q?k�q>�1?��C?.X�>�Ϛ>Jw�>܁���	?p����
�X��k9����뼎;���m>MS>[Tb<�[�EdԽ�'��O>=��<%�>�:F>��@=B_�=�R<]<sH>B$�>v,?5U������ ��<�n=?�S�>�yl=���<*e�>�,>���>�,?�>��Z>��ž�X; Iξ�G�=��?R�>��>?��=솽�����g�^=�i>��t�:���p!����þ���=��>+T��l>�^?�c$? C6?s�"��B��\��W����zܼ4��Z�%>��>�+������/��i���m��@>��r��h�Y��<L�_>�c=\<>�'b>���>Q�������q=H�1=��׽f�>�h?��>��=F>=+���J�yCb?���U���ܴ<����SVo>�j������?%=��������Gc�n,?""�?���?�9?1���D�D>�Fo<jz�ڽ=��f>��;>w����5V�R؅>b�X>��:,	���=�~_?���>
���#|�:5��1� >�
����A�5黗q��B���4������[�����1t�($׾��f����d}Y��[P���a�wK���찾]ӄ�8{�?�|?Y�a>=>��2GE�݁���y��g
�R�	�+l��`����Î�g���*��?\�\�3����ܬ۾�D�>��������{�G~�f	�J�>�e?��Ծ�Xu��[�1��rk>|aa>(��u������a���c?�'*?�ɾ@�Ѿ����2i�=�(�>z��>2;�=3I�;#�Q�0>�A@?�M?Գ��Q'��Z6��E<D�.��?3?�?��Y?����7g��O&�ݼr�<�>c^?��>����מ��R�	��=��?/�E?_�<=9����K�T�>�Ԕ?B&��	q�>�o�>s_`>�Ft���������=��$>ڕ���g�s��<�u7�b�ؾ��:��,=b��=�{���~��_�>4��t�M���G����P�!�왂<hl?���B>�@e>t>�)�����������L?���?�S?7D8?���������ό=a�>"��>�9�=%
��0�>�]�>0��'r���_?r$�?���?*Z?A.m�\ ��������o\���>=z�c>e����=�G>`^!��7�˫;=�|>>`��=j�>���=v��=�L>(���v��ځ�������'��S)�Ik���ξ E�����};3��پ�!ھ�&2�m�����5�v���t���=B&g�GM�AB?-��>�?�����=�����WX��I�)�^�'��N"�����l�Ti9����<	�==T��xbK>�W���N�>kEs=VY�=�vZ=8�������v�=�>F�=�eE�!��=��h>�s�>�m�>�`k>��>>��=��>fK��|�鿇���O�7-���>�A?iٽ��G��� ��.�����xf>��*?j��>�,6�ŕ���D�~a�>c~I�Y(�Xr�|�:>d[?�P�>J�R>��=<�5�:�����)>�3?PZ>S����l�lK��եG>���>�U��FZ��G8>��5?L�d?(�?��=s��>���=/#�=�	�=��>S?>��>x?�^??pB?m)�>!E >��U�5T>�F�=T_����8�!��4�:��^��sk��5���[=W,=��t;���<*>� �<���;6N>dK�>;j9?Y��>	[V>��r9�K.���r@��?�=��<�X?��)>(��>K��>@?wx>NʾU�Jt�k	�> v�>f�U�����`>�>�>L�w>Y]A?��?;����b�����.�Uu]>kV?/�6?��=Eα=�h�{��m5ӿ֒#�hs!�Q��]���~l;ʻ=�@N����\�.�{Q�� 4�<NA[>��>L�p>kE>I� >�[3>f_�>z�G>,܄=U$�=��;�"�:>E�y�Q=�H�'mA<�rP��λxUʼ���K���B�C_9�;���	ݼ*W?�?��Sڐ�Q���U�|������>�3�>b�><��>U:�=�A	�D�W�u�?���B����> �W?l�>�rE����=a�P���<���>mT�>��7>�U���ٽ�c���<<ѿ>�
?_:�>�,�a��j�����>�=k�<~�?K�i?�9��Ic�}���Ɏ;�g[>�r�����������R��~u���n��`�/�&M1>ʑ�>��?J=˽��b>V�!�z�����D��3cȼ*Y>h"?W:>7v=,�fվ*���K���6Q���>8C��
?,=�>��>ʺ>A�?5�>s'M>�U?�1>�K�>"��>קW>���=�7z>�R���P>���=�,<=��:�۾�H5>p�F���#>�]>�I�=_j̽�^y=��=m�=�{��6�����=�HH<����i�<t��=��=}��>�Z:?�����D��;�\=,L2>�4a�>`�>��E���>��2���T<>�>�z/?��?/�	���A�� ��eؾ�� >�?��@?�Ӯ>���=�>��|�n=`k�=��>�;���3���M�<���>���=��->l8>ɤs?�/?d�N?dcH�h	�:�h��Z�dTy=f�='L�>b�R>:��m�޾D ���[�J+O��j:�uf���S���=��=���=��>�,żh=>�*W�ݬ���8W�]�=�}��4�>��>+�>�,"=��ི쬾Mz �I<?�q�]�ھ������Ue>)l�J>V>��_?�>�T��b�Y�灢�m�7����>F>�?SI�?dH.?PS����)&0>^�6>[�>l����v��S>�;j>�73>�m>ق��)�þF�h<�u$=��2��j��ɥ���꾝>��J��<F��:�=񡫾:�t��K�Ki��'����Ͼvhl���
�P���1U���P��X��| ��z_������"3��8�?�?�u�K3��.=������\x����=�s��6`��X��$%���l�<g�rʽ.�ݾ%� �oI(�k����>��	�E1��$�C�Z�ھS�����>��?������=[�.�Ҍ�^��>�պ>�U���X�{���lPX���{?�C/?��7	���\=�(�>ʟ�>}��>�H>�,ܽ1�[��Q�=�;|?9ĉ?��Ƚt���쳌�����?��?z�^?�w9��~r��� �6x��=��>�RD?I��>�%���O ����<!d�?z��?9
*?�u�t���z?>jS�=RÈ���z�4<?�Ք>d�=+�*�� �������X6�CG��@��<;�<��T��堾��<���=s��>2�L�9��59�>)�Ӿr5�uV�d��H����$>�n�>w�
���>��>Q�����#��������^)>�m?�V�?�??g~N?�������r���Q�<&C>��>%��>ݬ����>g?��u+X�����;(?���?���?աv?��d��/޿�����u��Լ���[�=U�D=
�,>眫���=�i=��a�̀=��>���>m�8>u}�>���=w->�jF>N����w%�n��(g���GH��.�ȯ��C���.���\���l���0\���Ӽ߽��Y�� ��O��>.�V�$��<�>���>�ō>��>�=�=j{�=jJ���þr{�����6�G���
���
*����f�|��;�P��e�>���9Ѿ�l�>B>񼔯">���>�o-�j3>_	�>���=ӧ�>��N>/~F>Ͽl>�ۺ:b�>���>��J>-а�]�{>p4�=s��8Q��k�7��<H�j�<�B?��Y�д��*�3�f�߾�է���>��?�N>�$������/y��!�>�zS��6Y�H����k<�H��>id�>�x�=�9u�V�;�v{�D꽛3�=xI�>��>4�l�~#���4�C��=���>f_���Q.=�|C>��.?��q?ҭ(?Q�=-#�>��U>�^>��>=pM>'�Y>c]�>��?��6?��/?��>�b>,+~�la�=�X,=�(Y�i��8v᫽�������eh��\��s
�=W��=�)�=+�=��<w��<
�^�N*0=�:�>�&?; �>�l?�1�6�;�ˋ�q�����Ͻ]�>��>�>{�)?n-?i�]>KB-�%�}��+����>\q >��=�c.]��ʢ=��=8W�>��N?W?"�_��=;={N>og��	�>8n�>�O�>��N>�g>]e��
��ۿ9{��	�P˾1�)��1>��X�3��oY>M �����^ۧ=�D�=�(=�*�>��ŻK�\>/�[>��>x�`>��>�+�=�%�<NI{<53ؽ�<+<��>���={v��e7����y��Gp��P���������N<��,?	��>)'�ܸ�����j⹾G���9?�^�>!��>�3?<��>G$��_��Yn�i�I=�?�=h?���>�f��Ԣ=Ƅ�������>��?ş+��q�=:��v �Ǘ��Ks?!�'?#N�>[{�����Ш�w�%�ǵ?�m��%𽖁�?�T�?c���10*�΄����M���D��G>z$����������:�̾ѩ��
��mF�����>��>��?D�=ҁ�����'Y����;�译��w���y�>C]#>�:��s�ѽ)nԾi����5�޿?=N��q{>�qD޽��.?���>�9�>[�'?�GH?�c�>#��>|�u?7����?$U>�c���3���ӫ>C�0>���8�*�|���Y|���r����=�J�w=S�p>���=hP��j=���=��9+�F�'�W=��=/�?�$6>=�I�= A�=�2f>Lb�>���>�T!��7T=�.�1 R�䦾�IE��
�<Т��P�Z��ĕ�5#>���>�[E?Bl%>�헽���f�ƾ��ݾj��>�?]?���>Eg��P�ܽYo˾�Q���zD>Щ�ǜU�p����W�3_��X�=��<��>��>��_>��?~�4?c?�Cƽ�A���h��5�c�=O6]���>���>�I�<�Cܾ�.#�Ӻi��dg��7/�]���C q��h�=V�>�\�=��>H��=}��=jq�=z���]����;�$�l�>E<�>��?��B>��=�}u�8���K�L?��My����|�վ���֯�>"�>���_-0?�����u��ģ��zI�,HQ>�?���?�V?-HW�Ϩ��nGG>��};�^�T�w���Z�:�>>P?O>�y�IFw���۽+±�4h>�$>h`Ƚq(��'c�_'˽��¿EVB�<�׼�^���e*�Vy���T��!��݆���"��ã���]����A�L�B��>��(Z��+!Ⱦ^Z���ѕ?�v�?���>��==��9:�����~��=x#�� P��������}����{ܾKe�R���B?�
�'��P��ܩ�>IK̾�O���l��XL�z����>	�y>
�.�U:���eL�R�=�/?�D�>�&��X�8�h�,�3���W?'�_?*�T�������T.>'.?��>V*�>��%=���d��>��f?�b�?aKL>a���򴘿�v)��М?�B�?j_?��%������*A����?���>�<�>ξ����~ѻޘ^?���?�>?��+��	��{i�t��=+�>�L��#�>g�>��>�~���(]�I���a����=u��L�����џѾ�*]����>HL'>.��>��ܾW	���>j��>5N�"H�����V�<��?ʎ�%�>ػe>�q>t�(��댿����� ��M?Vp�?�R?s8?�|�����8S���ґ=���> ��>֯�=��K��>�s�>�s辗�q�K����?��?.p�?��Y?h�l�,ؿ<�=]��7����q�=����bl>Ni��>"�>�?���=��_�=��E>�H*>��V>��="�>`�>�
���+������2��l�1�����׾����Ⱦ;S��Q���ŗ�	���.*���?�a�n<a�j��o4�CzQ�)?f���=>��?a��>F^[>����،�ǕB�A�¾�������4��@���~z��`*�f&�=�!�=j%~���;�z��?��>��P�
�d>,��>�;���=c�p>��>��>�-/<Q�l�	_>>U_�>?�>D��>�,>�z~>FI�=Tᄿ#����5���B�e@�;��C?��A�/j��d@.�Nݾ x��~=u>�N?�L>�&�-Ҕ��t��M�>iW.��?P������k!�̠�>3k�>�֯=Q˹���z�>l��yw�=D"�>�$>�,O�Q������e�=��>P����ߨ=�k�=�?�O?H?���=5�>��S>�/\>��<���=/r)>r:^>Zr?��7?��;?��>��>��u�k$>(/>**A�`���5��F��<��/� &�=HL�;/ό<k�<��<`2W>_�>���;����>W�>��"?;�>]�{>�Ž�]��ꀿ ���s�o��\���	?��>��>�	?�?�ƛ>�q��Nn�=~�o���>�>�]?� Od�?��5b>��~>�#!?ٮ?@�E>��&�����:\=�l�>��K>jk?�s@>���=_�=K��ӿ"��2Ȭ���Ӿ�x��ܲ>jg���*}=�? ]S��B$�������=��/>~��>�F���`>��'>=��>�$.>A>�E(>o	F�!'H=C˽m8���?+�ե<��T=b������}=��>�����v�=�o=Z�?��?���-����K��ƒ:�g�۾�t�>Kz�>_V�>>N	?��>U�龾�S��4˾�F���>$�L?�?��,��6�>�W,�Q�;=Ϝ>\�>l��\�[�b��=)�'�k>"�,?��8?%4�>�<E/T��뢿�<�G�>a����v��K�?f�g?������wD��'n���-���z>�	޾%]ؾ ������4����бھ��R�3�=~� ?܁?�^��J=[ݾ튃�\�M�~⸾�a0�&�>�2�>��> ��=R���s�ܾ� ���ݬ�<�<���>ޒ�
K?���>Nt���~:?�j?�C��E�>�7?"&�=��>��=����^�=b�.?��4�Gb���p���>#pٽG�����=f��=J;>`�>�SZ=����F�=ф8=e�&�[m�"b�2G~=�L3=ms(��=��<w�C>��>?`R�9]�=�����y�� ��8K>�|:>z����>�1�G�rS��Fՙ>Ђ?���>�B�fd��
��]�&>��?¬�>�1>�7����=���=DM��<4	>b�h�t������J��!y齿�`<�ذ>x�L>qR��/l>�4{?�D=?��?�κ�k�$���y�9Z*���4�Y6z����>Z�>Z;�=׌¾*�kl���^��U,�W׼j�B��ݣ<K��=Q�,>�?>2��=U7	>%�`=��[�i ����\�񶯼��>� �>�h?��_>	�W=54�����,?P�v�[\���:N��*ƾɾ̽�|>GW>�YW��'?D�S�#g��;���DHC�q8�>-��?�f�?�DE?�O���2="Ъ>����5𠽇s��߳=	F �����h1>��
>����(�7�`U>�{�=`��>�M<�ܾ���w=}���JD��)=<ks��;髾�f��	ɾ��	��9��|QͽW��b&���`���]��L���-ý�Nt�����I��A�?x��?���>�>P�9��G�t����:7��&־��ܼ������������6���$�������t߾�
��1�>I�Ⱦ23]����0!���\j=�h�>�>�%�nha���D��)�>)Q?e��>�U����k�HO���}#��*\?�Xk?|�W���K���̽�o>� G?�v"?n�&?ǳL=U�Ͼ��>W�a?��e?�5>�[���Į��|g<��?�:�?'�c?�;�zn�[�½k��>V?]�??נ�>'̓��A�'��>�<h?�ɑ?�p?�뀿�p��j>?8Z�׬���w|�!��>��>�}�=u7;� ݾ��W��R��*fԽ2�"�G~��ta]�	���*�t뮽��>���>m	���|����>�š����&�������F4ƽ�0�>8z��p�T� ���ϼ"�C�����Kq�`�ѽT1R?E­?'�+?�FT?ODȾ��'��Cw��&����>�9�>�r>*�%�[�!>zg�=W�'�%�b��X����P?;�?�%�?��D?��H��ϿTॿ�S�˧���6>d�T>�ӷ>�M�@2�=�陽y�4<�=�]>�1�>�h>��v>��">l(h>�C�=�:��x�&�U���Y���:����=i��w�߭�SQ���龓[��ک�����x�O��� gν��;"I����>z�>~&�>e��>��>+��>g�	���߾�j8�=�߾��D���"��p�ܽ۞���Jɾ˾8�澶�ڼ=����>Z���0�X�>hz��O��>�h�>!R=��>\F�=��R>v�>,�=��=�6>��s>ju>�Ϸ>��=Օ��.���q���P=���=�=?2���R1><?u@�C61�W�쾕��>Q?�8�>�Kھs���2G�6*�>�\*�NӰ���c�CF��i�>�G>8�=��ݼ�
½=����;<�я>���>O�>w�!�F4Z�>�}�q�]>��>]Y羪e�=��#>�{?'~�?)?1��=d��>W�K>��>/�<x�->n^�>�>��?��?�?f��>G_>����-�>�/>������Ἔ�� �"=w�n�̗U�Fv�=���=�3=>�w8��W�g_���ɻwK��<s=[`?^� ?X��>� ?�w��{�[�l�L��9�>୭=��>o�>�>��B?D�?j.>=ͼe�H>앑��C�2�?Le�h.��S�v�������	>��@>���?_S?���=��`������=��$�>&�?>RI?��9?�?�D����e*�A�)�}'�u�`����=B��>��P��`�Sa���A޽R�={ѐ>#�>�'>�R�>�c>V��>=��=B��>���>��]>(3>����]H��$̽�}�;�[I<��*=�8�ִ��<2<�12�}��c�ǼsfX����A�	�l�1?A*?�_����7=N"$�]붾U*'?�F�>�`B?!��>&Q�>�꽾U1��$�>k��S�B?���?�ck>�r���U>.��={��=�U�>�$�>}�>`Ծ�t�=c���㌽=]��>i��>è�>"��F%���w���9�>�x����Dd�?�Q?>����V��.�9��
���ٽ�~>��D�cr��;� ���7�=�)�K�(��ܙ�5x�=�ؼ>B0�?�W:��:> �9+c���䑿M���$6�<[M=]#?+�>�2��Z-0��}L���о"J~�Aa�>ц>��6>�7�>x�&?��3?'�?�?R^P?�U���-?��C=U� ?3�?d�1?t�?F�>��{>�:|>t�>ڳ!�y+�r�U��,=��P�L�=��a>Y~i>�Q7<2F=d�?Q�<�C���.>��=���=�M�=�G�<v��=j��>�?Q?��B�4���SD�S͔;b�=��=u>�Zx>�@��"�"�`r޼q��>�T>?�P�>Q�>%��}l����!�B>�o?�FZ?6�!?��}=���>+e-�&�ڿw�Hj`>�>$P�����,@��>����7�V>`E���^�>�M�?�6R?�=?��Z>6�@��ˊ�[\M��Թ=]Nm�߷$?�G?�Gj>�T�\Vr�%���Fl�.����L>����x����p>�>��<r�=sb~><��=b蟾^�!��.j�uEܽ	N�>���>"��>N�2<D�>�ľ�G¾��F?�ZV�E\i��%�i(C��q�=#Ш>�2X>VzL�i��>*���/����)����پ!<?���?�˹?�^?��->�~V=��I=�ӈ��m:<=+�=Kt�= 'ƻ��@��=��>Ւ=�Pþ�t��3E>A��><�=%��u� �CB>s1���^J�]G?��c_��Ez����1����s�(e��;(��Κ���'�HI���;����)�D�󡭾��g=���΅?��?s�U>��%������7���=r��D��ξ��M?ƾ^�ʾ��ƾZS.���A�&^4�UD��q#�>05\��4�� �|�Q�(���l8�>>�?.?�\��� �����{C=pE>�p�<"꾇މ�-��B����V?��9?X�5񾠷Ͻ]>��?��>/>-푾|[ �*`�>��2?��.?uY�6��o���N�t��ں?v[�?��@?�CM�%�A�{������[?3�	?NO�>6找�ž5+�US
?7,9?��>ȉ�,q��"�����>E!X?RN���a>Ǣ�>���>Ȥ�\���'�!��甾����=>�P��9���q�(�C���=,�>Ly>S�4������>�š����&�������F4ƽ�0�>8z��p�T� ���ϼ"�C�����Kq�`�ѽT1R?E­?'�+?�FT?ODȾ��'��Cw��&����>�9�>�r>*�%�[�!>zg�=W�'�%�b��X����P?;�?�%�?��D?��H��ϿTॿ�S�˧���6>d�T>�ӷ>�M�@2�=�陽y�4<�=�]>�1�>�h>��v>��">l(h>�C�=�:��x�&�U���Y���:����=i��w�߭�SQ���龓[��ک�����x�O��� gν��;"I����>z�>~&�>e��>��>+��>g�	���߾�j8�=�߾��D���"��p�ܽ۞���Jɾ˾8�澶�ڼ=����>Z���0�X�>hz��O��>�h�>!R=��>\F�=��R>v�>,�=��=�6>��s>ju>�Ϸ>��=Օ��.���q���P=���=�=?2���R1><?u@�C61�W�쾕��>Q?�8�>�Kھs���2G�6*�>�\*�NӰ���c�CF��i�>�G>8�=��ݼ�
½=����;<�я>���>O�>w�!�F4Z�>�}�q�]>��>]Y羪e�=��#>�{?'~�?)?1��=d��>W�K>��>/�<x�->n^�>�>��?��?�?f��>G_>����-�>�/>������Ἔ�� �"=w�n�̗U�Fv�=���=�3=>�w8��W�g_���ɻwK��<s=[`?^� ?X��>� ?�w��{�[�l�L��9�>୭=��>o�>�>��B?D�?j.>=ͼe�H>앑��C�2�?Le�h.��S�v�������	>��@>���?_S?���=��`������=��$�>&�?>RI?��9?�?�D����e*�A�)�}'�u�`����=B��>��P��`�Sa���A޽R�={ѐ>#�>�'>�R�>�c>V��>=��=B��>���>��]>(3>����]H��$̽�}�;�[I<��*=�8�ִ��<2<�12�}��c�ǼsfX����A�	�l�1?A*?�_����7=N"$�]붾U*'?�F�>�`B?!��>&Q�>�꽾U1��$�>k��S�B?���?�ck>�r���U>.��={��=�U�>�$�>}�>`Ծ�t�=c���㌽=]��>i��>è�>"��F%���w���9�>�x����Dd�?�Q?>����V��.�9��
���ٽ�~>��D�cr��;� ���7�=�)�K�(��ܙ�5x�=�ؼ>B0�?�W:��:> �9+c���䑿M���$6�<[M=]#?+�>�2��Z-0��}L���о"J~�Aa�>ц>��6>�7�>x�&?��3?'�?�?R^P?�U���-?��C=U� ?3�?d�1?t�?F�>��{>�:|>t�>ڳ!�y+�r�U��,=��P�L�=��a>Y~i>�Q7<2F=d�?Q�<�C���.>��=���=�M�=�G�<v��=j��>�?Q?��B�4���SD�S͔;b�=��=u>�Zx>�@��"�"�`r޼q��>�T>?�P�>Q�>%��}l����!�B>�o?�FZ?6�!?��}=���>+e-�&�ڿw�Hj`>�>$P�����,@��>����7�V>`E���^�>�M�?�6R?�=?��Z>6�@��ˊ�[\M��Թ=]Nm�߷$?�G?�Gj>�T�\Vr�%���Fl�.����L>����x����p>�>��<r�=sb~><��=b蟾^�!��.j�uEܽ	N�>���>"��>N�2<D�>�ľ�G¾��F?�ZV�E\i��%�i(C��q�=#Ш>�2X>VzL�i��>*���/����)����پ!<?���?�˹?�^?��->�~V=��I=�ӈ��m:<=+�=Kt�= 'ƻ��@��=��>Ւ=�Pþ�t��3E>A��><�=%��u� �CB>s1���^J�]G?��c_��Ez����1����s�(e��;(��Κ���'�HI���;����)�D�󡭾��g=���΅?��?s�U>��%������7���=r��D��ξ��M?ƾ^�ʾ��ƾZS.���A�&^4�UD��q#�>05\��4�� �|�Q�(���l8�>>�?.?�\��� �����{C=pE>�p�<"꾇މ�-��B����V?��9?X�5񾠷Ͻ]>��?��>/>-푾|[ �*`�>��2?��.?uY�6��o���N�t��ں?v[�?��@?�CM�%�A�{������[?3�	?NO�>6找�ž5+�US
?7,9?��>ȉ�,q��"�����>E!X?RN���a>Ǣ�>���>Ȥ�\���'�!��甾����=>�P��9���q�(�C���=,�>Ly>S�4������>�š����&�������F4ƽ�0�>8z��p�T� ���ϼ"�C�����Kq�`�ѽT1R?E­?'�+?�FT?ODȾ��'��Cw��&����>�9�>�r>*�%�[�!>zg�=W�'�%�b��X����P?;�?�%�?��D?��H��ϿTॿ�S�˧���6>d�T>�ӷ>�M�@2�=�陽y�4<�=�]>�1�>�h>��v>��">l(h>�C�=�:��x�&�U���Y���:����=i��w�߭�SQ���龓[��ک�����x�O��� gν��;"I����>z�>~&�>e��>��>+��>g�	���߾�j8�=�߾��D���"��p�ܽ۞���Jɾ˾8�澶�ڼ=����>Z���0�X�>hz��O��>�h�>!R=��>\F�=��R>v�>,�=��=�6>��s>ju>�Ϸ>��=Օ��.���q���P=���=�=?2���R1><?u@�C61�W�쾕��>Q?�8�>�Kھs���2G�6*�>�\*�NӰ���c�CF��i�>�G>8�=��ݼ�
½=����;<�я>���>O�>w�!�F4Z�>�}�q�]>��>]Y羪e�=��#>�{?'~�?)?1��=d��>W�K>��>/�<x�->n^�>�>��?��?�?f��>G_>����-�>�/>������Ἔ�� �"=w�n�̗U�Fv�=���=�3=>�w8��W�g_���ɻwK��<s=[`?^� ?X��>� ?�w��{�[�l�L��9�>୭=��>o�>�>��B?D�?j.>=ͼe�H>앑��C�2�?Le�h.��S�v�������	>��@>���?_S?���=��`������=��$�>&�?>RI?��9?�?�D����e*�A�)�}'�u�`����=B��>��P��`�Sa���A޽R�={ѐ>#�>�'>�R�>�c>V��>=��=B��>���>��]>(3>����]H��$̽�}�;�[I<��*=�8�ִ��<2<�12�}��c�ǼsfX����A�	�l�1?A*?�_����7=N"$�]붾U*'?�F�>�`B?!��>&Q�>�꽾U1��$�>k��S�B?���?�ck>�r���U>.��={��=�U�>�$�>}�>`Ծ�t�=c���㌽=]��>i��>è�>"��F%���w���9�>�x����Dd�?�Q?>����V��.�9��
���ٽ�~>��D�cr��;� ���7�=�)�K�(��ܙ�5x�=�ؼ>B0�?�W:��:> �9+c���䑿M���$6�<[M=]#?+�>�2��Z-0��}L���о"J~�Aa�>ц>��6>�7�>x�&?��3?'�?�?R^P?�U���-?��C=U� ?3�?d�1?t�?F�>��{>�:|>t�>ڳ!�y+�r�U��,=��P�L�=��a>Y~i>�Q7<2F=d�?Q�<�C���.>��=���=�M�=�G�<v��=j��>�?Q?��B�4���SD�S͔;b�=��=u>�Zx>�@��"�"�`r޼q��>�T>?�P�>Q�>%��}l����!�B>�o?�FZ?6�!?��}=���>+e-�&�ڿw�Hj`>�>$P�����,@��>����7�V>`E���^�>�M�?�6R?�=?��Z>6�@��ˊ�[\M��Թ=]Nm�߷$?�G?�Gj>�T�\Vr�%���Fl�.����L>����x����p>�>��<r�=sb~><��=b蟾^�!��.j�uEܽ	N�>���>"��>N�2<D�>�ľ�G¾��F?�ZV�E\i��%�i(C��q�=#Ш>�2X>VzL�i��>*���/����)����پ!<?���?�˹?�^?��->�~V=��I=�ӈ��m:<=+�=Kt�= 'ƻ��@��=��>Ւ=�Pþ�t��3E>A��><�=%��u� �CB>s1���^J�]G?��c_��Ez����1����s�(e��;(��Κ���'�HI���;����)�D�󡭾��g=���΅?��?s�U>��%������7���=r��D��ξ��M?ƾ^�ʾ��ƾZS.���A�&^4�UD��q#�>05\��4�� �|�Q�(���l8�>>�?.?�\��� �����{C=pE>�p�<"꾇މ�-��B����V?��9?X�5񾠷Ͻ]>��?��>/>-푾|[ �*`�>��2?��.?uY�6��o���N�t��ں?v[�?��@?�CM�%�A�{������[?3�	?NO�>6找�ž5+�US
?7,9?��>ȉ�,q��"�����>E!X?RN���a>Ǣ�>���>Ȥ�\���'�!��甾����=>�P��9���q�(�C���=,�>Ly>S�4���ܢ�>���'���j���+�1l*�P<M��>ߕ~�G��=�a�����@�G��L��]�d�b��;M?�۫?��J?��3?ٷ����f����
�=�U�>K�>��5�G(K���j>�q�>�B¾6.R�)*��1�>���?���?Q�a?�`�}�ƿ����t�'uԾ��>M7>�}M>y�[���=_z�Zh=���<��n>�R�>���>��r>��n>;:6>ɡ�>/&��48*������Ɛ�x�3�h�ؾv���'��׾&����:Ҿ1���bѩ�_w\�����]���ђǽz����U�����<��?4v�>k�F>��>+�=1	徆�+�/ꕾ��⾕w'��]
�1�
��l�fCi��#����+�8#׾��f�վ��>��<G�=5�>��T���O>��1>e(6>�]}=0 =fg>3��>}�]>XG�>m>� �>��f>9y}>n�=�-��d���9��T�Qw<<Z�D?��^��`��hn2�,�o���8D�>V?r/T>2&�n&��n�x����>�E���b�}�ӽWD���>D��>�{�=�2����Hw�MB꽑z�=q��>z=>��X���D�+�=,�>8�����J=�=�{?��u?��3?3����=�ȑ>��@>wh>� >n��=	7�>�<?�t=? 6?F@�>O"�=A�����[>���=]L]��*`<\0W�>�>�#E��Z�~��=���=˦=�E+>r�=7-估��P�����>a�?(66?�.|>��?O���l���I�t='F^��U>��>��=>�$?
�#?!��>ԙ!>�ɽP������{�>!k>�.����{�0����S��%�>q�?�~9?�w>�F>��m*=c��=ҁ�>�>�>�3??@?�5�>�4&�����翅L��;%��j��?Y=��Z<����S��R��=n�ҿ�	>��>��>�~>\3o>�y">��>���>0�=>�>>��,� Ճ<�N(��1��"5O�Y����yM����8�M�Ž0v��!|�0D���c�yb=O�?��?�9��~,��FV����`Z��,�>�'�>���>J��>V�=��
��2T��i-�#�/����>w�W?>�>��y��A�=�&�<4Y=w?�l�>��L>�X2�᥇�i㮾5��=&��># 6?��e>"�c{Z�_Ǆ�t����u> Nѻ�78�J��?�gw?�����Q�c.�D�Ͼ�
�^�R�ļ4>�w��;����Ǿ>5��K��������G�@>	��>x��?� ��W�>i+N�C����RV����
��>ĝ�<v�?6�='�l�}���[J��Ⱦ
���<�<�>g�>�ޟ>���>� ?�"o?`�??�:���m>(�j���?��1?��/?t_K?}�?�>;aܼ������:�p=s���=�=#au=h/M>w�=7���,�����`��Ҋ:<�=�v�=;�>>Հ�=^t�����=�?�@1?�����<��=�R��D�x>��>��>o�7>Iw�����yN>U?��?2w�>W��=�y����ݾf)��I�=��?ξ	?Q�?m��=9�>�[��Mk%�Ϸ�=�z-><�">�闾^l�7���Zq0�u�=>/�>�o>�w~>�H�?#�>�?���>�O�ƻ��"�ٲ�>1� L�>3`�>��>(�����槓�n9���j<���">SxҽX��<���=����֞�>L�$>�>(u������̶ּ<��R�;�W�>���>If?���=C#�<�n���
���-?�J{�bj�r5�Ȇ\��=����>��x>f�>��>?�6(��pP�;���r�v�ZK?�ѽ?Ƃ�?�Ɣ?�����C���lk>�&>֟T>�Q�;݋	9<w{<�x �Q{/>���=��ʽ�)���=�>>*p�>��@��n����۾���/Ŀ73��B<>.�ؾ:���� ������^ھ�Kɾ�-� �����~���ҽ].��~Ο��ȣ�D򩾞�e����?Jx�?Go>�w�<��*����%�ؾ�T�=��\�@���渾8E�_g���g徭�J�=�J65���%��t�����>YY����T�}��)��-���#C>QO0?��¾~������V=z!>���<M�����w�����$�V?�Q:?pq쾧k����s$>�g?�d�>��)>C���޽�4�>`A6?�H.?Ԑ�{������4�z�G�?&n�?�hD?ap+�*:��|꾾[���:?�	?���>���0��$I��a
?�;?,�>f� �A@�����>�hG?�9��mh>!3�>�?�>��������ɽ?����^Ag>.Hs=������@��S4�uq�=�X�>j>��j���;ܢ�>���'���j���+�1l*�P<M��>ߕ~�G��=�a�����@�G��L��]�d�b��;M?�۫?��J?��3?ٷ����f����
�=�U�>K�>��5�G(K���j>�q�>�B¾6.R�)*��1�>���?���?Q�a?�`�}�ƿ����t�'uԾ��>M7>�}M>y�[���=_z�Zh=���<��n>�R�>���>��r>��n>;:6>ɡ�>/&��48*������Ɛ�x�3�h�ؾv���'��׾&����:Ҿ1���bѩ�_w\�����]���ђǽz����U�����<��?4v�>k�F>��>+�=1	徆�+�/ꕾ��⾕w'��]
�1�
��l�fCi��#����+�8#׾��f�վ��>��<G�=5�>��T���O>��1>e(6>�]}=0 =fg>3��>}�]>XG�>m>� �>��f>9y}>n�=�-��d���9��T�Qw<<Z�D?��^��`��hn2�,�o���8D�>V?r/T>2&�n&��n�x����>�E���b�}�ӽWD���>D��>�{�=�2����Hw�MB꽑z�=q��>z=>��X���D�+�=,�>8�����J=�=�{?��u?��3?3����=�ȑ>��@>wh>� >n��=	7�>�<?�t=? 6?F@�>O"�=A�����[>���=]L]��*`<\0W�>�>�#E��Z�~��=���=˦=�E+>r�=7-估��P�����>a�?(66?�.|>��?O���l���I�t='F^��U>��>��=>�$?
�#?!��>ԙ!>�ɽP������{�>!k>�.����{�0����S��%�>q�?�~9?�w>�F>��m*=c��=ҁ�>�>�>�3??@?�5�>�4&�����翅L��;%��j��?Y=��Z<����S��R��=n�ҿ�	>��>��>�~>\3o>�y">��>���>0�=>�>>��,� Ճ<�N(��1��"5O�Y����yM����8�M�Ž0v��!|�0D���c�yb=O�?��?�9��~,��FV����`Z��,�>�'�>���>J��>V�=��
��2T��i-�#�/����>w�W?>�>��y��A�=�&�<4Y=w?�l�>��L>�X2�᥇�i㮾5��=&��># 6?��e>"�c{Z�_Ǆ�t����u> Nѻ�78�J��?�gw?�����Q�c.�D�Ͼ�
�^�R�ļ4>�w��;����Ǿ>5��K��������G�@>	��>x��?� ��W�>i+N�C����RV����
��>ĝ�<v�?6�='�l�}���[J��Ⱦ
���<�<�>g�>�ޟ>���>� ?�"o?`�??�:���m>(�j���?��1?��/?t_K?}�?�>;aܼ������:�p=s���=�=#au=h/M>w�=7���,�����`��Ҋ:<�=�v�=;�>>Հ�=^t�����=�?�@1?�����<��=�R��D�x>��>��>o�7>Iw�����yN>U?��?2w�>W��=�y����ݾf)��I�=��?ξ	?Q�?m��=9�>�[��Mk%�Ϸ�=�z-><�">�闾^l�7���Zq0�u�=>/�>�o>�w~>�H�?#�>�?���>�O�ƻ��"�ٲ�>1� L�>3`�>��>(�����槓�n9���j<���">SxҽX��<���=����֞�>L�$>�>(u������̶ּ<��R�;�W�>���>If?���=C#�<�n���
���-?�J{�bj�r5�Ȇ\��=����>��x>f�>��>?�6(��pP�;���r�v�ZK?�ѽ?Ƃ�?�Ɣ?�����C���lk>�&>֟T>�Q�;݋	9<w{<�x �Q{/>���=��ʽ�)���=�>>*p�>��@��n����۾���/Ŀ73��B<>.�ؾ:���� ������^ھ�Kɾ�-� �����~���ҽ].��~Ο��ȣ�D򩾞�e����?Jx�?Go>�w�<��*����%�ؾ�T�=��\�@���渾8E�_g���g徭�J�=�J65���%��t�����>YY����T�}��)��-���#C>QO0?��¾~������V=z!>���<M�����w�����$�V?�Q:?pq쾧k����s$>�g?�d�>��)>C���޽�4�>`A6?�H.?Ԑ�{������4�z�G�?&n�?�hD?ap+�*:��|꾾[���:?�	?���>���0��$I��a
?�;?,�>f� �A@�����>�hG?�9��mh>!3�>�?�>��������ɽ?����^Ag>.Hs=������@��S4�uq�=�X�>j>��j���;cN#?P��t3��:�.�*��m��>~|�>T��>w?���>��>���U��i�����[y�=�d?�!�?/r?L#!?����쁾��)>�f>�_?��>f8���*�����>�'�>2C�癆��@��?2�?<}@�G?}ⅿb�̿�6���%Ⱦ2�Ծ�:==��='��=�1H�n��=r)�=�@ν��!<c-b>sƯ>�>�j>0R>�!>d��='Å�(X#�ʫ��I:��F����]��(�v�վj��%A�f��!�ξ�����Џ�n�ٽ��K�tU�>G�pڬ<�����(9;�?��>��?��=�%!>�.[���������۰��u���þ}Ѿ�H���Un��	���1��Fz��	���b־��>�����=G�>iY��>wH�>;q#>���>�p����O�'z�=���<��/>`/>�u�>A�3>��>IJ>� ���`p�K	4�����,����&R?����ھ�rJ�]/̾٤��*��>�"?z~M>,e3�����B��hK�>m	ռO�����+�f**=kC�>��>�s�=��=�" =������<}=�->��>ג!=��8�~�e��ia=�8�>��׾Ú
>�@Y>lo/?�^g?�.?�=I[�>��^>�u�>@*�=j�D>��,>�S{>Q6	?��!?mj%?�g�>xl�=me�┼<5�=
O�E���ڽ.a�0��N��<��U<�K�=Z�T=�,I���=�`�=T�P�c3;�^=Ң?'�Y?���>�;�>�Du�2�%��j�D�<V��>+;����>��?p�>�)?�s�>G���ᚾ9�=��<3��S?���>G~��T�t��բ��#�����>=�r?��f?:҉=x!ʾ��W��n�>9�!?g"?E�G?�bd>�̱:��d��ؿP��:*�3�z��c��5�=����������>�\����Ȼ�JI>i��>�Jx>��E@�����=��>ǎ>L�]=�>!��=��6>� �U�=d�=#x�Ȣ<(ț;"�T;�i=���}�;n�l9kw����Z��w�\n ?�P?B��>���>����Ϛ(��𙾶��>�do��'�> #�>Fә�H�V��lP�8�o���i��?�V?w��>�7���e�9��Q5�z��>��Q>3�H��=2��5Ģ��g�=tD+?Y06?ڪ�=�����_�芋���$����>�>������?ǞG?�O��I���V��E.�׸���4>�ޔ=4������.�2� .����iҾ(7f���=���>�?j�eC>*OC��掿 d���< �=(�>G�?xr����]�[�
��N�����=��>~��=iZ8�^>n�?��?2�?�g�>A��>+p�=߰>此<}��>P?K�>!�?��A?kؑ=����2н'���\�������4�=��x;B��=fZ>��=�#�8������=��^=,/�<���0�ɽ���=l�=B��=ہ>-��>��?�e?��ž�>W"F>D��DW<>�??Zx	?E܃�/���V�H>G/S>�{C?GM?�Y~>h�k�~�ܾX 8��2�(ܽw�*?*�E?�w?Tĸ<��=�~��gt����>O7�>��~=?�-���˾��5��>��>��>�r�>rY�>ȏh?�+s?��%?�9�cѾ������Ҿտ���Ǿ��>`�>~{=J\ھ@�9�7-���~j��G��<�A�?���;B [>���<��8>�S�>���=�rH���?>��5U���|>	P>�7?]�-?��=yԼ6����Sq?v����D�"���ܾ*ȿ>u�?��ɾU
;�V?"�%�虲�j][�4	��^{<7i�?!e�?P�q?��>�|����>��>r�W>�?=cf�ꊥ�_zB��>����y �r8Y���:���y>��>�>��6x��q7�����pq����[��;�z*;�r{�߻��$�׾0@��VM��*��qˬ����<�lp=2=�i=8e�/žѶ�lj���h?��?ȱ�=����4\&�:C��*)辤��<_�������x��9F=�~���堾m�ݾ+����"+7�:�T��>�*$�S���k,r��,J���y����>2v;?cܾ�u�������y���>��>�)���Pk�+�p�X&>R�w?*��?i�5���O����������H?��F?��>�$��:ǽ�A>b��>�τ?����P,���}Y��yY����?���?C�??y�N�~CA�Q��D�h�?3�?VL�>#���?:̾V��G�
?��9?)�>83�,8��'&����>�n[?�LN�׶a>���>�ח>��d���[,�gǒ����m�9>�X廞��s�h�c�>��Ȩ=��>�4x>R�\��箾���>���H��?�R����=����>&�K>Sj�سs>��>Nk����ҏ��玿��=���?�-�?��?:�x?��&�IK�%4�����Y?�a?o�=�����?5?�4����#p���?���?���?Z�>?xK��xտN��.s��-���C��=�.�����=1%��Hy�=M;<kߟ��%%=�>���>+�>A�">>�=���=|l9=�n��D_0�+����M���O�p�5�x��UAA�d��e���wj��Z�J)z��מ��3����M��sC��)\�%L!>��?��>4b!>�v/<���=ǭ�
\��ZQ�K�+��w=��~"����ֻ���4���$�!�w��_ǽ�ӷ�#✾t,?��8>��<�V>K�<��I=�3�>�j�=���>Y�׼�/=�'J1>�D���V>X�W>癶>��=pdz>�2�=%G���g�� �8�Q�O��E�;��@? ^��4����5���߾!n��N�>E�?�T>@'��d����w�'L�>�&:�F�\�sν�&�+b�>���>���=c�.;���ѓw�&��̚�=�>i�>���ȍ�����EC�=s��>d�Ǿ2��=�"{>��%?+�r?��2?%�=9x�>.+\>��>O��=^�?>��U>��>�~?![6?�2?��>��=8`Q�w��<��<�j9�0iV�DE�� ��k�.�&|�<U��s=��I=��<9�(=�=���cp�<���<�K�>vTD?[�>%�>h*���$�3W4�����x>�7����>�<?�1?�(
?�ֽ>�=�)+��BӾ�ݾ�o�>(�>]_f���X���н�>렲>*�O? ?
�������4�!=� >Hf�>��>(�?P��>�[>��+�����ؿL.0�?q8�_r��`���~�����;H:=��>�>s�y=����<�>�]m>�H�<[?>��]<&��=���>���>�= >>mn��T�K���轉`%��&y�J�=��:>�����=z�ٽ" �MY����	�}i �b9�=�?c�?:K�>-�>!�ܾ%\��Ll���U>��>�g�>�9?޽ϼ�	F�:�B�|_�`�1����>B3d?��	?�0��@,>O*���҇=>==B>إɽE�=�"��=`�+��/>��>?E�)?4��=�B>����_&q�hW-�
��>o��=3��	 �?Fib?�n�r���B��~?�H���=���D��=-�Q��TN:�ꭷ�%�Ǿ���|�>V�>�r�?3�ȽǦ�>��ľ����qh��h��䔱=���=��?[m>N�Q��ρ��_|��ЊȽu=�E�>A�A>JG?/?�*�>�4W?  ?k4G>ތ�>ɠW?N��=��>�j?��"?�l�>���>.����Jb�t��=Lu�y3��R��TH=�/J��S>�<9>���=��<�:C>m�	>��)��{�<�ʽj�6�=�>0��=$z�=�-�;	�?s@"?�F/���=��潈�ҽ�!T=���=Gv=X7�w����➽��>�?��?�a�>���=�tݾ��2��
,>��?��?�S�>5!=Z鞼=�,˞��{%>%g3>��=o�a��F��
�>���m,I>A��>��>y}{>`u?ۭ>?`pZ?T�b>����J}������^�>Oy��>���>��=l9��{-3�deT��y��C��-��T�x�=SXH=|͓��^t>��/>��\=��=�޺\̃�[����H>d��>�C�>D�?��#>�&���t��;T���4k?;���c�&� ���뾿F?Ć.?�{��ы�Y6f?��%�Ì���i�mYU��G?4L�?���?*�6?��=g�,�>$��>���=a92<�s��u0ʾR�=�̅>-�c�Dy
�&�?�<m�N��>R�?�8��������;�I��mN>���j��̾Μ����p}���Y��Mo������w}��-
�n����C%�����u�Ӿc�;����_?�9�?-�{>�7A<;�����Ux��?�����;���(��=������=�d��o���⾥3־���+,"��l׾u0�>ɥ���,6h��俾��=ܴ�>�D?�	;0�3_-�h��>���>Q��>����������>�g?�M0?:龕G.���8���K>�E�>���>s�>Y��5����`>m1?��J?�u�=P����ڇ����<`Ȼ?��?��G?P��`�'���i>.�?a% ?�/E?n8��ǂ<��h�)FB?I*�?:�2?�Z߾D���d��??F?iv?����">2��=N�>�E:�>ʅ�!1��i�Ҽ��+��}�<u�q=��ӽ=���16R��R�<�+<>�>�p��:A� �>�����\����G�
�R���4�5�=}DJ?�  ���>;ݵ��:k��@쾧���|�9����<�~h?iݜ?�da?��q?�����Q�����bn�ҏ�>�w?��5�V�>x�2?�s>x�����A���>���?)@�?]$!?���Sÿi���u�����k�=�>'8<\�M=ק)��<�=����x�=�l>�;`>���>��>��/>��>{$N>:��=��}���+��Q���]���<�.C2��2�����+o��*ξ �쾲���	ɾBM�;|���	��&�a���*���m=�%\��:>|�"?7b^>G6�>���=�y���ؾ�!R��ӆ�eq �5� ���K�>�Ҿ\K׾��/��I]�%�<�m���*=��Z��3?}>��:��@�>A޽)r�>
�>V�<��e=Ng>�z/=��,>vҽ4�+>؆�>�}�>�^U>^p~>���=�ل��Ā�_�:�<�P��3	<mD?�[�3x���c3��h߾JW����>g	?�_V>{'�����?�x�K��>�m>�7fb��ƽ;���N�>'��>d��=	�ƻ�
$��^x�VM���=��>��>Z��	J����m-�=�:�>��־���=�o>�#&?Hx?��6?8�=�8�>�k>�Պ>=��=��H>h�F>���>q�?�Z;?p1?=�>c��=�[�D�=�(=6�:��I��`��j�ϼ����H_<x->�B \=�e=d</�c=��D=���b;�9�<$�?H]>?���>�%�>�P����w���0�,8�=�=K>�PO�ǥ?��>�#?M??��
>k4C���7pL�cJ��>�"�>��c��m;�#�8�T\�=a��>V�]?�a�>�<����
�j>$<�>�5�>��>�AG?Y+�>��=)_��x��!@ۿ�,e��u)��M�>�P!����RǪ�$���9�����2?�=��=�K�>d]�>��J=�8�=R�d>�Մ>U��>��V>Y~1>�d���n=��=>�4���y�P╽!��=����'�½��H��L�:1'���N��T�Ž��{�>�j5?���>7<z���'�����ɾ��>��>"@�=(�?$F>�{V��c�Ԋd���i�+m�> �V?�`?��=R��Z��i>��>�h�s�(4>zOX��
�>K�$?3�*?g�5=�����<b�*N����w�>5e!=@w����?��O?��(b��� �aB�0�&�0Ep<΍���
z�/�ྈ���s6�{x�gu���S5���=���>7��?��M�w[b>��Qы�_t��H�?=�����=I��>0�=�FZ�[��v/��v������H�=Oj�>��h=� ?$?�l?J�]?�E�>Z~�> #=k?a?��=x�>n�M?�GK?�$?���>¸���ݞ=�1;�z�<>y�sN��έ�=�{��>]�q>��=�!=4}O>��=��w=`+;aF��7C<�w>-K=ນ=�%'>���>Wu
?��$?��ͽۦ�=�>?�eƾE�>-x�>��>�q%�-����{Y=!��>O�?��?,0�>���=pɾ�J��7�W�f>���>O?#�=?�
b=��<���֩9��V�=!o>�S$>J�������}����Ӿ��>��>|I>k�P>��`?,�4?c�$?}v�2į�9�a��� �{�&>�Y��6�?���>�A����Og�x��c����n��#�S��Ij�v�>�^>�>���;� >��0;o�9���?�e�$��x.�`��>�?L�?�S�=��m��q0��H��t?T����r]���/���"�+�%?�7?1h&�*�&��y�?�$�LB��P���s�̯?���?x��?��)? �_>�ν���>]Ag>������>7S�:C)�R�e=�a">����	@*��0g�!7�o.�>��>���� ��8�i��������~J��ȽE5���I^��/S��J�Y�¼����P�4�9z�������6�f��_�[7��l���$�� �y��?���?Jp�>��>�7��	�����>~�'�+9<;�v�A�u���ԝ<��^澩o����k�	��9��a��>3�Y��@����|��(�#�����?>�5/?�`ƾwϴ�]��1�g=�`%>���<	;�$���⯚�l��bW?��9?}Q쾞*���Ὤ�>~�?�s�>O�%>�(��Q5�'�>�84?8�-?�S����:��(���+m�?-�?�??�jO�ԕA��������?F�?�>������̾�5�-?7�9?�Ӽ>��$\���3�1��>Id[?8oN�Pub>���>CV�>��<�����%��>��a-��n�9>��
����Xh��->���=Eˠ>N�x>Y�\�NԮ����>k�	���~�������6��4 ���?Y ?e 3��N�>�Y"?͛��]ؾ+ؑ�`ܨ� ��Po?���?��*?֎A?������]��A�>�k	?"^�>6�r���'�ֹx�-?�]ϾE7������ ?�t�?|}�?"E�?�w{��ֿ����Y��V�}�I<>]GP>�@J>�k~�M
�=MN�=�b�;iH�.�M>�+>��N>�-@>�.�=2>Z�~>D[��X�0�)���*���Q�?��,%�����6���$q����-���Ǿ�O+�y���^jT<n�r�=Xn�J\�;��X'>Y�%?~Y�>���>}B�>"���PC�`��rI���2�����)��4�۾v����7�A����[l��c���sM���پ/k?�,��e��;ϧ�>X��Z.=�6�>�A=�hT>�w">(>�=�RK>��N=���=J��=a�l=8Ι=��>� >�����:i�,,:�����P_�=L3L?U�ӽ�ƾcZ ��	���'��]��>�[?�h>{3��ǚ�K,��Ƭ�>�Ĕ<k/�� lڽ���:�t>5T�>��=`=�=�z�����x�;��(3>��B>�N�<+�\�!�
�^�\>�A�>j�Ⱦ���=�un>�?��p?�S!?��=�>��H>V�V>�W=��=GT)>6$w>��?+!=?��.?��>��=��C�B~U=��=0T���ʼN����C�5N����<S��i��<,]=���;yo9=kW=�ǻ�ht���H=Z�?�y<?�һ>���>vw��*&-�����!�Z25>��0�>�̢>�<�>��E?S�X>;8�7��� "�l�:�;"�>�({>�1����J������=S�>�5?�DG?He>�fPo�<�>�:߽�J?�x0?e�?�?> M=��Y�ey�B�׿����Z���kr<�@-�u�d��j����F��=�~�N��<�O>��=Ժ�>�4�=���<5��=�>`��>)a�>ZB�=`�=��k=.x�=�ƭ�+b�=���x(��(=z�0>�M=�'�=D���\����>�ُ;��M�t?�?)�I=��(>`�q����پ���>WP�>�7�>�H�>V�;�H
��
Q���E�I�Y��;?��K?��>��r�:>���=�\��� �>���>S�E:�K=<6��+&ž0��=E	�>�SA?:0�>��/�
���+���"��G�=��=N����ʙ?�V?� �+^2�p(�1�9������췼ez��I�q��~��
5�<QG�'���澢����'�=�b�>�1�?,ߌ�2>��پ����OF�jG����>j�_>�B ?�r1>��<�ԟ���+����l��P}=���=f�?=��>13?0v?�ʟ?�{?�Ԑ<�E3>:Z?�X��+�>�yY?�9?���>?k?NZH�!���?��}���rLR��.��9
���Y��U�=ޠ>��Z=���=R��=���=�(�<ZZ���μ4�z���"=h��=n:>�C'>�d�=|v?�*?�x�4
>Z���k��T��HS�=�&->랾��Ͼ &��1ľ U#?�%@?��>�)�:�v��H�߽��'�>
�?:SE?���>�Q�=�����پ����!D>��>xd0=F����Y7��:�(�4�)1�>+vh>'Ш>�V_>�҂??J?�(2?�+/����O�d��k���VR=/�Y���>���>Ź>#*�������s�G�X�
3;�A A�xQW�bL;�T�>��ؽ�-�>�ׄ>��~=c��=�/��&� "W;}��=�,�>}��>h��>�{�=�Uݽ�_�Oy�7M?0�Ǿ�'�1\����۹�<�^�>���=(��� ?��}��t���Ռ��X��98>���?	��? }y?G�^>��dV�>V�>(ڭ>޻Q��V~���ž��T��>���/HH�
���ģ;��
?/�!?�8�=�#o �<��=[ĺ���B�ܶ���ʾ�=y�e��o$׾ùM��b���ͻ��Ǿ��L��&��[!�:���^�t�}�%F`�γ�����?�?���=����r�x�n�X�Ԯ��
�a>����K A>څ��a�ܾ�k����<��8��~3�����ա��&�>_�]����}�| K������>o�5?��׾r�<
e��J��� �>6�ڽg�#�^避���/���q?@#l?��,�mm��#o��G�?�
B?(
�>�9龮<�9]�>�?�58?�3߽��R}���I=��?���?�@?KL�(B����y�?�?7��>����ʸ;B��Æ?|�8?���>gg�~L��Z�����>�JZ?��N�x�c>��>M��>J�6k��*$*�瓾��`���:>���^O�x�h��@�CƩ=t��>��x>ڐX�����D>gj�����JH�e'"��-�(�4>,��>���(e�>u��=��ս��ݾJr��Q�L���½@8x?�
�?"v=?';�?��!��uV�e�Y����6?�/F?ǱO>-V�=��?�] ?�@������S��`�?���?5�?�}3?��g�T�п����T���ު�����=Z��=8�G>_�����>�l�= �����;e_>�"�>e>��U>�J>�#7>�>�N��I+�ꁢ�����=��Z�l��Ĕ�\\�y�g�
�!��uپ���ڻؽy����E����Y���*��
��nb��� 2>k�?�E�>���=�v�=u��)���-#��5��5�G�/�����)�݁����>U�
<�'���=�*
�6���\�>��=[�<���>��+�8� >�a>6jn���)>n�v>mSm>�=ZW�;/�N>' > �>�>���>z��=�ɏ�"V���9������=�"v?y�%����������}k����>|G?ξ>�1�;�����z��>��=�����n��=��$>��>���=��Z�j�����"���G<�=��>#_>�þ��~�������+�С�>�p��}�
>�Dk>�G?W�k?<?L	�<�~>H�b>Y�=~e��Q�/>y��=��a>�0?��:?�,?��?�=f�4���,=3H=��[��H�;h경^�.����1�H�=��=�S?=`���<y�d="f����<c:�<�
?�MC?&d>��^>�8����I�lG��6=���>�P��?�?�;?o ?��B<9���I�پ�L��¸��#��>�ө> ���b���%��N�A>VA�>�s?!x?]l���P���>D>>�\?�i?D�?Kp�>���F�x�����ֿj��K���^���n�>'��p"[�[	ռmJ�?"�>H˽gp6�Be>�̂>e~R>�61>��>�&>�9�>�
^>�@�=�>�Ω��x��VQ�c���R�o�<N�_�̻Re���bĽf�н��M��C�L2Y���;�+�>��	?fW>��>�$����l��˾�*�>n�>r;�>?��x���.��6�JrM��\�>��>��]?�$	?˄�`��<_p1=�M(=+�?�\>�2�5s�=�|�=9U徚�?�2?
 �>���>n�������灿md�޴.=ظ�<�t}���?��B?0j����-�H�/'��{ܾ΃B���=�F�uB������S�D����)�UIF�ss�=�g?���?�}پ��ٻ�X�M[���7S��T��	�\>��>O��>y�>��=�Zf���/��� �"ɦ�R��=���>WB�u�$>z�?jXB?�ʘ?؎G?�(|>�����v?��޽�2�>]�I?ɱ�=��?_�>s�B��ؿ=�>�=���=�I��3����w�<C ˽��=�	G>-��=��K=�>м��%=�~��i��?��9w;��=8z�=�F2=�Q�=DX�=1?Ҭ?P�羙g\����b�ݾdr>݊>$�������?R�͛>��?�?��I>Vo�=4��{@�b���+>�h?#2?�0�>�@I�i�
���"�>>�v��>���=���,s�T�ܾѺ����<�>�1{>�ҵ>�>Ɔ�?�<?�G?��=�!��cG�ܐ����=�J�7,�>>�>:ӼJzd��2���m��cY��M���G�W���(fr=%��>�	)��ݓ>��> �L<�;���=�;��J���=�=�>�#�>���>&I>�����y�œ�u�_?F�+�oiV�� �n��4sZ>�b?�Իw�W�טr?��������=�T`��0?���?�ʮ?�&?�������(�@>��=��=�C,>����(r��e+�=��(>�r�����)X��hq�L�>UX?����5�n��¹�ܿ��c�u��=H���i�f�ʾ�Th�|��|����=����������U*��y�L�SR�~Մ�n�;�56R<���?D�?t�> P�}�:��q*�J�¾A��<.��"�p�;a%�}9��0��\ѾѷѾ0^̾����+���>��X���ߝ|���(��ܔ��i=>�/?F^ž?g������j=K�&>�~�<V��ᤋ�Ú�4[
��W?��9?���������L�>��
? �>7�&>:Ē�O��Pё>�I4?�.?�׼^��*)��kP����?/��?�J?!�޽S7R�0���Z����>ڔ?;[?��f�U{ﾹU��?�7I?�%�>��۾|�r�&�4ȟ>��*? �]�p�>1��>qw�>���񯉾c��<�N��9�;���>	U�����\\�;��)�6>J�>f��>G]��$��R��>�*꾪�N�'�H��������Ď<�?��*<>�i>�L>?�(����͉����m�L?���?ÌS?�h8?:����������=d�>���>��=��l�>!��>@k�G|r�����?wG�?��?HVZ?�m�>~ɿ�|���!_�ȇ��w��=�L�=o�=\���$�= �=�ly=�蟻[�=�E�>�Ǌ>NGV>�c>>~9>a4�=8��ہ��9��x ���$_�3]0�����`����LɄ�m��b���:�Ҿ�6=�!�4���ཤ&��k W���O�	�������>�)>��>6�w>��>>b���\%�?*̾���K<�]ھ$�����Gf ��D���H��OlI�����;$���>��)>�4�>A� ?B��hʮ=�#�>��˽�_�>�*=c=0=BOd>��>��>C2�>�o>w�>�����=
���@��+�M�`u�w)#>�r]?	�3����c��̾�#�D��(d?[��>�F�1�������%?X$&��R���� �ES=}?�K?!QZ>[��eH>��-����v�ƱI>��->�aK>�3�<9��U�i��k�>=j;?�09�>_H=�+3?1V?J��?a�>?�<�Y�>b��>��%?-��>9��BŽ��>{�"?��X?�q^?�K?���=��ν$p�<���=�S潽�
<��=}�ȼ����߽O�s���3=(˔<�(�,NQ�]��=�0��m	7<Mɇ�j%�>�A?��>�q�>^�(���Q���P�;+��y4�=iU1�&�>1� ?Ĺ�>/M?��>���>;�=w�k��V��ȍ�>�Ĕ>�h*���o�� ߽��<��>�j?�h?(X�<-$\��s�=�e����=�>�a;?BQ?��>΅�<O��� Vѿ����E7��b�l]�=��a�
$�!Z��G��)�-��V2���ʽ��[>��V>Z�6>fx!>�=m�M>F��>���=.�>�Z�='na=r
�3O�,���BQ����=�0��o=��|��o<�P��+=N)�=����lQ<��?��S?��;�.T�A!��o��Ƽ�\2�>�Q?�g4?�f�>PNa=Z��J�Q�/`3���i�]�?�.z?�Y?ν�"�<\n5�mv��·�>���>3V>�/�j��=$�&=:�>N8?�M�>rH��v�����t�;���כ>_�><�ؽ?b�N?�@���d��'0��G���C\�<�w<��%���K����6�Rx޾ � ��v����x=���>;ܭ?��o�*�=��ľ9ך�(���%���-5j=3��>�>�O�=;y��Ґ��.�됿�������ʌm>���=��>M�?�~?U�U?�S�>�	�>@.�#?_p�>� ?�"�>�?�4?�&�>y">:v�>���=�t�=e���Ȧ�ɐ�=��=4�H>Pg�>�a%>����g]��5��=��J>d<�<	��P"��֢�%��=���=!�>��u>\{?�(?T�����B���:�ӽ�rü*�>T��>��=w�-�8�8��$�>7!?�t?�<�>p�=�lԾ��¾������<_.?��9?���>�=3"�=�o�V��B��=.|�>��˼�S���:ݾ�x��!�����>�m>��=RC>�Fn?�n?� ?`��!S2��M���S`�����~�_�%>AV�=��>u޿=��oPU���@�G�W�N0��ft ��N�=�=�O�>��z>,�S��>8�1�4�q��jB���>$7�=_u�=�� ?��?��.=n)?>��I��M���H?XY���S�n{�� ʾu�J��K
>�B>C�ѽ#�?�t�%ux����s>��A�>��?���?�ie?�o5����>�m>��L>���=['���D� 6�B��S>)}�=�i~�r���ɝ��IG>�q>9��UǾ�[ܾ�T^�R1��s�,�vr�=��ھ�i���aݾɤ��<84��K��aG�I���r�����߼rp1��?(�YP���Qƾ��پ3;?�n�?$`������S��o?�u8��D�E>��)��Y���!$�-����I�hB��{8��1�� �W�\�Q��:�� �>�I�=���0���!P�+�^=�T�>��s?F����V��D�	C�z�q>WT���焾aǊ��⨿kXM�1�1?�.?=˲�G\[�F�M=���Z��>���>�:T>
�j��=t�>
G?��X?�[ >���U藿��]�3��?�M�?'4)?����C����0���(�>�b-?��>E��B&���<���5?�s?�ͨ>�>����u�C�<�>|M?u����s>�1?���>��8��H۾����)��Ȁ�wg�>䐩=�Ȼ1�����ƽ�w����>��>q���DK���͏> Y�c#���>���*���㽘��<��>!O���=*�>9�>���Y�{�I������	?�z�?܆U?_ ?�A�X8�?��x��>�:�>��n>Ksr=�lE��k�>Gx���P�ukJ���Ⱦ[,?�X�?���?!m?\m���ҿ�q�����r&����(>��N>C}L>���v��=c2��M�R��G�7�=N`�>5�>Ǌ>�W#>��L>S�>���h>��6��,��,�2�����q(�"���+�`�y��@	�H˾a+��Ј������`��/+��ͅ���z�M฾�O�>�>�>�?N>��>Lu6>٥>?�N��X4�A���]9���=�U6!��9�I��l?�����˼�C�m<��%�����>��u��_�=.�?��ὠ|>��?\����&�>���>���>�l>�RI>]�l>T��>�˅>?i=�Su>�؏=�������?x;��`��S<��D?�p]�Cm����4�'uؾ}*���P>&�?MvJ>|�(��$��@�w��2�>P�J�4�v����Z�缃a�>7p�>�=I��:|"+�e�{�׋�g�=�H�>05>d����␾{��w�=7_�>_�/Jo>mj�>�t8?]�d?"�? �U>�]�>ĄF>̼�>�T���D����>Ӌ�>nW#?YX?��??O<�>Q��=�#�rh=��F=�N�@\��v_��*�=��<��=���q㽶׺�0i�=��=�֡<��Ľ)���5	ünn�>0<?&s�>�,�>Z�ν�C�t�I�9`Y��V>���=��>���>��	?g�>���>E��>�<>=�η���K�>��>?�<���~�������O>���>1L?�V?GX�=>���U˽#���&�2>�W�>�?��>�s>z�i;���fmӿ�$���!�,���?I��҈;b�<��M����7F�-����͜�<��\>��>�p>,E>ٮ>=3>�R�>	IG>�ӄ=g�=���;�;Y�E���M=���CG<k�P�����2Ƽ��������I���>�[A��Hټ7� ?ʚM?�3�,�g��,7�"޻�`���|��>gG2?j�Q?��>�?g�����<7�e���dX?�d?#��>�G"����=�Ҏ�k�)�nW�>�w�>�Vm=�]
��$���ɾ��P��?�m�>�>y>�	���A��y�������> ��<l�V�
}�?�[?��־�Pv���%��;�q�վz�u�p��^!F�&޳�i,H�Q=<��3��W �����\O(=���>(_�?������#>��z�����փ�0��ю��'��*?��:>
W�������w��l0���R̼�N>�k�>�"_>;��>�X4?zV?�7'?/x�>���<q�?�J>ȝ?e�>5X�>?J�>�+�>�
?�G?҅K>������y�6c�����<!�$>8�=��>�,X>���=��5�<�	�= ��6�.=B�=V�A=ҧ,=�>AH�>���=dS?H	/??	�{< `)==�������Q��Xi>%��6u,��x�=|�n>�~�>�A)?s� ?V1�=jT������ᾙ�U<��?�Q9?6o�>q��=�2>i簾��9�f�@=�~�>���7Ƭ������r��}�::ݽ>�8�>��>��=�N�?��7?y
?gO�N���D���^h�2�����ٽ$�0>��>�8>eV�� ���@F�HK�_5�Wx����$���> c=�e���->�S>C�=�/��ٽD��j��-��=ߏ�=:�?/_?�$?��>%7�=RN��)��J?SI������D���Vξ�#��>�fE>��Ľů?0��(k~�x\���;�>��>��?�:�?L�e?8F�����l>��N>?J�=�;/:�,ۼ�Wa��3J>�H�=U�q�JԖ�
@�'9U>9&]>�3ٽ�/ž�?߾R�0 ݿ�L���=�N������,���%�p�ʾn��٥W��
ξV��2=_�=�P=�^5��3Ⱦk�A��{�b�x?T˂?�#�=v� �.H�6w�!��j">ϟ����Ļ6���U">�e�.����?��k4�!�9����%��>����Q���s��=�'��ʾ��?̂?%mȾ����A��L�>s9d>C�c� ��� '��,���h���%3?�fM?���,C�}��S�;>��*?\1?��>ޖ���Ƚ,�
>=H�>�R,?�_�<����Qz�����?���?��=?���b�Y�[!�:��#�/>��,?9�>�
�O�H���y��q?� ?'�=�������U��?�׍?����I>��H?i>�>�~����t������*�6�>�w�<* T�	����C�O�Ƽ�ï>���=06u�L�¾R��>�*꾪�N�'�H��������Ď<�?��*<>�i>�L>?�(����͉����m�L?���?ÌS?�h8?:����������=d�>���>��=��l�>!��>@k�G|r�����?wG�?��?HVZ?�m�>~ɿ�|���!_�ȇ��w��=�L�=o�=\���$�= �=�ly=�蟻[�=�E�>�Ǌ>NGV>�c>>~9>a4�=8��ہ��9��x ���$_�3]0�����`����LɄ�m��b���:�Ҿ�6=�!�4���ཤ&��k W���O�	�������>�)>��>6�w>��>>b���\%�?*̾���K<�]ھ$�����Gf ��D���H��OlI�����;$���>��)>�4�>A� ?B��hʮ=�#�>��˽�_�>�*=c=0=BOd>��>��>C2�>�o>w�>�����=
���@��+�M�`u�w)#>�r]?	�3����c��̾�#�D��(d?[��>�F�1�������%?X$&��R���� �ES=}?�K?!QZ>[��eH>��-����v�ƱI>��->�aK>�3�<9��U�i��k�>=j;?�09�>_H=�+3?1V?J��?a�>?�<�Y�>b��>��%?-��>9��BŽ��>{�"?��X?�q^?�K?���=��ν$p�<���=�S潽�
<��=}�ȼ����߽O�s���3=(˔<�(�,NQ�]��=�0��m	7<Mɇ�j%�>�A?��>�q�>^�(���Q���P�;+��y4�=iU1�&�>1� ?Ĺ�>/M?��>���>;�=w�k��V��ȍ�>�Ĕ>�h*���o�� ߽��<��>�j?�h?(X�<-$\��s�=�e����=�>�a;?BQ?��>΅�<O��� Vѿ����E7��b�l]�=��a�
$�!Z��G��)�-��V2���ʽ��[>��V>Z�6>fx!>�=m�M>F��>���=.�>�Z�='na=r
�3O�,���BQ����=�0��o=��|��o<�P��+=N)�=����lQ<��?��S?��;�.T�A!��o��Ƽ�\2�>�Q?�g4?�f�>PNa=Z��J�Q�/`3���i�]�?�.z?�Y?ν�"�<\n5�mv��·�>���>3V>�/�j��=$�&=:�>N8?�M�>rH��v�����t�;���כ>_�><�ؽ?b�N?�@���d��'0��G���C\�<�w<��%���K����6�Rx޾ � ��v����x=���>;ܭ?��o�*�=��ľ9ך�(���%���-5j=3��>�>�O�=;y��Ґ��.�됿�������ʌm>���=��>M�?�~?U�U?�S�>�	�>@.�#?_p�>� ?�"�>�?�4?�&�>y">:v�>���=�t�=e���Ȧ�ɐ�=��=4�H>Pg�>�a%>����g]��5��=��J>d<�<	��P"��֢�%��=���=!�>��u>\{?�(?T�����B���:�ӽ�rü*�>T��>��=w�-�8�8��$�>7!?�t?�<�>p�=�lԾ��¾������<_.?��9?���>�=3"�=�o�V��B��=.|�>��˼�S���:ݾ�x��!�����>�m>��=RC>�Fn?�n?� ?`��!S2��M���S`�����~�_�%>AV�=��>u޿=��oPU���@�G�W�N0��ft ��N�=�=�O�>��z>,�S��>8�1�4�q��jB���>$7�=_u�=�� ?��?��.=n)?>��I��M���H?XY���S�n{�� ʾu�J��K
>�B>C�ѽ#�?�t�%ux����s>��A�>��?���?�ie?�o5����>�m>��L>���=['���D� 6�B��S>)}�=�i~�r���ɝ��IG>�q>9��UǾ�[ܾ�T^�R1��s�,�vr�=��ھ�i���aݾɤ��<84��K��aG�I���r�����߼rp1��?(�YP���Qƾ��پ3;?�n�?$`������S��o?�u8��D�E>��)��Y���!$�-����I�hB��{8��1�� �W�\�Q��:�� �>�I�=���0���!P�+�^=�T�>��s?F����V��D�	C�z�q>WT���焾aǊ��⨿kXM�1�1?�.?=˲�G\[�F�M=���Z��>���>�:T>
�j��=t�>
G?��X?�[ >���U藿��]�3��?�M�?'4)?����C����0���(�>�b-?��>E��B&���<���5?�s?�ͨ>�>����u�C�<�>|M?u����s>�1?���>��8��H۾����)��Ȁ�wg�>䐩=�Ȼ1�����ƽ�w����>��>q���DK��<�>�q��A���=�}���.����� ��>��׾qwk>��q>�Zr>�4��3�� ���j���?�P�?��[?;�$?M �c�r�Dk�=��&=��m>,��>n����7�xR�>�1�>��d䅿`R��!? ��?{�?\J?7;r��ё�߾z�'r��1Ʃ��!�=�+>�>�>_���6�=A��;��¼1p};��>���>w�><$�>l܀>M��=3�&>�����,x���餿��Z���.��?о1\���v��#��Cj$��%¾��ξIJ��� =�޽�'ھRޫ�<��7*���>T��>ƌ]>��=d�
>q��=,��7����z��D�=?!�l����o��0��
����Y������`Z��*ڼVj��\/�>���s�
>'��>���<`(�=_p�>��=Ee�=�v>^8�>L��>��>��5>�dn>�q>��>ЮN>-�r=<b��s����`K�亇�V3y>�Z?ᆂ��uվ/�@�ػ���Ἶ�S>gS&?�5I>�67�a2����f��>���i��S��)�=AG�=��>��B>}��0DG�nk�doN����W�=�\.>��3�;�E���J<�>��UJ>�O�>�j;?Y.v?��?�1ػ3��>�!�>$l�>޹d>���>	j�>n�>%H(?�N?o^#?���>�,+>}�ɽQ��=���<g�.���	������x���!�=��=a�?=�;=V̖�O=b<k��=��=�7�=R�?��E?���>�F�>��JP��wF�bi��;��>hY�=Q��>͹�>,�?���>��>z$�>	�3>�VF��>�����>��>hF�C�q�&7�=�|�>R�V>űv?��a?��F������Xx�=M\?uQr>8?�d>��=�]i�����ӿ�j#��<!�6'��������;i�=���O�8�y;I1�)���游<~?Z>L��>��p>̴D>|c>=#3>:?�>6�F>�Ԇ=�z�=��;�=�:��E�w�F=�	���7<��X�������p���sh��O}@�n�>����=���?��?���\����g�]�����x�>@/�>�B�>4��>r��=+���.T��A�xWD�!��>�"h?���>?�8����=��&�ם0:�r�>�2�>��>�I��4��S��XL�<��>@?��>�����X�� m�
��>�>��ɻ�*6���?;U^?Ȯ��6ϊ�ʌ ���S�kE��H�=��t�p�~�l������ξ�z�􇾈� ;4A�>��?�M��%=6$;*_��7���4��P�=M/佈�>?@>�L��F\A�_r�^{˾��F���T�ّ6>��	>r#�>v�?!1?��w?�G+?��R>0���?	vO>��>�t�>�Y-?��+?"��>�?�c�>��μC.}�tf<��龇����=��>BE�>:٧>;�/�	q���>�4�=�>p	g�&n(�X�=|��=p-�=�7[>a��>p�?��*?�鞽ɱ1�u����}�$V�<�
>+?x>~P/���g�KGڼ@�m>6
?'?+4�>��=��ھ����L�r�=��
?��*?P��><X�=d9�=(ؾ��E3�=bk^>X�w��v��
ܾ�ñ��(�3ǃ>���>b2�=_��=�l?�22?N	?Nt��5L�)4l�Y�;�>���7�1���>�҅>��۽�X¾?�)�kQ[�yR�k�������}��[>�c>�)>+�h>�0.>��>���=	Հ��l�%>F�4��\x>J��>�) ?��j>��o>����
���I? 衾�S�۠��yо3���>^�<>��?�����}����?G=���>ez�?���?d?�C��'�Ư\>�6V>�>��2<�>������y3>���=�y�LB�� ��;�\>�ay>Yɽ�ʾ;K侈�J�e8����n�
PI��Չ�V`��L|k�t���G߁��g��1b�=|\!��;��p#���]�⠷�:J��ty�����׉�e��?'�d?��0>0̈́=���͂����ɒ;����j�z��c��ց���Y��⵾�I�����
��+�b�+��N�>Pً�݆���6���޾�I@���>��Z?���,��� �@�սUd�<3�r���t���e������5:?<�1?rBҾ",Ҿ���:·�=� ?��<:c�=�R����ӓ�>��;?��I?Ҹ���s���֥�A�=U��?��?$[3?��d���]��"�8���0�>u��>�(?Ջ��о�{��?ğ(?)�(=�?�����X�6���4?��{?h�V��J�>��?Y��>MG�� N��������w�v=���>I\�=�fF��۾�"1�4��<�a�>��B>r6轚����'�><E��SMk���^��4�����=�?yu �G�p>H��=�j>j����������g�r_"?���?�H�?��?�伾}�ѽ��>.H���&>�>�� �ִ��ei?|�>�'�?����C¾�>���?�V�?4�d?p"��Z�ܿ����签¼�����=��>���>���p�=�RF>2�>�z9<���=6y�>�͖>T�|>��A>{+Q>��9<�ȁ�s�T����܈�:�@�:b'�}��ǡ�؋�hV��X��G�C�;�[�ŹM<(���f�J�y�W'������+�=�V>���>w��=��>�^�>�W��8�qMw�c���;H��</�&#侞�5���%�P��
ؽ2�q���g��W?�Hڽw���h?���G�={4?������>wL?�n>E+>�>���>![>f��>2��=�A/>GT>����"��B�:��Q��cr��An?8牾�J��^zm�0��������/)>��?M�$>�9�\�����q���?gn#����'����Y+>3�>�#?�>$Ž��ͯ���\�^,=O�b>�B>��O�������eV>���>��
�,rU>鴩>���>+z~?G�3?[Y�=VD�>��e�#g�>��7>u�=厶>Aۅ>��?�?B?L� ?$��>�%>(�m���}=%��=��~��+��X =ܳ�O6��z�;t�0��}b=%�=O��=�R�=&R> �3��	>@V[����>@�M?,U? ��>�P ��H0��[�\�%���>Ǒ�;��>�
�>D|!?��>���>`�>E�>�\���^ǾA��>=�>۹6�����M��rlt;W��<h0L?�<]?,Y=�$�����=�d�>�ͯ=��>s�?<��>��?>�G�?Q���տ�� ���S���S6�=s9�9M�ͤq��F�<�k�f������:"�f>kE�>:�n>��B>` >�L>7��>L,|>��=#�=q�ּ�\�*��+S�z(P��ƼWx���=9<��
��o����0���Z���A诽BD���? +?t̂��4�xǾK��"����>�S�>��d?���= �!�`;��e��b�O熾?�>�k?N?,���{L]=�޽k� >���>7��>��}>ˆ�;K���¾^a�O�1>Ք�>�\?�����|��1C�l:��u�=�H=@f<�H��?^�Q?���z� �jD�T�V��B�|�x����@����������O=��]�������=MN�>6��?���6�4>g����U��e���u۾�ϙ��Bj���>�4`<�&;�Vr�|�� �־�۪��B߽�k�=��g>A�3>!�?�41?ėy?�9?Z*�>�b	���?AA�B��>��>i�>��?��?+��>���>ӱ^�3o߽| ���<��o�R<վ>j[V>���>I��>T��:~⽄��;5A> +�Ȅ�0����;褳=�� >��>�D>��?g�1?]R</��;�W�= ��q�ky>vǦ>p�����X�y�<�k�>��
?�).?���>��=2B��>�����M�	=��?�.?�Q?��>���=e¾�P����<-
@>�5ۼe��X��j�s�tϽz�?>ٻ>�x>�eN>�j?��(?��%?A4��Q6���v��]�����H����>:��>̡Z>��ӽ���m�C��
]��#��������.��=!�>�$>��5>08���?��6�=oTu=axl=P�2>1�=v�?>�>A5?U/�>9$G>O �����#�I?�U��N=�������Ҿ�{8���>��;>9I��X?.��a'~��6��>�Ɲ�>Ţ�?��?�e?=?������[>��\>��>*^�;�6?�!��ܮ���2>���=W�z��4���e4�F3^>�w>��ʽb�ʾ�L���`��ȿ+@?��b�ۺ��$ �U.�8g �!��	Y��L_��Gо��=>�{�x# �*8T=�R�h~���������$�?�(�?�Qg=e��^"�).��_�kxQ>۹�n�c�)�5"2�R�L���Ҿ���o����D�9L3�t����>\T���˷��I���/�����>B�>k)o?�.��	�+�W��$>��>��q��˰�����|��R�S�}�Z?��6?������	��y�5>�=�>!�>���BN�@j���|�>�&F?��<?�����Ի�+�����=(��?���?�B?d�H�*mO����[��j��>�
?�>�T���꺾��!���?}�7?~�y>���}I��B����?��p?N�E���c>ј�>��>��@�\�����>�����h���D��>�-~<>:J�4Ώ�!�@�%�D<�n�>���>���3����a�>�Y־�R{��A���G�L!�6�+�z)(?Ԍ����=��>�:�=�kO������8���z>�Z/?c��?
$C?��d?B�4�i�A����̈́���"	?6�?���x��"i�>�t�>���}vA�{2����>d�?���?K�t?;
_��7տ�H��r���]qľ )�= 1>�YL>��O��=P�> ��=+ �<�d>�^�>7�^>{�3>��>���=k��=u��9����چ�53�������T�CO	��
����4j��ҾKw���$��X��F�V�S�$�h"�������s=��P>� >v�>Ν�>�ͽݴ��'��V㺾9��ic,�x��n�j�
�@};҈��Ḿ�����f?=���G��>��'=ց:=,;>uy���I�=<�2>JJ�;��<z�>�����}=�G�=�>�O>In'>Ƭ=�U�>�SU=������c�;���R��=|YE?�N��� �6��v�vձ�1�>�
?BFf>��"�G��Gs�ī�>�Ƅ��9E��ٽ�����}>Ԣ�>�q�=��W�a{�T&뽸�=~~�>��>c�¼M��}X!�ŝ�=k��>��ȾB>$�=>�K2?�v?G7:?���=��>��>1]�>�N/>���>��>*�>��?�=+?��-?�{?W�=��]��0��:�=ĬF�Ϟ���ݼfS$��O����)�y�;�b��=	��%�<���=rBe<�a�,鎽��?p�G?8��>���>����]o���[��׻�O�>��O�8�?��#?�E?+�?j�>zʡ�~��/"��/�����>�0>XD���w�^��ѻk�>�HG?]"&?�ѽ���]U>�t�>�F�>��9?wD?!�>���Y�����ǏƿY8"�±� �k��/e<Gݣ�RG5��������88�a8��=��=��=|�=���=���=-�&>7��>�d>�Ѝ=箉=��!<��ż��v�!o=%�5U�ħ������X�H,��y����c�5�C�Q��L���$?�V>?-Z���>L��0˾o��خ�y��>-�=CV>��+�/�:���?�Q��P����?h8�?���>�F���d=*�=��>�5;>�k�>O3>^��<�Š=">��RJ >tv ?� ?���>�4�&�<��^�����K/�>�fJ=5P��"ǆ?�MC?��sGq����=;�<2�}�F����搾�m˾�p)�%�-�����޾rQ�g��<�?���?L��N:>rW�����>�h���оo��Dgֽ�o�>�в>�fֽ�Užce���q��3=zu>l��> �]��b>[�n?Pӑ>N�?.|?�_T?0�,���=��$?�>?�dG?�D?�KZ?h)?wVл����!W>��.>�|ý�rf�i_!��ý��=5�>�@>��Ƚ��W��Bv=6�|=S�/�kIx=�>wX����T�v��=��=*6a>��?<�&?*u�琎=�콩����'���=�>�6�mh����=�k\> 1?�S?vu�>���V����K%���c>}�U?��>�T8?��x>ZH�>g�;��ƾ�Ǝ>��>��-�r�/���I�a������>1�>�$}��
�>��|?ԓ/?�J?ڂ��	�A^c��|��u>�����g�>x��>l�>����s4���T��}q���0�P�i=O.����[��y>>��*=�=������<ד>>�֭�@=^,I>+��=G�?� �>.��>=�h��阽KҾ>���<e?ݏ'�i�L��K�L�3����=>��>��>3B9>��?���!��d+q��渾�8
?��?�0�?�/7?�
<_Dؽ�>5��>�!�>s�=9������1�=G�d>s/�<�lҾk�ھ���<��$?x�?�C콍���x'���S>/Ͽ/�Ta��U�������7�ț���$�����" l�K�޾"�ʾ�nؽ�۾C����ٲ��o���蘾���Z@}?��l?�#�<'>tFϾ�� ����yV';-2f�@�w�kv;�x��]b��'���f��xξOU�7"�0+���>Q3Y��-����|�;�(�?����`?>�/?�wƾ��б��f=� %>��<�,ﾄ���ۗ����
�b<W?��9?���̉���Fཥ,>~�?a?�>�%>���݈7�>JE4?�-?�&����; ���Ǎ�:l�?��?��??8�N���A�������n?�?���>N����;5���x�
?C�9?u�>G��5������z�>�Z?&N�z=b>�I�>� �>D��ና���)��/��m?��6:>���=�fCh��=��=�x�>_qy>��\�4>�����=����C�H��W'�-�H.8����ŭ>�׾�JQ=���;�9�������2���ש�:�i?���?FQ;?:�r?�B�T��VF��5̾.��> �4?�ǲ>�5>SE?��S>����\�({G���?>��?�<�?�M?�.O�N�ѿ�H���|�L���dfW>>o�=��=�1��=���=Bԓ��O�aw�=�J>�s,>T�6>�\">P�P>]>zd���q �5�����A�N����.�X%��R���W��W�:�8�1 �{#��w�����&���c�i�t���-�-υ�����0?�-�>��(>�>b
=��9��1��=��������">�H����s��|�"���q�,��!̾3���G��b�>��=)�>�t?^Ç����č�>R��=��>��7>Oݯ=��=���=\�>f�=R>`�O=ag>rsE>$��m����)�]�W<�� >v�@?�*ɽ2|U�Mn&�$Q��C�?���>�w?�?:>S(����,�}��?�>\��vd)�.� �G���m>��>�@�=����i��6A�;ҼmL�;��=��X>x�=u涾b�g�:��=v��>&�ľ��=6!m>O&?a.v?�U6?���=�o�>��[>]��>V0�=�?H>��Z>Ԅ>4�?�5?�,.?�c�>��=)zV�=�<�>�<�:6�9Q&�/���[���+��5=vt�u��<�c`=ؐ�<�w~=�.=��ϼe��;,'=8Q?�B-?�&�>���>�3�j�(����;��>.�<���#?#s?�$?�?o��>S
�l[��ڹ�Gʾ�ڔ>P��>��I��T������[>�A>,(8?�d?[�d��S���0�<���>u<?{<?f?�M�>�g�<i>t��J	���ѿ*!������'�G}��NK��*M�/������˃=�b^��Jc<u�H>�Mh>hX>`�8>�>�m>���>=�J>u=Ch�=�1�:Z$�:u�R���E=���N�.<4B�s�q��#�0��菥�;xR�͋E���'�������?A�?��= :�=�۾%����G�>��=�ݨ=d�
?��f=t"���f��C��[���>(�[?*�M?�W�,�'��*�=Jp(>��A>��>8�
>�u�=o�l�槿�;�>M�*?ڮ? �>����8�Ҡo��&��4�>n(,>���J�?uEs?�7ܾ����⾐�\��02��Z��%��7�����%��:����,��W�ƽʉ"=ܚ�>�`�?���9>7ϛ��ܓ��}��a�� ������C?�e�>�k>�ͻ��~
��t�D�*���=���>�M�=�� ?�x�>�l/�G=Q?>OP?߼c?�=���>�_�>�>-?T�j?��k?�D;?躽h�D�������T������{��i=�ۥ<���=��=�G�<v���}�8�|�>v�b=	藻qG=S$Z��c��������>t�=>�o�=7D?J %?�����[�=ꧼ��ӽ�[�=f)>&M�>�Qg�m�8>�S�>��>���>�PL?3��>r*���o�.e�4��>�>?ʅ$?&�6?9�F>�o�>_��.c�"ر>���='����ULɾ�'����<��g>5��>�f�=���>�W?R�B?>L?��k��e�DZ�|�*�)�ʽ����i�>aE�>�\�3�㾄�)�ƳQ��@M�6A���>A���R�A�̮=$C8>�,�>?E�>#�>�	�V"=<b]��>,��x�/����>B,?�A?Ó>�'���O���#� [?�5B�jn��0���K�%�ھ���=-�8?{�>�o?�־_~��T����_ܾ���>��?�q�?ol?<?C;<��ы4>$�?�$&>C�>=���:�����w3K;�S��a���а�c4>�V�>:3�����`Q�ۅ�{T㿣z\��'������L>�<���{�E�˾	Ⱦ�^����^�����/ʾ���ᾙ�����߾4h��a?�?A?�_���}������ĕ��p=2hM���H�Cu�wH]�G���%���4���׾�a����|֮�S> �w�.����{f��`�Y��L���*�?�iþ���*��f�<�>�ν�#��Ċ�6����R��?V?��;?�T�� f���齚�D=���>X��>�s>��y�ݺ|���>:U.?.�1?WĽ��h��{���������?PY�?WV>?H�A�7A�M�
�|�e?�?_2�>�[����Ⱦ���0�
?S@;?F-�>"� �b[�����5i�>�vV?/M��Mb>��>3e�>A��������3����j���6>����T��&ai���E���=���>7�q>�gc�&\���_?u�߾4C�������Fa��m��5O���$?�C�-G�>��y>��S=�V3��_��U���΃^��W?Ly�?�`?�>F?�$�>-����b̾��?L;;?���f�1G=���>��]��� a��-?
k�?�@ES?14E�]�ܿO��g5���=�O�>�N=�3$>�Y��|">^Ѻ=�8��o��hC&>�+�>eQ>b0|>:�>4<>3��>A���� �Z����p����*�]�����A�����ލ�=~��;`B��2N�����S���q���0��l�=O�ѼY�>�??R̟>ifw>؀�>���=J���P����ﾒ5D��<����_�[�޾Mo�^�#�O&���!ܾ��T��S� ��>���<`9�;ф~>:Ŝ�q�b>���>)��=�ʉ>\��=�&>��>q�p*[>�k>��v>�X>����#
>�T�]]n��T
�*���׾4.?�ņ��ž#V⾂x㼎�y�z)�>�@w>+�����1��봿th���}�>�ɔ=� &�Z�g�d�<�g�>�J^>���3����=Z�F�N�n�;/�=�1<>ren=�|�u	L�]�ܼF
�<���>0��l�?>TS^>A�?�"l?�c??��2=��>��#>�mz<k�꼳��:f�=>��>1v
?O�-?ak ?v̤>f�=^�r�Ր�<M�I>�,�Cr�(�k��1m���G��<��q�/�"�yH���R�<�`�ً�`k��Fw��S >'C�>F;?�{?-�?p*�x&+�� W�/�S=�L�>��t��X?�X�>�?�L?a��>�a�>[hT��о�����>�V�>
�\�_��z���w%���=�� ?�
?��2�A�p=[	�>X��>}�?p�?�
�>d��>xg>�4>6���9ݿ#I�5LD���μ��W:�e�<�L"��0<J)u=�m+���	���=�$*>��>3dr>�w>&�U>dp�>��>o[�=ܑ�;�>��_�7KA���<���=Η���{�=
�=�^�=��:�1�1��󲼀����d��ry����?}k,?��
>y8�=#��:��/���9��>�׉>�>}>���>&�M=�:�ݵ`���I�h��w�>XLH?R�?�x��'Ũ��)��81�=-Q>���>H6�?��=�p>��!�Y>�1&?&�?�Qj>���HC�����5�b�>���=_䑼��?9�\?Oݾg�*�ƞ�=�-U뾖�׽����3���پ���S[2��>澾:پQ#����,=���>�7�?P5 ���>O%��j���!���������:_Ƙ:��?��>���;�0���]	�/�¾�&��|�=I<�>���<$�N>[9�>�I?J�?�^+?A�T?5o���Q=�
?&+�>y�??���?C�J?!i<?��<0OƼ3h�<"���-�1�`���l�4��m
�Ɔ=t)R>�i�>�������=�>���:���<�s��=>;@=#Vɼܗ�=��q=6s(>��>a6?��v>Q�\>f97���j�d�A�g>T�>��?��f�=�+>��>wa ?��<?���>/	j��퟾�lƾ�C�M�?=�3?zN?-?f�l>���>J���ᾔ��>]=Gxڽ�I������۾�����%<>p֖>�e�� �`>��[?�!?�#5?��>�w6��5�t��`��>���b�>W��>T�ü��#H�v�a�G�m�NeA�����������"<�?;���<>$�>��=�!>��=i��=��}�8+���������>�ٖ>��>SEw>��E�h�����þ1q?$82��^�[W�T4���ǽC��>��>�NӾ3��>P�;o���oh�������?��?r��?��y?��%>��k����>��N?Q
>��>�rC��cB���e��p���]=���l���!+>��=CM�>Ņ��-$����p�~���ǿ
wK�� e����.v��:���zоqN�G�0�"\j���T��~�V≾m[���b��E���ʗ��8ܾ>C&�v�?�t�?禕��R=jm��FB���6��G��D���d����u��`�=�o��H�?�����J	�<\7�y�m���<�IAX>�T�+���g�� �q���+� *?_Nq���	������=|q�=�5̽v�9�7-������\*��:^?��H?(�;�9���v������>$�>�s?���cd����(>	�?\
�>�4�}�s�hl��w=����?�?��??��O��A����/��-1?Ъ?���>k���s�̾�6��M?e�9?߰�>L�7]���/���>}|[?�.N��Fb>���>xW�>\F𽣞���&�MD����9>��	����Sh��>�;k�=��>�sx>a]�ா�И>�У�`v�J/;�X��_�r2�v�?(��?>��>a�v�*9��Y��rM��������I?�ǹ?��o?a q?Թ��~/��W����Ͼ�^�>�}?&TZ>��=��?��?��׾S�������l3?4�?7�?�Wv?P�^�_�п+���G����Ǿma>wV�=s�J>�H���>�;�=OG�<��=�K>���>�Yz>V[>��R>AQ>�J,>R���wc%�X���m��Z�:�.b��P�p=9�l���{�ǋ�ly���K���r�r�[�x����9��y�z/>���Ѿ��w<r�>D�?>�.�>ai>|Y���s�u^�y�{��`��e@����V]�R ﾜ��ч��%z��/�K�E����y�>��=9��=�!d>j
�!>� �>�R��#6>�d�>	��>?�>A�=EД>P>2D>�>�[�>�5=��n�A��F�8��cӽV��<��L?�1�������5�����2oƾRx�>�E?n�\>����ۑ�WMv�;��>���\��)��@>����>oC�>C��=�T =�Ѧ�U`k��G�� �=(:�>���=![K��]��IH���<
G�>��
�d�j>f;�=r�?$J�?�?^�,��H(><��=���=R��=�5>�s�>�ŭ>�$?{�+?t�>'�?���=[���\�	=?>2���.� ������j�_�=;��s�뽛-N=xܤ=B�W��C���[�=�UC�z8B<��E>e�
?��,?I �>��?�ܾ�B^��]y�X`�9y�>��޽Q6?m�??�4?F�?�Ԥ>��Ӎp���(�)���>;��=��9��[�7���j=��Y>�I?�#=?��:>H�����=yn�=��>?� ?̓.?<?f��>V�l����kӿ�$���!��ނ��B���;��<���M����7P�-�d���~Y�<�}\>��>�zp>�D>*�>E13>�S�> IG>�ń=��=#^�;�3;��E���M=*��@G<t�P�Ф���4Ƽ�������1�I���>�*G� &ټ�*?�=?��l�=?<0���q���~�ͨd>$�>�l�>3��>(X=���Fe}�xu6���g�Ƶ?}��?e�>l�x�]��=�c��X:>H%�>��g>7-->B7�<���<Jx�u`p>D�?�e�>0��>e۽������_���sU>9�=p�s����?loG?�v�@��*��:����zC���R%��K��������+\�g���ݫ߾�曾V8">���>�u�?�1���H�=!���)x���?��I�达����
���?�5�>�ܺ�#슾g��^ֹ���Ἧ�4>���=3#�e_�>��#?�wk>��V?'P�>�&D?U^����>�;�>��?� R? j?�
5?�-�>��"�l멽<�>ra�>�;F�b���!����ɷ�;��>�*p= y�`$f<�:8=�N��h>=j`�=�%���^<S�h<���=��%>cq>�q?&��>L
��`� >B\W�uSk����<�>�3�=����k9���_�M>љ?ŵ=?�5?	�>ޑ����m���T�>۝#?ӌ?,OM?�[<>�G�=�m����v��D>L� ����$'����C��lE>�,>�<�7>Ȏ�?��+?�j?S~)��K#����1���C=>��ž��>*(�>yM�=�7�����pe���~�������+���i���C>�>j�>�5>$�>}�=>m����>;H>O�=r-�>+��>���>yɦ=�W�ڣ�{I���k?P��F�d���A$��E�=�%�>�I>#��=�$�>������;��������?f��?�V�?S'=?= ����R;�=�G�>�c=ɹ��T��$D���KA>��>��">�3޾�[��%>)̊>c6�>nb��]�� �{�ż݉ۿL���ӽl[v���=��dnǾ����E�P�l������վ]���3UӾJmþ�6��mξR��?�+|?��<y��=[���$�������8䱾��z�^�ξ�V��
�� 8����#����W�"�Ne���$>�BN��ܑ��Y������򖼓�?۱þ@,��,-����<N	>H�������T���ј���-�c�[?��7?rɱ�b�ؾ���<G=���>��>�p�>��Ng�랝>`�?��1?C�˕{�U�t�;+�=#�?z��?T�??�P�|�A���6���K?8�?S��>������̾�`�<$?��9?�>w���D������>�[?6N��gb>,n�>�K�>��TD��'�Af���	����9>�F�9���g�$>��=7۠>dx>��\�����a�>�Y־�R{��A���G�L!�6�+�z)(?Ԍ����=��>�:�=�kO������8���z>�Z/?c��?
$C?��d?B�4�i�A����̈́���"	?6�?���x��"i�>�t�>���}vA�{2����>d�?���?K�t?;
_��7տ�H��r���]qľ )�= 1>�YL>��O��=P�> ��=+ �<�d>�^�>7�^>{�3>��>���=k��=u��9����چ�53�������T�CO	��
����4j��ҾKw���$��X��F�V�S�$�h"�������s=��P>� >v�>Ν�>�ͽݴ��'��V㺾9��ic,�x��n�j�
�@};҈��Ḿ�����f?=���G��>��'=ց:=,;>uy���I�=<�2>JJ�;��<z�>�����}=�G�=�>�O>In'>Ƭ=�U�>�SU=������c�;���R��=|YE?�N��� �6��v�vձ�1�>�
?BFf>��"�G��Gs�ī�>�Ƅ��9E��ٽ�����}>Ԣ�>�q�=��W�a{�T&뽸�=~~�>��>c�¼M��}X!�ŝ�=k��>��ȾB>$�=>�K2?�v?G7:?���=��>��>1]�>�N/>���>��>*�>��?�=+?��-?�{?W�=��]��0��:�=ĬF�Ϟ���ݼfS$��O����)�y�;�b��=	��%�<���=rBe<�a�,鎽��?p�G?8��>���>����]o���[��׻�O�>��O�8�?��#?�E?+�?j�>zʡ�~��/"��/�����>�0>XD���w�^��ѻk�>�HG?]"&?�ѽ���]U>�t�>�F�>��9?wD?!�>���Y�����ǏƿY8"�±� �k��/e<Gݣ�RG5��������88�a8��=��=��=|�=���=���=-�&>7��>�d>�Ѝ=箉=��!<��ż��v�!o=%�5U�ħ������X�H,��y����c�5�C�Q��L���$?�V>?-Z���>L��0˾o��خ�y��>-�=CV>��+�/�:���?�Q��P����?h8�?���>�F���d=*�=��>�5;>�k�>O3>^��<�Š=">��RJ >tv ?� ?���>�4�&�<��^�����K/�>�fJ=5P��"ǆ?�MC?��sGq����=;�<2�}�F����搾�m˾�p)�%�-�����޾rQ�g��<�?���?L��N:>rW�����>�h���оo��Dgֽ�o�>�в>�fֽ�Užce���q��3=zu>l��> �]��b>[�n?Pӑ>N�?.|?�_T?0�,���=��$?�>?�dG?�D?�KZ?h)?wVл����!W>��.>�|ý�rf�i_!��ý��=5�>�@>��Ƚ��W��Bv=6�|=S�/�kIx=�>wX����T�v��=��=*6a>��?<�&?*u�琎=�콩����'���=�>�6�mh����=�k\> 1?�S?vu�>���V����K%���c>}�U?��>�T8?��x>ZH�>g�;��ƾ�Ǝ>��>��-�r�/���I�a������>1�>�$}��
�>��|?ԓ/?�J?ڂ��	�A^c��|��u>�����g�>x��>l�>����s4���T��}q���0�P�i=O.����[��y>>��*=�=������<ד>>�֭�@=^,I>+��=G�?� �>.��>=�h��阽KҾ>���<e?ݏ'�i�L��K�L�3����=>��>��>3B9>��?���!��d+q��渾�8
?��?�0�?�/7?�
<_Dؽ�>5��>�!�>s�=9������1�=G�d>s/�<�lҾk�ھ���<��$?x�?�C콍���x'���S>/Ͽ/�Ta��U�������7�ț���$�����" l�K�޾"�ʾ�nؽ�۾C����ٲ��o���蘾���Z@}?��l?�#�<'>tFϾ�� ����yV';-2f�@�w�kv;�x��]b��'���f��xξOU�7"�0+���>Q3Y��-����|�;�(�?����`?>�/?�wƾ��б��f=� %>��<�,ﾄ���ۗ����
�b<W?��9?���̉���Fཥ,>~�?a?�>�%>���݈7�>JE4?�-?�&����; ���Ǎ�:l�?��?��??8�N���A�������n?�?���>N����;5���x�
?C�9?u�>G��5������z�>�Z?&N�z=b>�I�>� �>D��ና���)��/��m?��6:>���=�fCh��=��=�x�>_qy>��\�4>��vr�>HO%��!#�b]�[ ���0����>uC�>�g6��.��(}?𼃉'��Ӛ�����cq��F�e? �?�e-?��w?���^-S�,� �ng�=�I?=��>���=o�;�vM>x8>?�@�d�4��Tɾg2$?A��?O��?�V?��:��տ
�������O�����=_��=k#>��V��3�=�u&=��_:A��[�!>���>h�I>�]>�1>ݠ>pU>�*��b5(�����mB���O�u��U�"��"������tF|�=��<X��j%��Š���� ������s;��6��n��r��ȼ�p8?z҈>l�>�
�Z�>����&�)'�M���5����,��O{��ψ���W��#h���}�2�R=O,�d!?�����E!=JcV>V����>�e�=|4>[�s>Z�>��]>��$=���`�=��h>���>�g�=���>�y>��}��������������7�N?C�Ž= ���8���ƾ�v��|�>��
?cVz>Z0�B܏�37�����>���<��b��z ���e=E�>�W�>/�N=��<Up=��[�	SνJ"G=}��>-��=�W=/D��/��dN��C�>�tҾm_�=�|>�)(?7�u?�6?�ɘ=�r�>Z�c>3p�>5�=�	S>�Q>擊>a�?��8?W�/?�*�>@��=�Aa�Ե0=�G=�4D�'�c��&��6R!�R���ו<[l=�ھE=�Lu=%� <1�W=h�F=*S����;4a�<�?+=??�T�>���> ~��r����`�czQ>�q�>Q~��~�>��?"�2?�?�a�>s��݂þ{Nﾹ1a��s�>���=E�̧��RS�>���>�|�=�o?�A?��ս�M�Ͻ�]>�V#?A?�M`?�>_���� �y������M��{�վ������8����a����d=ա<�靾:��}	M>���=�kl>�>�=�H=��=�	�>��=p悼,V>|T��`{=��<{� ��頼2Z��!w��Y�9��c�A�k��ݷ;ݨ�A�����;3��=e2?^�>a�=�F0>)I����,��M޽�b�>�>6�p? & ?˻>������p�aC�����>�Ƅ?RR?�,>�ʩ>7��j��>?��=�+�=H�X>�F��
�N��T�=VB?#�)?��>����t�6h���$�A��>	;�<�6?�(/�?@�F?u���y���	�VW9��!���0>�|#�߾��e�ܾ�8/�i�4���߾R�ؾ��Tl�=��?@}�?g���aG=�����ꊿM���n���> �>�)�>g %>�\������-9��վ��K=���>���>���8�?
n*?^+F?7�s?���>�!>`Q���(!?�����Y>N�?�y7?��?w4�>�~>FE=��ƾև��T�p��M����=������<���=��>���Rֻ���W3�=����LP����r?�������A=�2>�>��?��W?чҾ9�����?��>;9���ur>(�>����r4���>7V?��9?.��>���>8�G�p���?��뾳`��U�>�$?E�>�Ke�{̷=P���V��<�<t�/>�B�=S���-�ݾ3�`�H�����>��">�� >��c>��{?.�*?lk\?�]���K�O`6�t�zG>k�M=n�>���>y>�J˾[�-��~��X�ln��F�=v�B�r�=ZT*>�'2>� >�Ľ=c)ʽ�A=��>�bh�O�h=�3 �l��>�{�>H�?�M>�����>�~b����S?��5��
>о[����=��>I��>���ȣ>���=���蕩�mU��I?�t�?��?aGY?��=E>>��>DuP>��>R�+��ξ�=�97>�1>��A>�-��$�c���>��>ԍҽ��ľ8R�;���G���DSS��'��J��~���<�;�%��fN���}�����i��~���z$���m����!��E~�<ڲ�X����h��xL�?�A�?��>�U�����
/������?5>�����=��m����|��~��r��&&���/�s-"��ƾϴ�>U�Y��9����|�S�(��A���u?>T//?Cgƾ�Ѵ�d����g=V%>K�<?D�}���-���N�7cW?�9?
N�6&��%��>t�?�z�>��%>f+���P�/�>�54?G�-?���\��/7��.Œ�%m�?h��? @??�[D��#A���,�qW?��	?n��>w���].Ǿ��N?	:9?�μ>�f�҄��A���>ZY?�YR�_>2��>�&�>����+g���#��얾'w��e4<>�0��]�>�c���A�a��=�7�>q�t>ڃY�烮�l��>�v��侖�_�(�̾��P��Z�>�{�>Z(���>?־>o}t���9��֌�i����4��n?�Ż?tYh?�}?ݢ3���_���ćD��bW?��>��>�/��e�>Ln<?`#����Z��e��2?�?��?��|?A�g�L�ӿ�c��������о���Y����%0����&6�=�缑��;�u�<�W=��j>K	1>?ob>[#>SP(>��B>B���,'��؋��ύ�Ƥ^��v)�"���C�����8&��侻�˾h�ľ|��%�7�i���M�i�Mc�BF㽽����>>�!?�<�>���>@��݁>d����&�����۾�w���(N���{ �,B�����c���ڲ��8=p���
?����C3>�#�>'e�<���<��>�rU>Z�>P�<>�;5=�">�#>�*>�ߏ>�:�>䑐>��>� ��!�����x��S�K����~�=��J?�����x�PA�w�3�ק���#?!�R?"˭>޾������F�en>�z>h���F�,�G=�*"�=[�>�ҕ=''j=S�5�����mJ�=JE>̷>�J�<ĸ�+����l�.��=s,�>�G׾>W�=zek>�'?��t?64?s$�==��>�;a>?B�>��=IRF>��_>p�>R�?Oh8?�2.?���>W��=�__�B|=!�:=�T�71��r�����jm'�. �;-�n�,d�=	<W=ƲF�!�!=}�]=�Y��,��<��K=,?n�?2��>��>P�ݾS+�՚�}�2>wC>
��=1�>8��>$p(?�~?�?�=y �=5�����!�¾k?�>|>�셿B���C|">���>��>f�?l�
?�fɾo�=��G�B�>v^%?h�?h�?�p�>���=���e ��f̿�Gw�ڈ�0���S.��G�� &ݽ'>�F=����׽��׼�=5s'=��>�e�<��>sɅ>(�>�� >㠊=��<��=�n�=���&X�0�<G>�=1u���H�<��<v�ƽ\>-�u�&�qI=���=�?���> {�>�^>u�B��N�ƮF��m�=�I?��?�>�<w>�:'���f���f���þ}��>ݏ�?��?�Se���3>D>Y<SaX>�`>�9�>�>���[���<�9�=��/?�& ?4��>!R��k��Mz�V�/��>(2�<nw��h�?�hF?g��Ο��_W�|E�
�	�P9�=�d��q5�޶ɾge#��J9�!��>��d�W���@>\?��?#�ͦ �,�ӾLG���X{��-l����]�<i��>0G>ք�T����#�勉�m���=�˝>�U��@�C?I��>�|?{f?9
�>���>-���>f�̾I#?��>?@O?�#�>�a�>?@>>��<z���ӽʖ7�!陾"T�=b�ƽ�CU;3��tyV>�, =.ro>��<�����T�σ��V��=?�,� ʝ=2�=B T=�BT>��?Fh ?H�����T�>n�>�ǡ=��>� =h7���}���h�#!�>�'?5�,?@˓>͕{��4��<�A#�^z>1D�>�O?���>�I�;�W�=(����k�=HDG>��>����z��ɠ�΀ �U�g>��m>u�r>>�M>ű�?6o,?�K?"��}�oS[���=��iT��OսJ@�>rl�>p*F>��ܾĽ�ni^��O��J�9o߽�SU��=|,>�s>FR}>nOa=���Cm�<."�~�E��1=B;�=-��>:��>��>̎S>W	=hܾ����VR?�T�������@�K����>�`�b'�<b�����>�u=銿�*��cf�m?�'�?��?��Q?��ͻ��=Έ�=�U=���=\c7�Xi羾9���>��?G�>y���h��aj�=���>+1�>��ǽ
���ܾ*�ֽh���'F�Euf=K˾���:�"����󑰾�	F�^쾶�;��ӏ��G��53Y���e�g�����ž�ܨ�t��?�o�?�5�>ɂ������u �5���Zt�=�#�/���y������j¾�-۾_��2�,�MU+�@g;�:8Ǿ��>��X��R����|��c(��-��d6>>�h.?�_Ⱦ�c��Y��#�a=#>L-�<���6�������� ��W?O
:?L��S����-�T�>�W?/��>,�#>����潌��>!�3?��,?m���������q��4Z�? ��?�K?o�(�-F��l�~�����	?�?q{6?�᪽���ʛ�*��>�`?*�?(��Oみ��-��`�>�;�>�A��Τ>�J�>�d
>՟=H�ϟ����|�>\v�=�����F��w��u�s�� P>�U�>M��=~IT�����G�>j� � VվH�9�����a��R�=� �>j"�X�7>J����>��a.�;ɉ�vkZ�ؒ��TTm?jʣ?�xS?�g?����<�幠��5�"'?lt�>�>3 ��{�>8}?Z���	O�;㈾�o/?3��?L��?�1�>��P�1�̿U��Kɉ�oYܾ
��<_ͼ��A>���]�=�<>�����C=�{=G>�[>A4>L�+>�b>�)></��=�.�D�������&�r�e�:�a�������6u;�~��L��ֶ����۽l%������zw�ɖ��ݢ�n���M��=��V?l�>2�9>��;��
=>�w����˾Ϟ���_��� ����9��==�k5=A�9=vE>�tܾ�	?���=���=�M�>��y�r�=�I�>	΁>Yy)���=>�~ >c:Z>*�>��?�G�>��=�'�>�[�=�H�����` ,� !0��� �N�E?gP�
ƒ���'��hپӯ��~N�>�
?��O>��+��ʐ�C�y��Q�>$½�E�X�x���� ��>ѽ�>���=8:���l�D���pAý���=*X�>��=�Ô��n���u���<���>��; ǔ>��>x��>�Yo?��$?��<���>pf>j�=�-=��">2�@>c&�>�?(�Y?�2?���>�S>���r�=�.>Bƛ�s������n 8>�=L��=�=ui�U
�����Ȏq>�C�>z_p>�mO=G�|�ά�>Kk8?%��>]��>�6�c�<���L�~���Y>4'�k3�>I��>��?���>�f�>�C5>͗o��#��*o侞	�>�YG>]�bv��:��Ju>�ah>#~N?��0?hC�-\����<G��=�Y�>a`?i)?�-�>2>����c��N�ֿwy �Z�!���U�ƻþ��,�0慾-z|<Q�!>3]����\��ɳ�|a)>��]>V�0>jN�=UH콌2�= :�>X��>_�V<'�}>	>|�=\Id����=uG�z�^����:^HԼa�d;q�o=5��;� <*�l;Ź�~$?���>ӿ�<rz=0�׾m��g��=`�;?��v>���>.�??�>!����e��z�cG����?�	�?���>��J=�	�=�<���r��?t<�>Aѱ>��>qdU�F}��T��>�`?�C?��>OvܾkI��X����̾bi�>X.=i	��Ù?��_?����-���;�LG�i+�`��<Ш���Y�9�����%�N�9�5��](���*Y�g�=���>?J�?}d^��z�=	ɲ��ݖ��������X;=�=���>�6>+&-�v�����,gѾ;�:�%�&=~�>�u�{e?l�>��/?fpy?��z>6�:�"$���j�?���>���>��>�s>���>l$�;�T�?�=̬���E�	���.����g<��ܽUܼK�=7�F>6j�2ۄ<=�>�Q��[K�*��<��<1D=3R��>�̓>�(>�?*�:?qXվ�M��K�f>:;��Pt�l	�>ժɽ��.=���=1��>��m>��>��
?][L>��:��˾��<Z�����G`>:G�>��e?"KM>MO���>T.�FǾf��=Kv=w%�8���Ѿ�/���\�Yx�> �=]�]>׭�=hܔ?V�>�qT?8d�>��Ͼ*�y����>>��S����>��?�>���x"�G���T������~刾�?�<t�j>��=Í�>igh=����~�|>�e<��?�����>�B>���>�}$>59!=�z�
���^8I?��"��_���J;�.��>�-�>��<V�v��2?�0k��Z�������b߾�oJ?ì�?s!�?��.?b��ҕ-;��=l�I�y�>�j�=W0�<��`���6���?>*��=�f�=�}��T%�;�q�>�A�=Ц�<l�"��~��������}a6�;39����>{��E����\$�V��̮��}H�R@/��@���Z���Ͻ�C1��^���1����A�`��?��?���>풼�Z�7�Xľ��[����
|��w�8_���2��(�����̾Dn޾����Eо�N�>b����f����|��
��14>&��=r?f�ξ@B\�]�!���0�b�>3��>{WS���d��4���s\��D?��-?������v����d=��>J�>�]�>��6�����wG=%�h?�"k?�g�=�������3���%`�?�W�?�2H?/z-�P)J��0��Ү���#?�43?"�%?��}��5�й�����>�&x?��-?�;P�v�i�9�Y����>��^?1���z��>�K�>h��=�q���B����!dx�}P9�7i�=��w��y�a���T��(ŗ>�|�>뜰;\mʾ/�����v=n��7[�e/��h�����)^-��n:<�� �9>h#����=TK�Qꏿ�n�����.�?M,�?�8%?��i?�2��E�p�{l�;�>��4>��>�s콗R�>�M|>X-���
ܲ�Y�I?U�?�X�?-P?؞R�_�Կ3���e�������=��W=s�>`m��">\��=���}��q� >
u�>�(A>�bg>�B>jj$>�>迆�(��c������c�J��������N����
�\�^�������������ݽE���@ ����d�S37���s��<�5�>���>��?f Z>����*��<׾�;ܾЁǾ����/�;�޾~��Gþu4���b^Y��T-�!5�7����?y$g���.>R8>�6��~��Qz>�C��'��>��L=?�=j�>=>�\�>iE�>-�>yb�>��0<����������`���zN�,2?׈�A�\�՚��X��B����Y�>�`?q�V>�,�pg��9r�&��>�����F��-!��h��y�>��>�=U��;�����i��/�[�>�Ͱ>@`�= P@�㮌����w��0X�>N����>'��=��>�vn?�G?�}x���>0n">2��=���p�`>]<�>���>�\?�w0?ʝ?3* ?P#>O�j�<��=���<M}�0,"�N�B���x=]Ts<�Gڻ��I�&[���p=�>�=�S�=�f_<��>cv=��>�Q#?Xk�>Z��>2o�j�6�$_?�����~>o��?t�>ZS�>���>�?���>?GS>��V<�i��3����O�>�8>7{Z�n�l��ǈ��+>�j�>�-W?�<?ޖ!=c�5��}���6(=_ƍ>��?:b<?�e�>��>Tý���lӿ_$�?�!�����O�AԈ;��<�C�M���7��-�-���r��<��\>i�>6�p>/E>J�>z=3>�R�>�GG>�҄=w�=82�;�b;��E�ޗM=]�yDG<R�P�疯�*ƼE���c����I��>��7��8ټ4�?	b�>��(=���=P��Z(���=��>��u>�K=?�Q�>���="ғ���c���^��;�����>Ō?��>��<�~�=�����彙�?��?֑�>>��������'] ?�?BJe?���>�Ӿ����lZ�Y6�O5?�6=,��`�?�_?���񭇾ȗ���B����I�k=���Z�ޑ����%�S�6����<���R�+_�=V��>�?4⁾��^=��(���g���ᦾ`D9=_�=W��>B>����̛�(��<�Ծ"X��>E=!�>p�����?^3�>��7?USq?�f>HL>>�>��?�{����>�>�?�>�N�>��Z>��
>s�
>o1^�c��6"9�0Ǿ
l<չ�P)P=���=Ұ0>rD�=r��=߽�=��;Zk2��눼�.�=9c=	���L�=���=
��=5��>��&?����창�>"#ս��"�u�>e�H��e����f>�&U>�[S>�E�>���>�ؔ>��6��s�[�X����[�7>� �>	�Z?3U>����=Ny��G׾��=0��Pm<&�j���վ��G޼�0��>�6>^�>��=�ك?� ?=U?��
=��6�"%m�i:�W�1�1C6;^
�>�1�>���=��޾�I&�1[W�^O_�g9H�&J�������6>@KL>��\>:g>w�=nu�=����Ȇ=?-�^=��;��B>��p>���>�=>@��=|C�s��ˑB?��aM{�p��%����伵��>1�$>���>�n\?���5���G
�������3?���?���?���>aǸ�Z��=u���Lq�ץ>�=#>�v�=�|�,�����>�&�>��R=�ƅ��QG1>��>�=��>`����n��{ӿ��5��f<�ם��֌�֭ �|�޾(���;n��0�}�R���6�t�����G�@̈́�J�r�����i߄�	2��i�?�r? ��>��=�L�iS�c:+���v�޾u�Q�|"�����Ҿ��� �B7��M]�/,��QG��36�>vc��S~���cm������>�'H>~?��l�����:�s�˽���>l�h>ڒ�{y��<�������3O?��'?��ƾ)�۾{�E�cU^=�ɿ>�p�>��>�Rl��!���xo>�L???H?c��=zҒ��a��1뼳��?eǸ?V�9?���e):�Ǹ��fҼ�nE?�l�>P�!?�4Q�L�����=��>cc?��.?�抾�X��^S8���>��a?�q���u ?̐�>��><�~��d瑾�d����!��%�C?@��J=i����Ӭ������*>�%j>����;S׾#����}>y�ھ�v޼2+j�����#����*>�i>���Ӹf>Ȅ�0n$=�]c�=�)�W���*�`n?�~�?;D?nu?�S��G�� �.�U�`#?��>LH>�V�<�*?���>�AܾV�L��ӾR`c?���?��?�?�D�5�ƿ/퍿6S����p�|��=�����>�z,�\�J>�VD>�iD���=�!�=.J>>q�Z>j�>;y=�>�S�5�,�<ܕ��Յ��mF������$�:���s���9@�����*�����M'*��s����>����쏾���P��7w>T�?Ƭ�>h��>@�=�3�=ͥ��۾x������U�����Lr�2���I���F ����SY��������	?o�����=nź>y�=>A>�q>���=O�>��>>��=h�>�3>��*>8�v>[V�>��%>>'�>z��=)Ć�������k@��oG��PJ?ʕ>��f��9'�n2㾙ؕ�P9�>ם ?�C>��7�:����0y�|.�>�a���A�>WD�qV���A�>�ϼ>p�:= .׽k>�;;�f�'�ɽX��=�id>s�
>k�m=:�.�6��1���d�>,�Ⱦ��K>��I>�[�>�v?�0*?+RU=A�>�TY>�� >��9<1>�r�>S��>�P�>Q�<?S\?�r?��%>"���{.>�]>�D޽!΃�4�p�<	�z��������=�+T=#N=m]>`�G>Heu<[���V<�-�?b�>��?���>聞��6�_{�P3�=>Q�>C{�#�=>��1>�K�>ee?{?��>�M$=���Mr9�x�>�_d=��q�~{�9�&�z��;�2�>�Ml?�A]?����-d��R$�,����g =ޓ�>�PO?��m>��>M�3� ��!��Es���Ⱦݩ]�doӾ����%��)J1��gU��)��}�>�#�<q�=�
>�C,>3r�=}�B�򦽾��>�hv>��=�<y�ȼiW��y�;�l�=;ɫ����xE\����u�2=�:����_ѼH6<
��;B�?Ø?#m>y5�=*�˾�{?7�R�>d��>�5?��>,b����i���a5�؝r</?.d�?�q�>�5���0>w�^��D��i�>�F�>;�>jj,>�~���;��4�>8�?�|[?�%�>t#뾏�]��hv������k�>���<\/��Ԝ?^[M?�����H���F�Q��l��4��$m��඾&���0���������C�T� >��?��?��̽���=�ޢ�i\���9s�փ��>�<���<���>��E>Uqb�@���"�����A�!��N?=�G�>���p|*?$0?��6?�]�?��>�O>� e���>lOL��>�_�>H��>��>��>�
�=|�=7y���pe���-�mv��g=!q4�zX�=�>��m>ku�=D��=�q�=�-�;W׽��w�'��=��=+9P=��=���>R[�>�?��'?�����<�z>�]�=L	#=�G�>k����.�hp>6�=�G�>$��>"c�>�k�>�`��]|�Z3����k�>�W�>�i?�y_>x!=]7&>d�=�����w>r��X��<%���[���F�����>į�>.�3>5�=q̛?p��>�(�?ߩ�>�����~������¬��@�R�>��;?��V>wѾ�'��J1��rA�>o��<�8\��g>�I>�a�=&�O>���a*��MM��]w>4�:g���ӳ�ـ�=5r�>/�>Kv_=3,q=�膾&����hQ?@��y����Ͼ�x�P^>��f>��P�J��>��?z������|���$��`A?�'�?��?�'?QnｑO;�~2�=�䇼���>�T>CM=/n�ɓ¾j2o=��*>��+�嵖���C>��>�?/>1t
�(����S����칿S�B�5������2}���M�,����U�<�����O���w.k��D��/��j�!�J�C�7:���ɛ�E���˷�?�e�?�H�>j?�� �@��$r����<�ʠ�Bf;��
�m�V��3˾@���M�cS��1�0���'/����>s������N�a������o>S�>	?9���n�n�~�����KL�>��
>,�̾�)m�lЂ�
��=:X?�&?D��9���[�4�M>�Q?�7�>�N�>���l���>/�K?��o?/��>Փ�m����{�9��?���?>�??�N����I�f&� �`=��.?IL/?B$2?�lU=��$��� >b^>�e?>3?����� ���!P����>$�o?=*G�|>KU�>m�=	���қ��W���:?��IN>E��=N��;�ž����s�@>�wq>,��=/8뾤���H�>��ɾ�S��DY��c���.�.��<`�?$h��&>��j>6�a>Y�/��ˊ�)��gݹ�x&M?���?Ռ=?`|-?��ھ�kҾA�l�`f�=2�>�%�>*=®��q�>�>�F۾�Hi��'���?L��?�l�?�!J?y-h�_�˿lo���]��>ش�|��=ϸ�=ĔL>W�ὠ̣=�}+=�<;0M<�	>��>ja;>�Za>��3>$�;>k�T>������(��t��e���W�M����9��c�`�
�n7y�2��ƻվAY���uT�8����G�>�7]�����`�5���C>LC?�{?o��>���>���>���o>ܾ��A�cm���o��͜��؏�\�Ѿ�_��4�Խn�{��%������	��8�>�q��qso>z�>C�4��d�=��>�C:jq�=R��=L_>Θ�>��>j�>��%=�>y=�>EFd�♋�?�T�-��#�u<T�r>�l1?p��������i=�Y�ɾҩ+>��&?~I�=bDK�<����;s�[�>WT۽'F����V���P�O�=�g�>o�{>�1���=ZD�=����/>/>&��9����� ��h>�?�>���yi�=��>3?�Ry?9�9?؋�<�H�>�?>7v�>�
�=�Ct>�JY>V�Y>X�>	"?=?���>�M�=H:|�����G�;�x!��Q���}��A;����s% �������=��s<f@�NF�=�$b=w� �D��u\(<c~�>��D?]�?`?b%��vJ�܌�����}fr>�8̾���>�g>�z<t��>�J#?���>�ƺ=���� ���K�>D�G>O�j��F��HJžgT >��F>�b?<�?�f�� O�l�ٽ��>�B�=WC�>}�?�ԅ>��Z>�>������T�)�#���z�����=c�l�P�<"OB=�IQ��S���1=���> �=��$��զ>��>C�M>�<�>Am>�l�=�T>�>�=USU=^|��u��ת�FC���;���;>pt=���<�z�=<���Uk@�i�a;)�/��>�?}(ڽ�&]����lc��d���4?��_>O��>�-�>�>�*��� �P�,��>����?�,h?Ooy>���(3���
��8>ɽ�>�J�>s_>�YG;�W<�v������#?�?pk�>�C���u�-�B�����>�.V�LЙ��Z�?�Ob?�}��ֳ��suQ�]�C���.�d�C<��T�I�W���
��7��;���8���TԾ'W��U�2>���>��?D��=��e>����d���Z������S���B�B?V&�<K���)yK� n����=Q�N>�<w>hG|>~P!>%r�>�+?��4?KX?r�$?��	?�c}���>�E&�h�>o2�>�N?�
?��	>�����>@�����\�S��I����3�<f�y>Ǫj>G�>ud�P� =5�3=F>ٖ��������=�Q�=cb6�cV
����^@���?��"?�=!�@>��q��4��N���uw�N3>��4>�D��@����B>�s=�6?י?7[��*V�"�+�q��J�L����>�?�u>��^��O�>b��Lڹl��CT�=�3���G���Y���
��N�=)J�>0o���>�v?\$L?�)?(>�����!GV���(���@==�p�O�">��~>�,>C���W���L�� T�C ���2�=G������y=>�l>���=�;>qf=��%�σ�ds>�s��9>�3�>��>�T�=h6�=��T���4�E?��<���4���7���'�z�5�f�>��=�h+?�6����,�)��[
o�9�d>ӥ�?�G�?Hw?X����=��=��<G�n>0�p>ʭT>��Ž��;>z�l�������>IM�}���L�>q��=��>B��ాE/��������P�Y��y���E�s�7���۾��}%/��Jr�l��h���E���PD�ϖ��E��M��-踾3I��:-����?�?h�>���=ut�����
��=@#��}�f4��n:~��yǾӸƾ`�⾏��A9�p�;�;�曦>�S"�����啀�ՇH�i�q�4>T*]?CS������������~�D�=:�>	&о�xp�܅���<>	�?0L?A�����>�����q�6!>?a��>��>�wӾ˭<��=� <?�]8?��I=���S��U��=�Z�?,��?�'?ғ��1g�D�?����=��<?h�5?Ct?�<��m����&>YMG?�?BF�=x� ��bg�IM'�z4�=f��>�N��B�>��> �6>q�ϽύŽ�,�]����>U>�Q�>2���Gt=y��������B�>N��=�욾ˁ9�Wʏ>C,��WN��|O�w��/���=v�?������=��z>I>�+�R�yy���m�8�N?#�?KMS?�r7?`����Ȕ��!ob=Dq�>�]�>S�=]-���>+�>�C��r��y�� ?<	�?-�?�
]?�%h��ܿ1����EҾ�.̾���=PV�=FkX>����f=fl3=x\:��э�F=�j>d�>G�/>�7L>�cx>�!g>P���|+��2��4V����O��$���׈2�yp��蛾d�������ڿ��Z����������?���������?p�3�<��>���>;d�>�N�> �o>Ť��k|��5�ֽ�>�B���5��7H������/�����f�N�`���}�i 	�೮>B�;m >Ll�>��$��=J>��>����.�> >=�P��gk>m/�=T_�=Rv�=R�d>z��=@p�>��8>�Ԅ��Zf�0'
�Lֽ�z>H�'?�%�`F�L���6_�H+���;��?�Ul>@�1����J����>�����̖���I��?��|�>���>��=6���'b�0��!��=�R�>���>�m�=c7D�Lv��L�u�U
&>k��>7b�:&��3�=�}&?x��?�S7?��S>���>�1�>���>���>ݱ1>2�>=�y>���>�8�>�N�>Mz>r�>�T��x[=�E>����p�>q&߼���<mJ�<5�n)������7:!�̽,p#��;!��=���-�<�(�>�dA?���>�?����Q�a<`��+�����<�1ɾmBP>�q<>�<�=��g>3�?��>s��=�<u�K����v�>c[�>B�v�ģ���k��{k*>o��>��P?��N?��>۸��p��L\>�3��$i=!T?.��>`b���w=�a��BֿXH'�j@0�x����6���=��z��������B꽷�-����=���=-�E>O�X>3�,>z�\>���>��S>�L�=�w�=�������;�:����<g`G�A��<��9p��<�?���[$�����6��<�=ҫ=~����Z?`Q?�~!��	�~<�����d��u��>xӸ>�+?�>k�7=�z�,G�:QA�n��"�?��c?���>2R����=�>:<(<���>�R�>�>����������� ڻ��>)?[)v>3���E�H�@|f���� �>0�-�c�ڽ�f�?go?8U��:�����@��,��P��`��E�=��s��{���F������+f����g=��=Y| ?�ʫ?� ��/>bƃ�ⷫ����e���kf���r����>�Vt>�'���y��j��і���|�=�X>��>6�>	aZ>�>j�?xMZ?ֹ ?��?n:Q�#,�>}]>ֻ>�Ğ>���>�?-�>�8w�h,�<�\ֽ���������=�2�na�F>i�>1��=���a=��=��<��
��:�kw�=���x��q�=*$>�ܤ=�+�>�!=?�V�=��B=}i�e����+ڽK�佌��>�ֽ���1�>}��>��>���>��>\D7>UzǾ�qֽ�-�F+����
?zo(?:��>�I�=��?>�H�)O�7滉��>M�"�l�"��'�8��<�d��5;�G�=B��>1�u>��y?��>?A]/?����'�R^��G6���<�y��\Bb>�V�>��}=B砾���C�Z��qO���7��&s=|K����2��=a�;>�T>���=�wg>=�<�/��vý�8>�M��#�>W�>�u?��=�d�;bℾ&	��P?�|��E���#�y�i�h����>b�*?��Z?�Ջ�Fǖ��ћ��Л�lR.�mG�?؄�?�2�?+�����y}>���=�k+����=��r�/!>3��*�>���>Km�-�߽-�>��z=WaS=~@���M��8Mj���оS�ӿ�,l�5��R�/~�����Pp�����R[�9�C��A��^��3fо����ڴ���<���CT�v��2�� ��?� �?3��>�Gz>:	#��x'�²,�����]!���K�C�A�[<�gԽ8 ��� ��������N�����W��O�>�k��㑿%H~� v&��SG��PE>��.?��žs��������l=+<>���;������!���u	���V?
-9?W羼���X6�GQ>�U
?��>�� >������콇��>ku4?J*?:I6�I���H��q�;m��?O�?�!?��پ�d��}���0>��/?B}%?/�>s#�Ž���=K�?��3?�M�>�V����.�;�R��=2�?9	 ����=��>��D>g�߽ԭQ�Si���_%�ጻ1_>�\�=��*�	�P���5�V>�5�>��z<���ޏ�Wʏ>C,��WN��|O�w��/���=v�?������=��z>I>�+�R�yy���m�8�N?#�?KMS?�r7?`����Ȕ��!ob=Dq�>�]�>S�=]-���>+�>�C��r��y�� ?<	�?-�?�
]?�%h��ܿ1����EҾ�.̾���=PV�=FkX>����f=fl3=x\:��э�F=�j>d�>G�/>�7L>�cx>�!g>P���|+��2��4V����O��$���׈2�yp��蛾d�������ڿ��Z����������?���������?p�3�<��>���>;d�>�N�> �o>Ť��k|��5�ֽ�>�B���5��7H������/�����f�N�`���}�i 	�೮>B�;m >Ll�>��$��=J>��>����.�> >=�P��gk>m/�=T_�=Rv�=R�d>z��=@p�>��8>�Ԅ��Zf�0'
�Lֽ�z>H�'?�%�`F�L���6_�H+���;��?�Ul>@�1����J����>�����̖���I��?��|�>���>��=6���'b�0��!��=�R�>���>�m�=c7D�Lv��L�u�U
&>k��>7b�:&��3�=�}&?x��?�S7?��S>���>�1�>���>���>ݱ1>2�>=�y>���>�8�>�N�>Mz>r�>�T��x[=�E>����p�>q&߼���<mJ�<5�n)������7:!�̽,p#��;!��=���-�<�(�>�dA?���>�?����Q�a<`��+�����<�1ɾmBP>�q<>�<�=��g>3�?��>s��=�<u�K����v�>c[�>B�v�ģ���k��{k*>o��>��P?��N?��>۸��p��L\>�3��$i=!T?.��>`b���w=�a��BֿXH'�j@0�x����6���=��z��������B꽷�-����=���=-�E>O�X>3�,>z�\>���>��S>�L�=�w�=�������;�:����<g`G�A��<��9p��<�?���[$�����6��<�=ҫ=~����Z?`Q?�~!��	�~<�����d��u��>xӸ>�+?�>k�7=�z�,G�:QA�n��"�?��c?���>2R����=�>:<(<���>�R�>�>����������� ڻ��>)?[)v>3���E�H�@|f���� �>0�-�c�ڽ�f�?go?8U��:�����@��,��P��`��E�=��s��{���F������+f����g=��=Y| ?�ʫ?� ��/>bƃ�ⷫ����e���kf���r����>�Vt>�'���y��j��і���|�=�X>��>6�>	aZ>�>j�?xMZ?ֹ ?��?n:Q�#,�>}]>ֻ>�Ğ>���>�?-�>�8w�h,�<�\ֽ���������=�2�na�F>i�>1��=���a=��=��<��
��:�kw�=���x��q�=*$>�ܤ=�+�>�!=?�V�=��B=}i�e����+ڽK�佌��>�ֽ���1�>}��>��>���>��>\D7>UzǾ�qֽ�-�F+����
?zo(?:��>�I�=��?>�H�)O�7滉��>M�"�l�"��'�8��<�d��5;�G�=B��>1�u>��y?��>?A]/?����'�R^��G6���<�y��\Bb>�V�>��}=B砾���C�Z��qO���7��&s=|K����2��=a�;>�T>���=�wg>=�<�/��vý�8>�M��#�>W�>�u?��=�d�;bℾ&	��P?�|��E���#�y�i�h����>b�*?��Z?�Ջ�Fǖ��ћ��Л�lR.�mG�?؄�?�2�?+�����y}>���=�k+����=��r�/!>3��*�>���>Km�-�߽-�>��z=WaS=~@���M��8Mj���оS�ӿ�,l�5��R�/~�����Pp�����R[�9�C��A��^��3fо����ڴ���<���CT�v��2�� ��?� �?3��>�Gz>:	#��x'�²,�����]!���K�C�A�[<�gԽ8 ��� ��������N�����W��O�>�k��㑿%H~� v&��SG��PE>��.?��žs��������l=+<>���;������!���u	���V?
-9?W羼���X6�GQ>�U
?��>�� >������콇��>ku4?J*?:I6�I���H��q�;m��?O�?�!?��پ�d��}���0>��/?B}%?/�>s#�Ž���=K�?��3?�M�>�V����.�;�R��=2�?9	 ����=��>��D>g�߽ԭQ�Si���_%�ጻ1_>�\�=��*�	�P���5�V>�5�>��z<���ޏ��H�>��ɾ�S��DY��c���.�.��<`�?$h��&>��j>6�a>Y�/��ˊ�)��gݹ�x&M?���?Ռ=?`|-?��ھ�kҾA�l�`f�=2�>�%�>*=®��q�>�>�F۾�Hi��'���?L��?�l�?�!J?y-h�_�˿lo���]��>ش�|��=ϸ�=ĔL>W�ὠ̣=�}+=�<;0M<�	>��>ja;>�Za>��3>$�;>k�T>������(��t��e���W�M����9��c�`�
�n7y�2��ƻվAY���uT�8����G�>�7]�����`�5���C>LC?�{?o��>���>���>���o>ܾ��A�cm���o��͜��؏�\�Ѿ�_��4�Խn�{��%������	��8�>�q��qso>z�>C�4��d�=��>�C:jq�=R��=L_>Θ�>��>j�>��%=�>y=�>EFd�♋�?�T�-��#�u<T�r>�l1?p��������i=�Y�ɾҩ+>��&?~I�=bDK�<����;s�[�>WT۽'F����V���P�O�=�g�>o�{>�1���=ZD�=����/>/>&��9����� ��h>�?�>���yi�=��>3?�Ry?9�9?؋�<�H�>�?>7v�>�
�=�Ct>�JY>V�Y>X�>	"?=?���>�M�=H:|�����G�;�x!��Q���}��A;����s% �������=��s<f@�NF�=�$b=w� �D��u\(<c~�>��D?]�?`?b%��vJ�܌�����}fr>�8̾���>�g>�z<t��>�J#?���>�ƺ=���� ���K�>D�G>O�j��F��HJžgT >��F>�b?<�?�f�� O�l�ٽ��>�B�=WC�>}�?�ԅ>��Z>�>������T�)�#���z�����=c�l�P�<"OB=�IQ��S���1=���> �=��$��զ>��>C�M>�<�>Am>�l�=�T>�>�=USU=^|��u��ת�FC���;���;>pt=���<�z�=<���Uk@�i�a;)�/��>�?}(ڽ�&]����lc��d���4?��_>O��>�-�>�>�*��� �P�,��>����?�,h?Ooy>���(3���
��8>ɽ�>�J�>s_>�YG;�W<�v������#?�?pk�>�C���u�-�B�����>�.V�LЙ��Z�?�Ob?�}��ֳ��suQ�]�C���.�d�C<��T�I�W���
��7��;���8���TԾ'W��U�2>���>��?D��=��e>����d���Z������S���B�B?V&�<K���)yK� n����=Q�N>�<w>hG|>~P!>%r�>�+?��4?KX?r�$?��	?�c}���>�E&�h�>o2�>�N?�
?��	>�����>@�����\�S��I����3�<f�y>Ǫj>G�>ud�P� =5�3=F>ٖ��������=�Q�=cb6�cV
����^@���?��"?�=!�@>��q��4��N���uw�N3>��4>�D��@����B>�s=�6?י?7[��*V�"�+�q��J�L����>�?�u>��^��O�>b��Lڹl��CT�=�3���G���Y���
��N�=)J�>0o���>�v?\$L?�)?(>�����!GV���(���@==�p�O�">��~>�,>C���W���L�� T�C ���2�=G������y=>�l>���=�;>qf=��%�σ�ds>�s��9>�3�>��>�T�=h6�=��T���4�E?��<���4���7���'�z�5�f�>��=�h+?�6����,�)��[
o�9�d>ӥ�?�G�?Hw?X����=��=��<G�n>0�p>ʭT>��Ž��;>z�l�������>IM�}���L�>q��=��>B��ాE/��������P�Y��y���E�s�7���۾��}%/��Jr�l��h���E���PD�ϖ��E��M��-踾3I��:-����?�?h�>���=ut�����
��=@#��}�f4��n:~��yǾӸƾ`�⾏��A9�p�;�;�曦>�S"�����啀�ՇH�i�q�4>T*]?CS������������~�D�=:�>	&о�xp�܅���<>	�?0L?A�����>�����q�6!>?a��>��>�wӾ˭<��=� <?�]8?��I=���S��U��=�Z�?,��?�'?ғ��1g�D�?����=��<?h�5?Ct?�<��m����&>YMG?�?BF�=x� ��bg�IM'�z4�=f��>�N��B�>��> �6>q�ϽύŽ�,�]����>U>�Q�>2���Gt=y��������B�>N��=�욾ˁ9�Wʏ>C,��WN��|O�w��/���=v�?������=��z>I>�+�R�yy���m�8�N?#�?KMS?�r7?`����Ȕ��!ob=Dq�>�]�>S�=]-���>+�>�C��r��y�� ?<	�?-�?�
]?�%h��ܿ1����EҾ�.̾���=PV�=FkX>����f=fl3=x\:��э�F=�j>d�>G�/>�7L>�cx>�!g>P���|+��2��4V����O��$���׈2�yp��蛾d�������ڿ��Z����������?���������?p�3�<��>���>;d�>�N�> �o>Ť��k|��5�ֽ�>�B���5��7H������/�����f�N�`���}�i 	�೮>B�;m >Ll�>��$��=J>��>����.�> >=�P��gk>m/�=T_�=Rv�=R�d>z��=@p�>��8>�Ԅ��Zf�0'
�Lֽ�z>H�'?�%�`F�L���6_�H+���;��?�Ul>@�1����J����>�����̖���I��?��|�>���>��=6���'b�0��!��=�R�>���>�m�=c7D�Lv��L�u�U
&>k��>7b�:&��3�=�}&?x��?�S7?��S>���>�1�>���>���>ݱ1>2�>=�y>���>�8�>�N�>Mz>r�>�T��x[=�E>����p�>q&߼���<mJ�<5�n)������7:!�̽,p#��;!��=���-�<�(�>�dA?���>�?����Q�a<`��+�����<�1ɾmBP>�q<>�<�=��g>3�?��>s��=�<u�K����v�>c[�>B�v�ģ���k��{k*>o��>��P?��N?��>۸��p��L\>�3��$i=!T?.��>`b���w=�a��BֿXH'�j@0�x����6���=��z��������B꽷�-����=���=-�E>O�X>3�,>z�\>���>��S>�L�=�w�=�������;�:����<g`G�A��<��9p��<�?���[$�����6��<�=ҫ=~����Z?`Q?�~!��	�~<�����d��u��>xӸ>�+?�>k�7=�z�,G�:QA�n��"�?��c?���>2R����=�>:<(<���>�R�>�>����������� ڻ��>)?[)v>3���E�H�@|f���� �>0�-�c�ڽ�f�?go?8U��:�����@��,��P��`��E�=��s��{���F������+f����g=��=Y| ?�ʫ?� ��/>bƃ�ⷫ����e���kf���r����>�Vt>�'���y��j��і���|�=�X>��>6�>	aZ>�>j�?xMZ?ֹ ?��?n:Q�#,�>}]>ֻ>�Ğ>���>�?-�>�8w�h,�<�\ֽ���������=�2�na�F>i�>1��=���a=��=��<��
��:�kw�=���x��q�=*$>�ܤ=�+�>�!=?�V�=��B=}i�e����+ڽK�佌��>�ֽ���1�>}��>��>���>��>\D7>UzǾ�qֽ�-�F+����
?zo(?:��>�I�=��?>�H�)O�7滉��>M�"�l�"��'�8��<�d��5;�G�=B��>1�u>��y?��>?A]/?����'�R^��G6���<�y��\Bb>�V�>��}=B砾���C�Z��qO���7��&s=|K����2��=a�;>�T>���=�wg>=�<�/��vý�8>�M��#�>W�>�u?��=�d�;bℾ&	��P?�|��E���#�y�i�h����>b�*?��Z?�Ջ�Fǖ��ћ��Л�lR.�mG�?؄�?�2�?+�����y}>���=�k+����=��r�/!>3��*�>���>Km�-�߽-�>��z=WaS=~@���M��8Mj���оS�ӿ�,l�5��R�/~�����Pp�����R[�9�C��A��^��3fо����ڴ���<���CT�v��2�� ��?� �?3��>�Gz>:	#��x'�²,�����]!���K�C�A�[<�gԽ8 ��� ��������N�����W��O�>�k��㑿%H~� v&��SG��PE>��.?��žs��������l=+<>���;������!���u	���V?
-9?W羼���X6�GQ>�U
?��>�� >������콇��>ku4?J*?:I6�I���H��q�;m��?O�?�!?��پ�d��}���0>��/?B}%?/�>s#�Ž���=K�?��3?�M�>�V����.�;�R��=2�?9	 ����=��>��D>g�߽ԭQ�Si���_%�ጻ1_>�\�=��*�	�P���5�V>�5�>��z<���ޏ�/��=m��ؖ����^��ܾ� ��[=��p>�"�?޹=���>��4>:	ܾ�?r�6,��8F����P?�? [2?��%?����q�,��qC߼��(>�ф>x�=E�*�u�:>1��>�`�����E�jU�>���?m#�?]@@?3m[���Ŀ˵��̀��򾎰��f5>��>�^�<SDy=�	Խ�;�=��d=���=�g�>�%�=<RO>�Jj>'Q>g�>�����-��ӈ�V����f���Q�a�*DI��0(�U���R9羢�~�����L�A�b�H��������<vH�R��5	>�m?v�1?���>���>��>�,<���̾5I��I�B�I��k��ھ�2�$���B�������Z��p��<~�Q!�>y���=�M�>
 >�z>E;�>�+�=7�5>�ɽ���=�F>�5>�y�>�o5���=�|�>��9>&��=�P����i���=��ð�.~��,�=?pt�Ryt�)"1������p0���w>io�>t�>���e��@���֋�>z��2e�ӑL��%1=i>Bھ> k�=��u<�F�;V� ���<:	=���>�'#>�e�v�J��>;��� >H�>.ː���>�v�>V:7?km?��;?�8e����>Bp�>yL�>;]!��緽��,<�e�>:��>��>�7!?[dH?�l=^���.
{>�Um=�t��q��Vg�/g�='S��a�A�Ҽ?��<z�y=�[<�]:;J
�i���8\i=eŬ�i��>�K?0A�>�?�>��j���B��M��'=�/(>J��<�����b>�~*>��>��>�F�>�ꀾ>n'��H
�xB�>��>�(8��4P�����6�U��(>7sE?�f)?� }>I.��G0��>����>lTU?�B�>���=ZEڽ�X���ҿK�*�n�$��֝�,�,���:-]c��N����(��۽X�<��S>2�d>g�X>�Ma>k7>ؼ#>Vs�>��F>���=�=����qj���a�@zJ=�f���KN�E*?��r�<R �U�\�n�di�x�Լ����?%�T?f�?e��?������P�� W
�ڐ�>&��>�?��?�t<�� ���P��:�X������>�?E?�e?Sn=�s2,=گ�<�>��>��>��&>�7��K�`�p#H>�k�>�"
?��^>�b���^���Y���4e�>ʥ���&<>r?^�-?аھ��뾮*1��';�g������r��x��M�Y�]���o��vH�Ԙ�a�k���Ƚ�!?�ϩ?�T��Ri=�3��,���_��HBþ�a�>���>@�<
��>�L�$[�=��-s����A�j��%���R>���>��*?���>S�C?�.?q��>ػ��+?�V8����>? 7>`�>�ۚ>q�> ��>A>jy�=��h=���[����=��=<>|ռ>���>��=�=#R]=���=�5��?�<�ms��g����2=-���(�;a� >��?��2?��G;�ּ9�P�Ug�.�Z�vӯ>�	?v�t=�3Ծ�i��R�+��->�N?f��>U*�=��從�w�l���ݽ}P?��#?�>U�>+�>;���?�����l�>�K�<Mľ��i�m�����:J>ݓ[>��>�ǈ>4e?(*?��?�y���Q�(�x��n��ʓ����>�?��=M���ݪϾyE��K��M�Sv��9ǽ9U�=w�\>���=R>ݮ=`}�=>@I>��<����9G�R�>�X>���>��?�v>Ԡ;��;����Ͼ��I?EM���z�ᒢ�s2Ӿh�0�f�>�H>$�Ľxo?p����������<���>o�?iS�?�&`?F*?�Z��hY>��X>��>�A�;#�3�9޼���!�3>�o�=��n�=-����$�F^>��n>}ٽ�ľ\�޾�K���̿�i��溾����n���U���9���'�����8I3�ZW�b��+�=�>Ȩ̾�)��O�%)�}xݾ��\?#Z]?@�8�|=�0$��X��O���@ ���rV��Ml��S�+Z��.[��%f�hM��	���#��z徴�}�?�C3��5��ZA�[v=��W>��?i��gԾO����r`>�J?S� ?4M�`م�.!&���>��>��-?f�e���_���Խ��>jN?��>���������Ž'�D>��?Q�?��*="�l�\���:��=��?Ƙ�?�;4?H}�%�;�[!о�=Ʉ�>�?���>pDW�����������>�N*??�>�ξz�u��
�`o	?&ma?�&��ŏ>aI�>.l>�.ݽ�gʾ
�X�멾����=��ӽO���u`�n��T�<�Ht> w>�j;�^^Ǿ_��>uB���N�i�H�<�����+R�<��?��q2>�i>�>>�(����Yω�(���L?���?ߊS?l8?"^�����R���~��=/��>�Ѭ>���=�����>I��>�e�xr�#�b�?�J�?���??\Z?��m���ʿ�Y����Ǿb־�-A�&��=�H>��F�R�=�Ν=�&��Y��'�@���|>�^J>�*�>f��>jD�>��5>�D���$�����������y�	W*���%������m�%銽�W'�����]�N4�����u ��5d������=��M~�ʨ���K?�2?�Hz>�|>�>�>6�)>����t�5��"i��5�oP�o�H�@o������]ž�;�\3&���>WS�i>h<?,�Լ��o>Zc?RC����>�ʇ��/8;W�>��=��>�զ����>�A�><�|><�="����s�L�>�QTs�����su;?��!����}0�H-ξb����H�>N(?1�4>k!�w���'{��F��>>=��_��E罃�s���>���>�տ=G�����c�DCl�1��1��=P�m>>e���:��5g���=K��>����� >��>��3?&��?�kL?��>~��>N�>�G!>�����	�� �'=�<�>:v)?��?;�1?c�?��4��5���?�=ѵ>�C����,�K�	�8\��?}����k<��k>h�K>��=2�V<'�=+%��$�=��=���>.|M?}��>�6�>���J�J���Z�"���c�;3*�5��>!S?��"?&2�>!9>��5��<��:�3��>�X�>�z��os����(>�/5>7�f?��#?NǼ=��J&.����|(<l�?f�,?0�3?gЕ=o̍=9: ��ҿ��s��w[��� ��I���΄=�����sT=+^�>�ͮ�����;���Jz=g�?�EQK=o@|�#=q>��>��>��7>e��=��D>?!r>�Li<�Ƀ=A>�o�:i ��H�3׵<�f8>_(>�~���@����Ʉ��$=&�?�d?�H<b�^p���߾ 耾���>��>}|�>��>��=���Y��+�������>��[?�u?J�E��]p=�ǟ=��=B1�>�%�>�"X>�1�a N�����*�p;���>�$?��>e1d�e��_��;��bw>ޢ���1���?.xS?�:�Bd��E��CU� ��P��>�J��IĽ�����R�Dc�T�C������k���&?f��?�s���j>ӣ��ε�����!N��˾����>:,?��?;T[>L|(��|����,a�㇠�O�K_&>Qг>�V?��<?�RX?ۺ;?�#D?='����>M-=S��>'+f>���>��>��d>���=P̍>�^�=������͛��R���^ý=�b=��>l�`>��=���v�=��,�e�>�uV���=K�/=0�̽փ�:�>��>=?�n'?E�����H�'>s��=9;���,>ȏ�=]�1��3þ���>��4>-1U>%�,?ދ>�b�=��Ͼ���Ѿ����/	6?̨I?�E�>�A.�
�>�J���I��y�> !>�/ѽCۊ��_㾀])�u6k���4=qi >7�=h>��p?�03?�V"?��Td7���q�{�,���A�%*����>�J�>�>�uƾw�'�`�l��[Y���?��qB��!��c�=F��=�$�=�u>�=4��=fπ=�)���0mμ�yy�N��>��>M
?�G>S>�=�L��E�EZ_?�|>�,�����-Ѽ��#���:�#? �>�C?@K�=�m������AZ��gJ?"t�?���?��R?���<����/�>�6�=�=�{>
�ĺ���>��n���>-�i<?/��:���އ�yM>.�O���&�x?���$:�\ɔ=ßɿЗj�h������&�z�Ծ�����E}��4�<pZ=70�������;�';�6��p@X��wA���w��s}�w�g?Z�X?�Q�<b�ͽ�?5�O����-�$=G7���'�</VC�Ne�����kȾ�y����+�f��C��,���>��Z��I����|���(�Ώ���?>�/?[?ƾ�x�����8!c=��$>��<��ؕ��e����
�(`W?/�9?5�4����0���>��?
f�>nX%>���J��?ۑ>|�3?��-?��㼭���"���ᑼ>J�?���??\K?�^��@C��4��Z��=O>?.-]?7�5>q3��Ւ�}L羄��>��{?o�g?���T1����{�m�3?��?R�޽vAD>]b�>��>�[g�O�T��!>~R�����w;���V=�p�=5�ȽY䧾�p�<@^�>�ӽ>	c�Z1�����>�/�_�N�c�H������(�<'�?�}�(U>�h>}>ް(�u��ω�=��L?���?z�S?�j8?�Q�����㧽&�=G�>ެ>-�=c��k۞>:��>W�;sr�:�֕?�H�?���?ZZ?'�m�j�Ϳ�������� ��&�����=��>0���j>ugH=ئ]��&F>��=���>���>�ڧ=�@�>owE>܋�=�V��� +�����ݨ� Rj�j#���&�ot������}4��)�]`���~žF<�=E�E��þ���S�뽞F��z��=�##?�$�>p��>z6�>f"}>�+�m�{ҽ��H�uf��!t����uL�����z���I�5gq��b0��3���>�<#؎=[%?���>t�?>sg��>oQ>�Z>3c�>�B =�p�=�uo=`0�>Pqk>�[ϼ�
2�4]���䅿8T��vX���>4r?g���K�F T��4�r���/>�?ۤ�>���7L��}XH���>�+=�X�A#���V��A�=&��>�V�=��5��Rb��zؽδ�=�j>��>m�>w������Ӝ@����=�'?���<z�S�>n�>QuS?q�Q?���>��>�"A?�b����H>��� �r�P���Zx>,<+?i???��@?�_?�I�=1�%�f��4��&�<��!��C�զ=��>�H�=C��m�^=��k����޽��=P��#���	>�U�>��*?a��>��	?	�����I�i�-� �n��������=~��>aXx>��0?z��>�~�=[���:�M����B%�i��>���>K1n�=�S��y�������v?&q?�`?���=x��r�	>�����=U@�>7Mk?9,?ۊ�>m�9�%���Vܿje��}��bx�[w>�^>'���B�����>���� ������=x=�B�>�>��>Ec>g��=�Ӿ>eB>fz.=q�=>��1>��#>����ߞ���A�.��O�U�}�����-�U' �6}&>2;��b׽+��<��&?�?��&��i���[</s�� :־Io�>�W?)��>??�>E���|��*��M̼oA?28n?ǣ?9�8�9ާ=�M�=��K�,��>���>0�>vJ�/�T�f6n��<>[��>?�S>ў%�݆j��j��
Ǿi��>�#�1*��A�?y[;?Fܭ��rA��=���;�w1�Y�Ž)B9>�D$������"�t�Q
L��:Q������>�L�>XL�?Y�;>���>&���W(���0�����r\ ��z�>��> ]3��H&=.�=�������]M��歾&\�h�>�(�>���>.�$?0W?�=?a�>�Sm��ޮ>�Y����>|��>�F�>��%?��?~M�>�?=>E�R>ٞý����b
����=!�ҽB>scy>�
X>7n�<A��=C��h�D���ؽ�������)�=$ƣ=a>M�>૵>��?a$?LqJ�]��=2QW��n׾�}�j��>��>u�!�U��zal���>�E�>
�-?�ɥ>��;>Me����Ծ���<�9?�!?ߦ?��=���XC߾&p����>�>��A�P���� �����*5��d�2>�4�>�3I<���=G4`?�LU?��#?�ꔽ �9�->y��
S�8�x^>���>&|��).t>͍��:�M��B��wʅ�g�X��ˇ<����ی>��=�K�>v�=Jo�2L
>\��<�1�y��҇�=8�̽���>���>|y-?��>C3R>_��J1���I?�՝���������cоX�6�y�>�^E>����2�?R����|�T)��E�=�w��>��?�,�?>�b?W�B����/Z>�*X>�s>��!<�k>���%��:����/>#��=p?v���� bE���X>��{>�Ͻ��Ⱦ�8��O��r���R���!���Ѿ`���E˾٭�N�ҽx����ܽ�cQ���~�����Խ��:�W����ѯ�ᥣ�9ߕ?L�?���=1EF���/��-�3��t��=����O�	�l3������
���п��c��	���0-���)�N=�C�>�[���t�c2e��D�kVS=N��>Y�*?ޅӾQǾK�	�d��=9�K>��Ȼw��]��0�����gB?.?�D�=�=���(Z>�'?��>"�>>����t��9f�>�;?w4?H]�<�������h嶽��?���?Yw>?�ZR��u<����*��/ ?��
?X�>�O��t�Ծl�н:�	?�@;?���>�p��Y�����x�>�\Z?��G���[>o�>Y��>��򽥻���hs�����h#3>b� �;��s�`��M/��ʢ=�J�>WWp>�$Z��P��/��=m��ؖ����^��ܾ� ��[=��p>�"�?޹=���>��4>:	ܾ�?r�6,��8F����P?�? [2?��%?����q�,��qC߼��(>�ф>x�=E�*�u�:>1��>�`�����E�jU�>���?m#�?]@@?3m[���Ŀ˵��̀��򾎰��f5>��>�^�<SDy=�	Խ�;�=��d=���=�g�>�%�=<RO>�Jj>'Q>g�>�����-��ӈ�V����f���Q�a�*DI��0(�U���R9羢�~�����L�A�b�H��������<vH�R��5	>�m?v�1?���>���>��>�,<���̾5I��I�B�I��k��ھ�2�$���B�������Z��p��<~�Q!�>y���=�M�>
 >�z>E;�>�+�=7�5>�ɽ���=�F>�5>�y�>�o5���=�|�>��9>&��=�P����i���=��ð�.~��,�=?pt�Ryt�)"1������p0���w>io�>t�>���e��@���֋�>z��2e�ӑL��%1=i>Bھ> k�=��u<�F�;V� ���<:	=���>�'#>�e�v�J��>;��� >H�>.ː���>�v�>V:7?km?��;?�8e����>Bp�>yL�>;]!��緽��,<�e�>:��>��>�7!?[dH?�l=^���.
{>�Um=�t��q��Vg�/g�='S��a�A�Ҽ?��<z�y=�[<�]:;J
�i���8\i=eŬ�i��>�K?0A�>�?�>��j���B��M��'=�/(>J��<�����b>�~*>��>��>�F�>�ꀾ>n'��H
�xB�>��>�(8��4P�����6�U��(>7sE?�f)?� }>I.��G0��>����>lTU?�B�>���=ZEڽ�X���ҿK�*�n�$��֝�,�,���:-]c��N����(��۽X�<��S>2�d>g�X>�Ma>k7>ؼ#>Vs�>��F>���=�=����qj���a�@zJ=�f���KN�E*?��r�<R �U�\�n�di�x�Լ����?%�T?f�?e��?������P�� W
�ڐ�>&��>�?��?�t<�� ���P��:�X������>�?E?�e?Sn=�s2,=گ�<�>��>��>��&>�7��K�`�p#H>�k�>�"
?��^>�b���^���Y���4e�>ʥ���&<>r?^�-?аھ��뾮*1��';�g������r��x��M�Y�]���o��vH�Ԙ�a�k���Ƚ�!?�ϩ?�T��Ri=�3��,���_��HBþ�a�>���>@�<
��>�L�$[�=��-s����A�j��%���R>���>��*?���>S�C?�.?q��>ػ��+?�V8����>? 7>`�>�ۚ>q�> ��>A>jy�=��h=���[����=��=<>|ռ>���>��=�=#R]=���=�5��?�<�ms��g����2=-���(�;a� >��?��2?��G;�ּ9�P�Ug�.�Z�vӯ>�	?v�t=�3Ծ�i��R�+��->�N?f��>U*�=��從�w�l���ݽ}P?��#?�>U�>+�>;���?�����l�>�K�<Mľ��i�m�����:J>ݓ[>��>�ǈ>4e?(*?��?�y���Q�(�x��n��ʓ����>�?��=M���ݪϾyE��K��M�Sv��9ǽ9U�=w�\>���=R>ݮ=`}�=>@I>��<����9G�R�>�X>���>��?�v>Ԡ;��;����Ͼ��I?EM���z�ᒢ�s2Ӿh�0�f�>�H>$�Ľxo?p����������<���>o�?iS�?�&`?F*?�Z��hY>��X>��>�A�;#�3�9޼���!�3>�o�=��n�=-����$�F^>��n>}ٽ�ľ\�޾�K���̿�i��溾����n���U���9���'�����8I3�ZW�b��+�=�>Ȩ̾�)��O�%)�}xݾ��\?#Z]?@�8�|=�0$��X��O���@ ���rV��Ml��S�+Z��.[��%f�hM��	���#��z徴�}�?�C3��5��ZA�[v=��W>��?i��gԾO����r`>�J?S� ?4M�`م�.!&���>��>��-?f�e���_���Խ��>jN?��>���������Ž'�D>��?Q�?��*="�l�\���:��=��?Ƙ�?�;4?H}�%�;�[!о�=Ʉ�>�?���>pDW�����������>�N*??�>�ξz�u��
�`o	?&ma?�&��ŏ>aI�>.l>�.ݽ�gʾ
�X�멾����=��ӽO���u`�n��T�<�Ht> w>�j;�^^Ǿ_��>uB���N�i�H�<�����+R�<��?��q2>�i>�>>�(����Yω�(���L?���?ߊS?l8?"^�����R���~��=/��>�Ѭ>���=�����>I��>�e�xr�#�b�?�J�?���??\Z?��m���ʿ�Y����Ǿb־�-A�&��=�H>��F�R�=�Ν=�&��Y��'�@���|>�^J>�*�>f��>jD�>��5>�D���$�����������y�	W*���%������m�%銽�W'�����]�N4�����u ��5d������=��M~�ʨ���K?�2?�Hz>�|>�>�>6�)>����t�5��"i��5�oP�o�H�@o������]ž�;�\3&���>WS�i>h<?,�Լ��o>Zc?RC����>�ʇ��/8;W�>��=��>�զ����>�A�><�|><�="����s�L�>�QTs�����su;?��!����}0�H-ξb����H�>N(?1�4>k!�w���'{��F��>>=��_��E罃�s���>���>�տ=G�����c�DCl�1��1��=P�m>>e���:��5g���=K��>����� >��>��3?&��?�kL?��>~��>N�>�G!>�����	�� �'=�<�>:v)?��?;�1?c�?��4��5���?�=ѵ>�C����,�K�	�8\��?}����k<��k>h�K>��=2�V<'�=+%��$�=��=���>.|M?}��>�6�>���J�J���Z�"���c�;3*�5��>!S?��"?&2�>!9>��5��<��:�3��>�X�>�z��os����(>�/5>7�f?��#?NǼ=��J&.����|(<l�?f�,?0�3?gЕ=o̍=9: ��ҿ��s��w[��� ��I���΄=�����sT=+^�>�ͮ�����;���Jz=g�?�EQK=o@|�#=q>��>��>��7>e��=��D>?!r>�Li<�Ƀ=A>�o�:i ��H�3׵<�f8>_(>�~���@����Ʉ��$=&�?�d?�H<b�^p���߾ 耾���>��>}|�>��>��=���Y��+�������>��[?�u?J�E��]p=�ǟ=��=B1�>�%�>�"X>�1�a N�����*�p;���>�$?��>e1d�e��_��;��bw>ޢ���1���?.xS?�:�Bd��E��CU� ��P��>�J��IĽ�����R�Dc�T�C������k���&?f��?�s���j>ӣ��ε�����!N��˾����>:,?��?;T[>L|(��|����,a�㇠�O�K_&>Qг>�V?��<?�RX?ۺ;?�#D?='����>M-=S��>'+f>���>��>��d>���=P̍>�^�=������͛��R���^ý=�b=��>l�`>��=���v�=��,�e�>�uV���=K�/=0�̽փ�:�>��>=?�n'?E�����H�'>s��=9;���,>ȏ�=]�1��3þ���>��4>-1U>%�,?ދ>�b�=��Ͼ���Ѿ����/	6?̨I?�E�>�A.�
�>�J���I��y�> !>�/ѽCۊ��_㾀])�u6k���4=qi >7�=h>��p?�03?�V"?��Td7���q�{�,���A�%*����>�J�>�>�uƾw�'�`�l��[Y���?��qB��!��c�=F��=�$�=�u>�=4��=fπ=�)���0mμ�yy�N��>��>M
?�G>S>�=�L��E�EZ_?�|>�,�����-Ѽ��#���:�#? �>�C?@K�=�m������AZ��gJ?"t�?���?��R?���<����/�>�6�=�=�{>
�ĺ���>��n���>-�i<?/��:���އ�yM>.�O���&�x?���$:�\ɔ=ßɿЗj�h������&�z�Ծ�����E}��4�<pZ=70�������;�';�6��p@X��wA���w��s}�w�g?Z�X?�Q�<b�ͽ�?5�O����-�$=G7���'�</VC�Ne�����kȾ�y����+�f��C��,���>��Z��I����|���(�Ώ���?>�/?[?ƾ�x�����8!c=��$>��<��ؕ��e����
�(`W?/�9?5�4����0���>��?
f�>nX%>���J��?ۑ>|�3?��-?��㼭���"���ᑼ>J�?���??\K?�^��@C��4��Z��=O>?.-]?7�5>q3��Ւ�}L羄��>��{?o�g?���T1����{�m�3?��?R�޽vAD>]b�>��>�[g�O�T��!>~R�����w;���V=�p�=5�ȽY䧾�p�<@^�>�ӽ>	c�Z1���6�>�r(��	���{��	��V�=�>a�t>�${���=�1-=��?F�,����q2N��r��ǇG?ҁ�?��A?h]?1�,�!V$��Ĥ���>+O??,>�>ai�>AL��N�>�\6?���j0Z��-h��i�>�?.8�?��?җ9���ῴߜ�f����.���X7>,cf:��;´�7�=>s���鶼�Il>G2�>t�>��C>�5>fmW>���=.p��v� �����%P���O�v�%�(�̻��?��s2
������ؾ����8��<���s���V����8����c�V��<~k�>���>�u�>���>�Yx>tڳ��v����J�%�辞2)�ξ ����?�x�^��慼ݵe�F����.����-�?P�׽���=��>��Ľ�m�=��>�~I=g�>Ӂ>%�=�M>�>Eh>ޝ�=�ڄ>d`o=B�>ҹ;>_�~�]�����Չ�
~޽�]?	;g�R��#�.Q��$��6��>v��>>�>e7�=���O��#9�>�1*�葽��#��2�HQ�>S��>��{=&�<y�3J��$?.���<�Z>Ē>�w�=╾x��?ؔ�)��>�h��	�z=/#&>�"?Vt?;�L?k��2��>�yl>��>ooļ�=c��<B_�>k_)?��8?˿?i�>VT=�D˽�;>�)����
���Gz���佺����ٞ��כ<7�;"��(7=��k=�O�=Ia��P9>������>��F?�S�>���>�K�_�E��@�QO<�HV=1�=�>r��>u�?��?B��>�m=��R����i������>ݜB>�VP��c�`�=��$>�s�=C�X?�>�>~�����=���߽lv�=�?��>Q�"?��>�t�:z�־?���9ӿ�@&���!�9�Z���M��ˢ�0�c��?u�u�=Q<����Z�k=�>�>�@�>c�Q>Ը=>�� >��->{��>��I>(tG=~��<jBB�Q<u�����;>�<���;�^y��ͼ�U���%��m��y�s�<�E��Z��1;A�>��8?kb�����2���J�{�Ӿ���>/�->'�>�-?~��E׾�9�s���_�>)?��~?4ɺ>�N��J�2=��
:�=�s�<ym=,��>�
1=~�$�н��G>M ?M%9?8��>����0����A����	���>�'1=�[�����?��P?����m��@���G����r<�N��Z�����F���<%���׾�{羓T9��u�=�%�>X:�?�Hl���=�����ɓ�ׇ������ބ=v�<��>-�>��P�C���̲��}�����F��=0U�>\VM�oP?�\?�1Y?���?΁?
Id>����:?����&�
?8K�>��U?�A?��?�)�>������"���=�C4��;���u��h��s�>ɇ >��=0�K���>�;�<�t�<̳�>�[���׽�׼��=��>){>���>Ѫ?�&�>��=xw�=�⽿-X��i���>j��A�_Ó��c��Z�>�J?��(?3w�>,SK��d�/�e����ԏ=��%?�D?o��>W��=|$%=Ԑ־쟭���ν鍍>��<�н���Ņ��i����>k��>3�,>T*D>��y?�j�>͆P?������$�A��Rջ�X� �VA��ޡ>���>a��>X���9�Y�	�m���d�{X�T �>�����=��<紲=E��>��=$�=QW�=XO���N��.Ƚ�L���L�>f��>CN�>��T>6���P���׼�t�Z?����/��Ⱦ�v"�չ>�f�>S:�>+��0?��=��P�%��R�*�:�9?ᐹ?�j�?�+??3�%�J\,����>0�\>�^�>�o���B�^�5�� ��p�=�=��-����>S`>�n1>� ���D�X]���ʿ>g5��2��񾫭��xE	�����T>ž�v��uf��|ݾ����b���M�4bB�f菾K����D��Y̠���?r�?@�>�ݗ��M�^D�jZ�K�F=���b¾�3���$�ʲ־HR��p߾��:���?�C�'�bf̾r�r=��7�lg[��ɉ�=_:��pi��),>�à>NC�����FF2��X>�=~�0��.�����b��cz*��Z?KA?�=���i���b��=_��>D�?��>�𜾦I����>3�6?��?�Yt��v������<%&�?9H�?�L??��<���A�C'�w����>�?���>[N���[ľ�C�~�
?a0;?z�>\������W����>��V?�J��]>|J�>D,�>����ܐ�8�0�ō�L��Z2/>�W|�<*���f��@,���=���>CMu>U�a�4ۼ���?O�r�{�c������8�>	�>Z�.?&����>� ?��+?C�'�s���>��!ƾ"pB?z��?�e?�(H?
�)�K�J��.����{>�A?zR�>�>�B��a���H?mu���}k��ﯾ���>���?��?��;?YJ"�ۜտ�U��qܩ��款��c>8I>��=ͩ~�%=3&ɼ'��[�~��3(>z�>\��>�bX>��s>jl�>�SK>�k���  �i��/j��]2W�w� �X�U��������+�@��A�����ö�7��m��)�������9��	`ڽ�����y�=�	?l�>9�>�$>$��>�)����l�|ľjo�ѳ����n��������ѽoE�΀��=�?��ȷ
?G����K(>�>�a��6:>DԜ>6mR=m�>�A>�I>-1Z>%C>�x7>�(�=y�q>d�=ef>��=q�x��Cv��7��`��'��6�8?5<X�������-���о�4�����>���>��)>�-����7r��m2�>��s��[������U�>7��>���=��	��_��x�[��~=�]>ɽ�=2�S�vݏ�X ὅu�=���>a�߾��\>,��=�J?��S?�YP?豽l�>)�>BN�=�|2��{Y=���=��>�.&?��6?�)?��>��=6;�b>x�=|�����S��=_������KἳG���=��Z=U?=�U�=[[���>�޳���?�O?3�_>�2?	�=�`BA��|4�ܑ�=dˊ>4�=�]�> B�>;(?-l/?네>��=c����i �{�����>�I!>�B_� 4k��<�=I�.>.�>m*Y?Q��>3hԽ�:�q񃽥Ƽ�:�?���>h,?&Y�>�:�=�ҿ���+Cÿ1�����0���Y��ܾf4�<�L����K�'m�=*��>l^�>i�z=�"7>�8�=`��=mR�>s�C>�a=���=����^��N��=]+>\[�;Qn��e�н��[=��=�����˛��lU�!�����8P�� $?apC?8V	�UW�g���?����#�?>�?��O?a�?H!H>���T��c��>{r��>�>+�}?H$?��&��A>j'<>����=�Q.>�=T:��"6��!��w�<���>��P?�[�>��3��������<�1��g�>�^=���R$�?KDT?�d��#\m���6SE�9����<	��#������ ���.��oվf
���G��hu=$��>�å?�C����
>�@þK��������A���!�<��=~.�>�>��A��֭�W, �!/��C.3���3=�K�>��G��A�>~�Q?�r?��?4V�>�#�>T�y�(?�]���>�U�>�|O?o�? #
?��4>N�>��@���>��5���>��>_�nH���>���=�,l>�jɽ�GO>�4=���<uVF=A�$���<PD��ᠲ�ǝ�=nX=�>9�?Zc?��Խc1>�{��1�8�),}=~�>��ѽ_���>K�9�:�[ګ>|14?t�2?s��>3���K�����Z��A6��TA?lW?>��>���=�u��R�����������=x�I;�$U=v�!���7���=ø�>w�>��>tc>�Y�?��(?�?<닾��&��T��}žt�>s��<�k�>�d�=��(>���Z��������]<� �>A5��q͠<p7c=�Y�>Ғ>�b>GeK=���=�'<��5�<��<W��N��>��>x�?s�m>ʇ��s���+��;uJ?b�����7�ξ�� �ie�>�>F�>��ed�>YA@���������I�x��>�Q�?��?�8e?P�|���4��l?�?>!՟>94X�����4��l0U;���>kp�>��־���\���Eo>Wg�=�
��X%�Z���d>o�6&���t�#[=�;q������{��3�����j����D	�T�=qS��Ľj��<��v�����Fd���7�	��?��?�,�>7�ʽ^9S����&7��T1�����T��y��v;u���J���.�Ծ+���M���M��dA�ϒE>���QGP�]v�ń2�y�I����=�>�Ҿ�l���3��"�=H�=ZCS�����������4'D��0?q�T?���x������3��=�?�(?�ž>�BH�s�>�`>��?�E?N��Tx��=�h�=C��?��?)�??�7O�ȠA�F����?+�?���>Ê��̾N&�s ?c�9?��>#��N���-���>wy[?��N�gb>���>2�>��ｭ���kh&��������f-9>�����}�g��Q>�Q§=��>�x>�4]��Ү�<� ?�d�3r��Ӑ�,�\�>�>Gn0?ˉ����=u��>�:	?����y�wb��9���QP?&1�?g	d?rF?>:���'�|u=�*�>{�?0��>�����K>��=�=!�3?�C���{}��
����(?@�?��?
�T?xpO���ҿ.�����Ҿ`ғ�v�>���=3x,=��}�=)���1:ǽS:
<��>�!�>ܙ�>�I4>�1>U,>��=P���Ћ)� 3��Z���}\�V� �����'���S0���r�3	�x��Ͽ��'HX��*���+�48���������6�лG<�!?�q>t~B>T��=���>�����N�^��!�����D^!�^b��7p������=fi��f��'8Ǿ�� ?W5	;��;>`@>%��<�78=O3�>v;�= f���<R��=K��>�d>��>��=F��>��bߖ>y:>�~��wp�0�'�V���)&��OdZ?� ����X��M)����B������>"�?�{)>1�.�����؈�Z��>�V<�-?��X	�W�=�ܘ>���>�S>�
=�_��g�V��~��w10='N�>�Z>8�2=Y@�֛Ľr�M=���>��վ��=��v>�^)?�/v?T6?�!�=E��>�V>�~�>��=��J>l�K>Q�>�?��8?��0?
�>{�=$�Z��#!=e�=�9�zda��e���_�wc/�oU7<�
H��LB=yr=>M<��d=>=��㼳��;���<!?�M?��>���>FDM���E��[��T<Q�=�.�=�O�>^�t>�?�/?�{�>b��=xJf�)���]��,�>�=>�3M��r��Θ=�B,>t�8>�]?�?�`��U�����9�ז�
2�>�X?xE/?d��>�;�<����� �`?Ͽ�MB�ժ�j��=#��={����-��K���ki=���0�*>��8=���=~�(>A5*����=���=KL��h�>�m>b��=��<V�K=^=�޼8��=��G�[��1�4��<`J��Y��t�o��<��(�@a>�7uǼ\m?�??�Pz�P�=q���WY���P���?���>�+?�.?�*���#��O"�f���C拾~
�>KbX?�?�>� ���=���i�)���>�̣>���>u�;��H<U��9�=��'?��?�)
?h7�@}��|˩���o���B?�]=P=����?<jT?���縕���
��N�]����R;kH��߄�F�ƾ��#��+4�s����G�-��vX=�>��?�>��r��=�]��]�����������<��p=�K�>�	>=�V�������������w�!C=�_�>5�ڼE��>q
?�s7?\�?��?,�=uT7�aMr?��ɾP�?��0?�eL?<�?�J:?|�>2L�R����;���"�S��n����(�b�a>�o�=f�>1e;��=���=�G}��ۧ=��8��<����]���D�]=��U>$3`=��?�-#?j=s>��@>�b��z�=��	����>@����>�b1�#v����>Y�B?7`F?ޭ�>��ȽII����z��_p ��5? ;?y\�>l,,>7
�=�*�i���CM&�^�+>@=j�>�"&��YȽ��=c�x>sפ>h��>#�>�>�?C	?\�=?T�r�W*2��=7���F>cǤ>��>�;>؟>f"׽�ZP��o���㊿�<�� �>�/-	<�q	>������=Y��=��m��?7=}f� ���j�=f���G>�d�>�&?��>�P=�� �PS�sJ?NOb���վ������%�ºA���?l���_�t^�=� ���t���|��J���Q�`>�`�?���?���?�b��fMT��?�	>�	?u��	
޾�W��눽��m��n�=�TŽ������ƽ��D>B���r��:��і�9�v��5<��/r=-m�`h��6t�������'�V�پ.+��F�ԂG�XQ����E��P���!d��í���ľ�Gʾ\�?8z�?J�>���G�M���$��~
���k>����F�(='~����@� ������ƾdi'�{ I��u9��羃�j>7'B��z"�cד��:A�N7%���?=��,?XZ�I�E�j�c�c���'�">	mU�+�����Λ���ѽ��N?Ss?�A�679�8T�r��?�.?��> s�=��=�x�>��<?z�?Z{�b���Yb����!>9��?�?!??�����B�C���(����>�o?Ѫ�>=�c�a��f��i�?T.;?zQ�>�i�)&����'��>`^x?X[���`>��>"�>˽�)c��DC��殾��i�>�p����������*�C�>�0�>��>>1匾/��m@�>����D�.�x����&頺}C?U�+?�����>�AJ=��4>���|���d��S�O�S?�V�?k�s?��y?]a�c!?� ��w0�$�i?X�3>�� ?̨r��?k|�>��	�[�����Ņ]?�=�?�@�$?��D��:׿�=����˾���=�U"=��=�=���$1=�=R�_����=��>��>�U>��2>p�>�R>��>yւ��; ��&�� f��Hsb���4���<�����͍+��G�)'��.t��-����ɽV�ƽ�6ѽ��Y�(�9�bꚽ/
��|��=��?�
�>O��>}/�=ЫG>�ʾ�����b�ؾ��%�8��R���)���<(*�9/��4W�Qr���d�u(˾OR�>X�<��&>�V�>+8^��k=��>���<�L>�>">F
�=���=[�n=O>"�Z>��b>��>�ax>��={ā��,~��@6�ai�����5�=? 2o�0X��i/�!ҾN����>��?fA>��(��j���e����>��U�	�q��ֽ0�P����>��>v��=AD&<\⼾�q��ݽ���=U�w>�o�=xLK�[��d���å=J'�>�\�m��=@��>V�?��e?;�4?7N�=���>!і>�>c��(>i�=��>��)?�^/?�/?ͻ>I�	=5��h�=�����O������=����5��n�<��:��?��6c�=�PJ�&=Sr.=2 ���任��<و�>ңK?��>{M�>~Kp�ݺ0��_d�j,��
�7<���� d�>Y��>,�?.?��>4H�=$�X���(�����.�>#�9>�b��u���&9�=�g�>FP?�e�>�蓽�[W���=���=��>��?��??ٜ�>~�=�M��;��|������8��
���M�M��a�Ǿ,j޾?�Ǿq���tu>��=?�i>�P�=��>Y��<f)�;��@���>�o>T�=��<q�����p<u�=զB>ԟ��j��d1V�E��;��B<�����P���7�<B����Z�x�w��??�2E?o晾�W�����y�H��h�>`E?�?�>!�'?Q��>���)O��耿�������>o�?�?�
�g�,>�>�|�H1>/��>���<�$I<9MT�5�����>�(?�+ ?� �>�����Ϗ�ℿW&��f�>5I=���?Y?�c��ţ��� �@hV��/���;�h��@���7��:�$�[{.�D�ؾ#:�eW_���=0�>-�?���¸�=ճ�zᓿ�]��߈��?%=�Z^=( �>�=*>�\�ხ�(��>T���V��y4=���>��;c�>�J?�q?��?l��>�Pk>�X;)�?͌����9?g�
?. 9?&6?�6�>�p>�C�=kg�<��&<��F��롐�ʂ�*�>B��=E?>_
U<�
>���lܽt,9<=z�=��<�@<jiE<R>��3>��?��>|��<!Z3>nG���c��Xy߽ٝo>��C<幬<�f��� ��Y�|>m
?�?���>�Y�=^ĳ�����XV�<:�=�>?)�D?�A'?���<�>�b׾Ւ�M>㼇�>��x;, ��|���ɾ3�p���s>k9�>�:j�gIb>|*�?Ǥ?l@$?X���f���B��� ���={����m�>o�=�l>	J����F�Rt���܈�����q�>Dװ�ͦ�<��=(z�=Ub.>�	�����9�+}|���ͽ����V��s>�;�>E�?W��>3��+��&�)@`?����.�|��N���W�>��>�u�>H/=�FO?�+���;��]��O���LA?� �?"U�?���>'{�z��.�?��=:��>*�D��4ľf"󽮋���@�>W%�=��o�ۅJ�v��=>3�>�<I�O�s�þ�3�Zۼ�͸��x��+����1&����\	��3����C���x������b9�QgA��e:���u��x������K��k(�?�%�?�h>{P�����ۅ)��T¾����4���?>��� L��<�ž����<��Cl�	b �-�C��?�1>D]"���[�};�������s�R>	f�>e��ZȞ��m.��
�=u8>)�����,b��H@���Y>���0?/iE?��C�;����J>#�?�%4?N��>��1�����r>��.?�1?Ce��^��ad���]�<6�?���?�7?�&��Z�9�ڢ���$^�>�*�>�^�>�Ɣ�������L�d�
?;�:?\��>4w�1���pX�j�>C=]?d�T�yn>���>�6�>mP-��8i��]���ы�(�Ҽ׶)>L�۽=�M�;���c�4��=�>��Y>�.y�/�i��Ů>҈��>�0��U���=|����>��?y��g�?�)�=���U���R��iop���Q��B?�ǹ?O�U?��~?�*�9[]� V=��=��\?���>{��>�]Q>��?}F�>�QݾV��ܣ��@TY?���?P@nD:?�U����-[��Z�ƾD�⾅>�o�<U��=i����T>
��<A���Ƚ;��>�1�>��=&G>,SZ>씢=��u=���r�#�ߔ��,R���0_�����-��Vs��q��e�wD&��E������Rw���L�+�����<����j|���%>��?�_�>���>�:>o!�=�����
��D~��ޤ����S�\����¾T[��k��0�`<����Ľ5�����>+׹<��	>���>+�j�"� >}��>�h|=È(>b�^>^g(>�4>��>�N2>�W->�l>���=3��>�O=)Q���x|��i>�$�M��Jn=.�E?X�*����8�w��/��;�>��?=r>zc�\���jr�H��>8� �%xJ�ѧ��g��|vf>��>Є�=7�"�>!F�5�ʦ��|>�!u>�;>\kA��∾�i����=��>�nӾ���=�!>�(?v?P�2?�/�=2�>�[>ϟ�>Y!�=�wO>�Q>���>"�?��9?[J1?f�>���=�][���=�C=�);���S����ؼ�@*�R�m<��9��FQ=�;�=f��;ϔ\=pS>=ˤļ ��;��=�e�>ï)?���>�5 ?"6I�[��r^��Tv��Ng�����?|&�>^�?��?��k>8�=B8��t����>n>��(
T�A,��O���O�>���>=�Z?#B?p=�y(��p�>!�>�h�>�,�>��#?$"�>� >ԧ�	�4ӿ,�#�<F"��9�ӵ���:�PA�)+Y�H�ͺ�5.�7C���p�<��Z>a̅>�p>ɻC>�;>�0>��>�%K>�ӑ=��=%�:u��YS���?=��O�<��X�3��.�ż=ғ�����L��,>�͈����<Z�>|�f?�4� �s���վlL'�sr��
�">#��>n�6?���>l-�<�[޾|�
H_�'��C�>�ĉ?��?�"�2F>��/�0��!%<��2=�d>�k��M3�=�����;�>�3?�7?d��>�2Ͼ�a���e��z@/��O	?x��<�d��|�???G�羳c`����W�K���''=!}�n���:1߾_L��������iȾd��=��=A��>���?��{�$HK> ?��ڒ������=1E� �H��=T��>q�>=����o:־ϕU�<��#�%w�>�%i>^5�>��=��?N (?W
�?zBA?(,���<�P/>y�徆D
?H�K?[�H?��?�Q�=��>!�>��>y��?�Q½�#�<���EA>b�]=h��=��W<6�<����h<�;=c������rڊ�%9�0�����h�F�=i�
?��s>N�	��>
׮���;���>�Ї>D��>B�����1���l�.<���>՗K?��?�+���߾�_ �M�ؾ�á=�l8?~�(?��?�<�=3窽<+�1���B"�M�]>�����Q(�<ܟ����&lt>K~�>��>-��=⨕?SQ?�@	? -��G�:�:<�*���m����R���	?^�]>Lz+=�Q�?�i��畿�@���pM�EU�>�b�����f�>��i>��>��7>VW�z�=>w,\�l#l�t�=�p���E>M��>4�?6�>B��=WN��`�G�;��?��;�����$������ͯ�>?�ֶ>$�b>��P?w�ǒ��Pʿ�݉���a?�4�?���?-��>�ຼh%	�D��>eC
>7J>ƍ&�sܾ��^kk�S
>�d����=%Ͼ�ܖ=���>٣�>��h�^x�	׾_�k<�ҿ�!)�K�r=�'�P找kl�L����_'�W���}�ݾ(A2�qA���'��[ݽ�Fp�S ��v5侥aҾE5�?���?m#�>��A�h^Q�$�3�I�Ⱦ�t�=��t�g����y��؅��kȾaXؾЂ0�T;���(Ŧ�~'&>g/K��u�����p)��4T�#J>�5?Q1������(45=�!>�|ֽq� �� ��i����?�I7U?wH?�����9�Ľ��=��?�?MO>HRq����=+_>8?�=-?E>4�Z���3���H҂<+��?�t�?��>?eC���A��������?�C?`�>�܆�CȾY콳B?o'9?U�>Z�Z���G���>�]?jUN�V(a>K�>�Ø>Ț��̒���F�(f���a��Ո(>bA�s��. g��G>���=LW�>o7n>��d�o����7�>rs*�`�.�C�{�̌!������s�=o1?�C*�٪!?X=�C�(��g���w��-�a�l?�?�1?@�?��{��kT��Չ�%��>���>$?�
r>��D=n?�i"?���?7����[�>=�?���?�`?�/l�9Gӿ��!������5��=�$�=��>>
�޽�ɭ=��K=�Θ�[=�R�>t��>�o>9;x>}�T>ۛ<>��.>n�����#��ʤ�2ْ��[B�� ����.wg��{	��y�����ȴ��񽾤���t���OГ���G�j��nT>��浾�"M>)��>K�?2��>�k���nQ����@R�P���׾��	�N$�����~[�T��������N�{ق��1����>m�0����=�л>�/�A��<��4>�7^=醕=�A�<��=�:���m=>PU=�����>DZ�>��>�>6#��������*�a�ֽ�l�=P&9?UcX��m��^'�I�wߔ���>>(?��&>�(�I㙿]&x�Pѳ>Q�B�i6��r��I��KWd>�ݻ>�B�=�XA= Ї�t���l�ƽD �<tck>�{v>����y�h"��X<�B�>��۾\��=#�z>̷*?�Pu?¦6?�@�=qi�>hj>���>���=��F>�cD>���>҆?�
<?��1?���>և�=��[�'�=��e=(YA���}������������G<�D�6�=�/O=i�#<�0�=0�W=���i}���=S��>�w5?(�>�\�>��U�#&>��cM�������=�+!����>���>>^?Q��>�5�>q�=,���q���ȇž���>��U>L�X��J���t��w��>2=�>�	P?Α$?1 =�g�S�:=,K->�o�>��>;M?в�>���=�1H: ��mӿ�$�-�!��>Q�qو;��<�k�M��7E�-�[�����<�\>/�>��p>�E>��>�<3>�R�>�HG>�ф=�={<�;)�;��E���M=�
��CG<�P�����)&Ƽ^��������I�G�>�`:�7ټ���>S$�>_�A�Û�=��P��d!��-i>G@�>���>�0>��<~� ��Z9�]dJ�-ı���>#:?f��>��a���X>�½�\=�;�>��>=,��ƽj�����}��3>�/�>j�?���>�'��8h�L�b�ھb�>"�{�\˽�Y�?�[Y?%������Ĺ"���<���#������z&��Y���Mg*�jPC�������,`P�fb>b?N��?�ዾ&o�;j���˓��s��}��Gi�=vFR>�&�>P)>��l������ojž��V^�=��>s�>Wda?.�>��k?���>=C�>�!���,?s�ܾ��?h(t?�!?�Oa?�*S?d��=4�4�]h�{���&j�-p��0̯�޲ܼHHc>9��=��
���N=
[\>`Nj=j���+^<H�Q^��0x��>��r>��>�)>���>�!C?V�����˾�Ԍ=���<�~�>#o˽���>�%w��� � �;�)\>��"?ީW?.66>vt/��:<�R`I�����=��U?�[6?��B>������M��������|�/=+�>�{������T�n�@���=R9�>�>1h=Jg?��>X�?̥���mh�
&��fa���㎼^iX�LE�>v��>
���';L�4�,�c�0d>�H����3>� ����4>�0>�M��
��;J�z>U-�>nm�����n>�������>�N>j�>��V=Hd�'L��>��d�p?a^�<�8�l>�<�澾��[=��>�R�>���=�RR?�\F�/�_�R��3)P�-��>EF�?��?(u?�8��k�־�?��>4{>����)�ľޯZ�����5�>L53�eP��oy��`�����>;jI>��
��ھ��޾5h��#ҿ�K?�]�=�]����21��M���ӽ�� ��t����-�rq��.m���Ӎ���T����k���)�y�Ӡ���_�?�d�?�n�>F�=""�^�þE���0�>/&�N����)�3�о4{_�(���j
����d)� ��.D���>�Iҽ��A�d�1�:�w=Y�2>Ӿ\?a���tO�*����<|��>}'<����:��:���A&��m?��N?,��SZ�-��E��=�OV?F�-?4iF>��þzm=��>�?��Z?�ѻ>���|ah�S�P�?�K�?�RN?���= �[��z=���-�-gb?|�L?1�?G�ʾ?aS�dJ>|LS>y�y?�?����u�.�9�gk"�Ծ5?
tI���>��'>��4=w;�=f!I��	�=��2->�,D���0={׎������->5Y�>r��>�>F��� ��S?�z�<.��0cU�-ھ��>��>F??��!���>I��>;�?>���skW�n��DJa=��p?�/�?�Gx?�>?����ܾ�W�=>�>�X=gN">6ڽ� �8>=�>�+>6�Ӿ�6s���F�u��>Os�?��?L�N?Bq��ӿኙ�Fڸ�i���G�\�|���-=��½4`=��u��V�(�=�>%?�>]�>��f>�Z?>�Q=�������>�-���8̕�*{f�=�1�t9��0y���"�>CW��M�)�;��ʾ���QGC��q��CJ�R�R����/������=H=?�,�>��1>�� v=�*���Ş�Gj��rXI����1���.��s��2���hw �ؿ	�X�ѽm���� ?!g�=��s�Z��>6c��e@z=��=R.�<�3I>�i>5Ӯ>OkA>��=�PY>�1>y9�>�L>[�w>�#}=� ������:���V�H��;3�A?�IZ�hᘾ��4��߾ī���|>w4?o�S>_�&��6���%z���>_�6��,X��Ƚ�'�-��>��>b��=_xr�����bv��K��=�>�~�=�>����������=��>K�ѾI�="ŀ>[$'?�s?��4?-2�=+�>��`>��>�:�=��@>RR>>P�>;}?\�;?�2?0�>ŧ�=�aY�?��<��4==���[�E�����Ƽ�� ���<���*�\=��N=<�0<KC=�`*=ա���6N<���<��>$�;?�>�v?�d]�u�'�z
r���"=��Ͻ��=��	?F߿=��>X}�>S�f>l��=Q�+<�G������>ׂq>sBn��ꇿ�� �K�_>�B>��b?�(?��'>ʓ���^>������=���>��&?���>f>��>����{�����VN��rվR��Joi��ұ�Z�E���G�D��~�	>K)>ˈ=l��=���r�r/v�:�߽�}�>f��>�`}=	�o>�կ:�t�=EY�=�d$����u~=��xA>\�1��T(��g����y��v�F��R�<vP$?�_?�p���O>�<e���)y�� ?(��>��f?��^?�5�=y>�p�辇�_�m�սZ�9?;;�?O��>�4�F��<��=�D>�7�>�&>�M=����5x��?;���>Fe4>��?a"�>lF�={Wo�g腿S�"��q�>R��=�½�*�?,�_?и�e��"��l9�w ��3K�Q%��+e������3�2���<����bp���=���>"�?PXv����=�G������7z�]����C+=�>�=���>~�%>8ڀ����LK�yuʾ)\�k�fW�>�D��b?�e6?b��>z��?��5?�s?mWN�!�s?�:W��Y�>ɹ,?I�F?�r?hU�?����F�M����%=h�&�j�p��
;���U�f=�'2>eȺ=R>��>��.�G#�l���K�=��=C�,=%��=0�=T��=��=�?�?���=�>����?,�����=I�M=���=�������ZG\��>�Ƚ>)��>��?�6&>�~x�J&�:�ھs��>G(�>�F?�Z?��<�x�=�ᾍ��>.=�h>m����;��� �־0m�͵�>�(�>Kh�=��t>T)�?�b?�iO?ժ2>�^3�se��N����=vu���W>��|>�Ͻ۸���۾U����c���c��I�t夾;��=��N>��=�~�=wS=ě=lX��_�����ς��ϕc�bn�>�>N� ?�[>>��䖾L�~+f?���3�S.Ľ�%����;U�>�b�>�<�pX�>i%Ǿ�"����s�P�K�&�>��?��?��D?��E=�M���=�>@,�>@��=�&���/���r�:Wݽɮ�>���;��ϾR~c�q$p�F�<c�T>0����������Ծ�߲��eM�&�������cҾA﮾��Ծ��0����V��d�i�)�:���F;�� �5TQ�����b�3蟾���?��R?X�`>Eᴽ5=�����w��>uw����n���پ� m�3|�s�վ��ھ�E��������QN�>��w��݀��ϊ�~V��!x>���>̴9?������q�侔tɼ`��>����}v��~|��Z��*�}?��?�#�j�T��о�=�b�?��g?� �>�!���������>$�C?8?
��>	��+�P��sw>֠�?˻?i�??��N�tHA��4�����?�b?�Y�>�犾+c;2�
?��9?���>��m�������>]�[?B#O��0b>�4�>�o�>)uｶ����.�[W���[���<6>��E�l>���i�MR>��G�=�\�>�lu>7�^�쮾#!�>ؕ,�C-��p`����zwR=���>�� ?�&�SXr>F;�>���=����D�U�!v���4Z�"�P?nq�?�O?C5?����|��}�z>�#���S�����<]z>���=Z�>8�>�����t���X�8��> 8�?'��?k�L?��;Gӿ�� ��������=%�=��>>��޽�ɭ=w�K=T˘��Z=�l�>z��>o>F;x>}�T>ۛ<>��.>q�����#��ʤ�4ْ��[B�� ���wg��{	��y�����ȴ���C�������VГ���G�U��&U>��p������B=?� �>��>B~M��>�������;���ܾ�K@� ��c�| ��1�����0�������+�ݳվ���>A�<F��Y��>G�=��⾽gV�>n=�8�=�i$>�a1>�ko>|�7>C�M>��t>��7>� �=��{> Ǉ=~�����f:�>oQ�]i�;��C??]��S����3�v߾i����Ȅ>��?y�S>k'�������x����>�zG�*c��̽����E�>���>��=��Ȼ��?~w����Д�=�m�>��
>��l�����-	�bG�=��?G�����r�
pS>��?\Ny?EG?	�\>5��>X�R>���>��l>AM�<z�>сc>�u?yD7?C�J?���>�.x=�K�qp�=�v�:�g���ݾ�2_ȼkH�VxἙ�>�`&��-R=(P�=�e�=,��=5E�yZQ�������=�c�>�R?���>Ĭ#?5���#9�h�N�P
��s>MH=$��=��T>���>}�>a��>��>�!>���u�ܾoh�>ڟ>�me�c�a�NY\<}��=��7>8[?��J?xad<P1,��r>&���H�> ��>�?���>��>q���'����ѿ�."�{Q%�J�d��r'�����KZ�ʛ��BEE���<�r�Ͻ~�=q�f>ū�>'�f>~�0>�V�=͗7>w��>��|>#�=��=�B<�8��-\��?�w=~����/�mo���(
���J�ڸŽm@�CN#�����jC �6;;��:?I�>����[�Y�J�t�0ȾN=���-?�x�>]�4?7�?���<~�,��M�O��Q<��v�?T0_?�v�>{݆��d�=[
�;J�=p�>+Ϟ>=OZ>]׆��xþ?e�89�>9��>B�?ȉ}>[��=$�>��y^�	��g��>��#=P5p���?n�h?����S��w���uP�[�8=d���ѥľ₞��!$�+�2燾�3��r�[�����>��>}�?{8־���>Wl�� �������q��k�A>v1�=��B>`0>����I����þ�B�
m�=b�>����>�N侁�:?�? �=sO�?3-F?v
?V*�0�?،�����>�]E? �d?�n?��l?Z���R������p�E��hK1�3�==B�A?�=%�>�$=�C�r�=l���Ā%��:�=�EU=sd�=��=_r�<쐅<'�j=��=���>j�"?9�������Rj�;��ڽ%��@�=�G>��˽�A�f<5�{>�) ?�E5?��>RG�<h���O��u�����	>�?�)?+��>�l��r�3=����K�� �p=˄j>_����+��ә��rb��B���~>c��>�i>�>���?��?.�H?��M>ё+�8�u���P!>������>ch�>���<�}�ؑ��߀�=�w��n���=�g���O�=%&>ك=��X>��S=u�={�<�C�=�8�M�G�̖Z��j�>�)�>�b�>D�x>Ly�=Ï�}�)��
D?��/����\�<u �f�ľ�cD��9�>�=r�?j���-j�w_���a[����� �?�x�?Or?�`����%{=[i>%~��
<�Ԁ��D6�j���̢H<$vڽh����A�Y�0e�DmF>�̽�<̾>�׽�]B��`��U�T�B�B�{O�0�ž�����;���E��;)�{Hؾ���5�y���۽��*�<3��n���K�t��H�q�oЕ?_�?��v>�:�c	M�������>��J�>�uƾ\�=u:��,�Ͼ����A��o���;}�P	�����v5n>�!��g�A���ElW��2�>8?o�&?��6�i�K�� ����;m�t>�O>E ����������M���?ϴ�?��S�͘T��=���Px>��K?��<?�=3jD��K=�g�>,�O?��.?��S>W���ʏ�ذ�=��?�^�?��@?��<���<�+:�_潾h�>3�?���>)����(��i��;v?u6/?���>ʮ�򑆿�V�@��>��d?����u��>��>Q��>n���!���Xt��ĝ�8hz��M�=����ߤ�ʘo���/��f�=1ʊ>�@�=Wp��:n���
?�p-�����i~�?r��c~�>}��>E?@N��6�<*�?^zt>�Z��X����]4��k?_x�?�q?��6?ۄ�*x��4�$>&-t>�Y��]�=�~�.՞<2��>>�>�2�[�[��k���>m��?!�?2-A?b�n�Ѽؿן��2�¾<릾y��=�E�<y>?����[;����T�E=-�=.f">�.1>�l>`[[>z|�=eZ=@�v<K���$%(��J��aϑ�'�V�+5<�h�����U�������S����V���F�����$=�����1����AF��y�=?G<?Ҏ�>۴�>�{p��բ=��q���ݾ����X-��P�E�澾J�v�����&��;w<�g^ﾴ ӽ�s����>� u>��M=j�>�-�T��O,>B��=�(�~p�;�%%>&�j>;>w��>�ݠ>!�B>��D>�z>)n�=���8����:�r�Q�I��;*�C?�J]������3��s߾�}����><�?>�S>��'�u���G�x�R��>p}G��_b���ʽ`!�RL�>�k�>���=�̻,P�r�v��O��ŷ=���>��
>�Mn�����-
���=7p�>�־L�=ǲz>0�'?� u?�x5?c;�=�>u)d>��>e�=	J>r�K>���> �?�9?N�1?R��>��=-tZ��7=4�F=��A���[�����U?��,%��*�<��B���>=1�i=>�<�c=�J=Q���F�;j�<R��>�,?��>�?t�;���E���`��o >�w�>��> e�>`Q�>%J�>:b�>
��>Qw+>aP�<C�<�m/z�hp�>��>�v��k�o=���>�ߠ>�E?R?��=�ٽ�ǁ>�ל<N�>���>�m ?���>A�|>qE�Z���7ſC�$��>��Ⱦb,���2�S1�����<V���4,_�0Os�N�7>�:>(I�>�6>��=��w����>�J=���=��=��0�f";W���7�>_v1<-	�=�3G>�C�&�H�B�=�����" �$NӼ��T����=|?/?>���=�'�	��s� �
�\?�q�>d$s?��>:�>�<a�}Q0���6�����)?I�v?mx�>i{f�5y�=�g��1��3 ?I�=ñ�=*mٽ,���_�E����=i1�>1i?��>P�=��V���Y����`?��M<���p��?�^?��I�}���%���?�Tz��N=`�k�𧧾uQ��pv��X8�G�Ծ�޾*��{��=kt?��?Y���}�<v�ƾ�V����\�-����K�=TR�= �>I�C>�R��z���#���׾���+�6>|?�>�h���Q�>�PR?Kћ>��9?�?z�>�I��H	?"���+�>]1:?�l?U.\?s�^?4`���ƾٜ�AYF�����rh��H=�`��pb�=���=�M�=;�=y!���~��ˆ�=���<��;���u�5>��u>R�1>ڟ=�'�=̷
?�!?�ı�P ������8.�z�<xC�=��d>�<�<}��0���;A>x��>�N ?��> �=��ԾsUﾦ�����
>�N?��.?���>!<�;�`2=���0�t�Gf�<�P2>�V4����v��]����8�N�>P@r>���=�BQ>��?�7?�c=?8�>���.@���1����>����O|�>(��>	]s>�*B�n�
�s��j���'S������~�߲�;K�>a1K>�g�=K��>T�>r�]��%_��8��S����p�>9��>�i�>2�Z>k��=9���/-���H?�����[�=H:�PR�R��>@��=̛��D/?����H��Fʄ����N��<lZ�?�ͻ?j�w?�Y��2[����>=\�>���=S<��Ǿ���VH3=;##>%!>J��^���j�ԾoRO=��4>b�:���ݾIb��J���ش��`\�\ᗽ�\��V|�������b����+���'����9W��=/���օ�8�q���q����W����e_�?zZ�?;��>��q�E���(��hA��2��1־N�.l��yR�a׽�X����l��o�"�\��)v���݆>q�4���s�����lX��<�>6��>�2?5W�_�L����<\n��+ >��=�S��;���낿P�=>q?m�?)-�ںX��(þ��">ބ~?a�h?o�>0ֿ���/�0r�>��o?
J?x��>q�}�J�|��B�>��?���?,F?nψ=�V��v��5��>7�>�R�>TE�>۽�s��(�=��?QQ'?�%?�����闿K�'�T��>��?�s��]�v>jQ�>�AR>iVþR5�����=\���U�>��9�8_�=����C=i����,i=APF>�`^�0GӾI��
?�p-�����i~�?r��c~�>}��>E?@N��6�<*�?^zt>�Z��X����]4��k?_x�?�q?��6?ۄ�*x��4�$>&-t>�Y��]�=�~�.՞<2��>>�>�2�[�[��k���>m��?!�?2-A?b�n�Ѽؿן��2�¾<릾y��=�E�<y>?����[;����T�E=-�=.f">�.1>�l>`[[>z|�=eZ=@�v<K���$%(��J��aϑ�'�V�+5<�h�����U�������S����V���F�����$=�����1����AF��y�=?G<?Ҏ�>۴�>�{p��բ=��q���ݾ����X-��P�E�澾J�v�����&��;w<�g^ﾴ ӽ�s����>� u>��M=j�>�-�T��O,>B��=�(�~p�;�%%>&�j>;>w��>�ݠ>!�B>��D>�z>)n�=���8����:�r�Q�I��;*�C?�J]������3��s߾�}����><�?>�S>��'�u���G�x�R��>p}G��_b���ʽ`!�RL�>�k�>���=�̻,P�r�v��O��ŷ=���>��
>�Mn�����-
���=7p�>�־L�=ǲz>0�'?� u?�x5?c;�=�>u)d>��>e�=	J>r�K>���> �?�9?N�1?R��>��=-tZ��7=4�F=��A���[�����U?��,%��*�<��B���>=1�i=>�<�c=�J=Q���F�;j�<R��>�,?��>�?t�;���E���`��o >�w�>��> e�>`Q�>%J�>:b�>
��>Qw+>aP�<C�<�m/z�hp�>��>�v��k�o=���>�ߠ>�E?R?��=�ٽ�ǁ>�ל<N�>���>�m ?���>A�|>qE�Z���7ſC�$��>��Ⱦb,���2�S1�����<V���4,_�0Os�N�7>�:>(I�>�6>��=��w����>�J=���=��=��0�f";W���7�>_v1<-	�=�3G>�C�&�H�B�=�����" �$NӼ��T����=|?/?>���=�'�	��s� �
�\?�q�>d$s?��>:�>�<a�}Q0���6�����)?I�v?mx�>i{f�5y�=�g��1��3 ?I�=ñ�=*mٽ,���_�E����=i1�>1i?��>P�=��V���Y����`?��M<���p��?�^?��I�}���%���?�Tz��N=`�k�𧧾uQ��pv��X8�G�Ծ�޾*��{��=kt?��?Y���}�<v�ƾ�V����\�-����K�=TR�= �>I�C>�R��z���#���׾���+�6>|?�>�h���Q�>�PR?Kћ>��9?�?z�>�I��H	?"���+�>]1:?�l?U.\?s�^?4`���ƾٜ�AYF�����rh��H=�`��pb�=���=�M�=;�=y!���~��ˆ�=���<��;���u�5>��u>R�1>ڟ=�'�=̷
?�!?�ı�P ������8.�z�<xC�=��d>�<�<}��0���;A>x��>�N ?��> �=��ԾsUﾦ�����
>�N?��.?���>!<�;�`2=���0�t�Gf�<�P2>�V4����v��]����8�N�>P@r>���=�BQ>��?�7?�c=?8�>���.@���1����>����O|�>(��>	]s>�*B�n�
�s��j���'S������~�߲�;K�>a1K>�g�=K��>T�>r�]��%_��8��S����p�>9��>�i�>2�Z>k��=9���/-���H?�����[�=H:�PR�R��>@��=̛��D/?����H��Fʄ����N��<lZ�?�ͻ?j�w?�Y��2[����>=\�>���=S<��Ǿ���VH3=;##>%!>J��^���j�ԾoRO=��4>b�:���ݾIb��J���ش��`\�\ᗽ�\��V|�������b����+���'����9W��=/���օ�8�q���q����W����e_�?zZ�?;��>��q�E���(��hA��2��1־N�.l��yR�a׽�X����l��o�"�\��)v���݆>q�4���s�����lX��<�>6��>�2?5W�_�L����<\n��+ >��=�S��;���낿P�=>q?m�?)-�ںX��(þ��">ބ~?a�h?o�>0ֿ���/�0r�>��o?
J?x��>q�}�J�|��B�>��?���?,F?nψ=�V��v��5��>7�>�R�>TE�>۽�s��(�=��?QQ'?�%?�����闿K�'�T��>��?�s��]�v>jQ�>�AR>iVþR5�����=\���U�>��9�8_�=����C=i����,i=APF>�`^�0GӾI��r�> Z�~��oq�����ͽPiľ�=0)���_����9�W�5W澸$��P{�q���f`?�I�?U�?��l?����ea��\�=�*O�x:/>���>.ov>c�H�l��=.��=��m��r��֟�t-?�K�?�n�?8�>?��R�+�ҿ�p���6ʾ�:ʾ7P=5[n=��!>$�C����= �%>gB�=��<(0P>��>��Y>�S;>H�<>{ i>Ǵ�>�p����.��ǌ����$��	�������;ھ� 	�J������Ǎ�{(�ֽ�"ǽm�E���=�X��Rĵ����=m��>ɠ8��?��$>+�`�]'������(����D�_�߾!���Ͼ�p��p����]����k�=�9�x�>� �>�?e��=��=��>�"ɽ��=��=�������7>��>��>��>��>���>�^>X���7yv��<�^pw�	��=��[?0����y>��:�[����=�?�9�>�'�|H���.��xg>�2��[)��;-Že��=瑴>�8>�� >�3Z=���93�*�j���>��&>�k>�_=�J����/���=~g?���ǻ��C�>��#?�Gn?�F%?<�@=9>��?>�!J>@�B>CH�<F�i>�E�>*�4?�-?��?��?.�=z<�?�Q=��=ӈ��i���<�}н�Y��ԋ�=��!����ɍ�<Z�=A�=��}=\2���4����o=]� ?��@?Qb�>�]�>{���J���Q�,�x)�р>C�>�3?��>d?�'E?~ݟ>8�ӽ�z޽s����vǕ>Z�=��+�LXH���<;a�>R�=�
K?��"?s��+�%=8��<�O>a��>݋�>n>.?���>LD'>P��<�D
�	z����*���Y�=&؃=zV�=���V�=>�g*>����8z�=15>d��>�5>�`�=7G>2`�=�{�=[��>iM>��_>;E7=�h=��#=,���>l��l��]�
�pm�9�_�<-��<mXC�ν�0@���<gfx��'����?<�?�_S�vv�=tf��T����<���%K�D�н��C>ܧ>i���iW���w��
��45?0�?�D?��{��=�(<`��z�>�i2>�G>�x���Y�<ť�Hc���D>U?)W�>V�Q�~�v�N�Z��`�����>�C�=~�����?�Z?���=:%�����;� c�����;g��;�=�����,�@l0���پ-��k4���=\�>4��?*�w�Ѡ>ؖ��E����E�3X	��Uh��[�8>�>y��>����N��j�3�E[�����3�H>c�L>)�z��N?x]E?��%?�s*?�L?���>]+Z>�h1?���>�?yi)?�9?.��>���>&�>�ꃾ�@��'b=H/����ꍽ_�H�v�2z����^�p�W��ܻD=���Iֽ�)��ŕ<��=��=
��=R�=�	>I�>��?��<>�Q�[ą��=�$�>j��>)E�+=�h = \T>�>?f��>���>ȶ=g+�������i��M�->��?�6:?	�?��?}b�>�x�u����S6����{6>�NŽ��$�޴�~�)�>��><W>8i�>��f?m�'?s�V?a�޾�oA���q����x=��(=Jg�>I>�	>�n{���~�z��[c�����̾3��&�=#�	>�P0�w�=�?�S�0�[>H>��9=��>�݂>*^=���>�R�>t�?R#>�(����/�n?.�S������׾�� ��҉�s��=��>�����m�>��P�a�܄��	
��I�<?I�?�;�?���>��>o���'�>�6�=k#>�����4�P�s>4�Z>��<>`�<'����!����W���+>��L=�JK�g�u�J�x=A ���k,��:@=��/�����þWy�,�W������,����G�3)�=I�/��s��|�I'�������� �q܉?��N?�C>��p��3�ښ �5iA��%>�:�˾�L�ィ�����=v�W����Ծ �@��
��v;����>���L��*v��9��3<�=F-?{��X?Ǿ��!�x��;/��=�q��Ͼ.[t����f �~�T?��;??���4�����[�'[�=s�?�k�>��z=�����*g�:�C>�>?�L:?WT�����*�����<@�?C�?b??D����!��{����`�Z`?�_'?y�>Q�о{ �UM�[��>��?��>6A+�{���j���'?ɨf?�f2��&>"�>O��>�W[�1z¾������xa>���>*��=�����_��x*��nZ>�>�x=,�Ͼ�����>���6�ό����B������6��𧿾�0��I������E��>e��J�^��E}?"G�?��,?��g?����h!�� ���<#s�>Bɱ=C{>𬑾0��=0�>�ླK\��� �Z`:?��?��?�W�?�S�I�ٿ'.��SS߾ܾ́�k=\�=8_�>a}�`��=�[>D?D�*����C>�O>@l�>�4�>�@>j{%>xL>�N��~E!�� ���Β��G7������7�H�^����%=�hþ�i��Q�ؾ��	�u��<�ţ=��]��P!�̴[�����B�6>��?a�>��>��8>��)>��s��⾔�X�\�������Ӿ�^��u�ž�ُ�;
q�\�x��S��@����W𾖽�>�|��>��>���<�>�b�>e��<ݕ�=�</>�� >�H\>�$(>�DK>9m$>��E>J��=���>���=
����}�̻�S���b��;fDi?�־�E��c�*�Y���)��
>�N)?_0�>M��D��>3���&>f�</G�����YY���Β>j��=p�>�J>MG�+���f����>݃>��V>�_
=�Y2�����9�7>�
?'!����@�>��*?�dQ?q+$?ў�=.Ȣ>��>��a>�(>��K>q�>���>6)?	�?�,?�^,?|n�=�*����=J�=|���HW���Q<s�������<y�w�d�����e>z�>�p�=Dj0�S����#��g��=�A?]W?U�>l�?T����y���l����=o>���\�G?�k?�ܯ>o�+?��H>^J�"9�=��'��:����>pY>0���O���>�w>�X�>u=?Th??mm�=G��;���=��=�C�>m{j>J�I?£�>�?�(7=W�	�\�Ŀ���^P'��k��&��3m��
{�F5���V>J�u=R#�<�W�=��>@R�>�T�>�c1>36�=��=��>L��>5˘>�=I>p��=�*��`:�D�<�D<O�<K�=T�=(h��G`<3鼽����Gc����ѽ7�Ľ�'?��!?w�<
đ=6}��sKľ�ʏ�\2�>�R�>�>�?CZ]=���ë5�QgT����@��>�u?=��>c _�|/�=��=_)�=���>��>}�:>/e=��Ľ��ڽp�輍>�>6�?��f>��YL�Bu����4�>�sL>n��=� [?�@_?��>�Oy&=� ��� I��^��>��sb��z]�����]�<�w�K���,��������U��=��>1 �?+���>T���6���S�$�����=��8?(��=�iJ����+<�	A��z�`�0u>#�#��s�>��P?�ɶ>��"?�?O?��S?���=;�??.��>�*�>b3?��I?d�>��'>cú�|e���>�#�4�Ͻ�cI��)�3L��L�=l�=c�>�~ �?��<@�<����f�=�<>�ʏc�J�=2�=/�=J�ʼ���=7�?-_ ?�ý��U����'���{<��>3�>LQ��)Q���T����=L?2�?�%�>�>z�.�־Ϋ�[/;��2?7?���>k��>@�F>Ep��?uV��fc=Y�>54��`�h�龺�����нxB>׫�>�YB>j�>�f?/�"?��X?��������k��C�i�5�b�s>�}�=���v�#��S@�mÕ�l�q��*U�Gp&=��c�Ǻ+=1c=�]�<Z߄>7��=ָE>��@>;�Q=�9|=����:��;Bv�>D��>�%?hC�>7�̫¾p�"��|`?jQ��X�9r���w��ሬ���˽&�{>���c.�<�Z־	���l�����1?���?H�?�1?�`)>��>�r=kE>��"?�X���|=W�j>���mAQ�*�5=\���iG̼!'R��� ��>];�$����Ҿ5��=���|�(�(�=����_=lM۾����ؾ�p ���a=B���h�[=+�">);:���\��e�_�l�� �KU ��ǆ?�Q?2l�=��M��tD����2���30���νz���j��Ҁ�� >�{�;U	� �Wp��)kӾ:T��t�>5ғ�`S����r�,��:� �B1#>4$?�齾#���%�P��=�J>׃<lվ9�{�󱗿i�����[?�<7?�a뾬��4Ե�u�>*�?;��>W�>r����$ǽđ>��)?�Z4?��C=T8����������ѷ?��?~`a?���[p����ݳ�L��>ܧ?u��>p7���3~�ٙ6����>�2#?`�"?�j�@�@�V(���>%,�?��2�y�>�|�>�!>�@��lӦ�\T�;)������=�=�¦� d��d����==Ȝ>9��>a����m�R_"?��R�=���[[{�гž� M>x]f>"^??�����u����>o֐>Ǽ��$-��K����ͽ��z?�w�?qze?��G?+���Z��re>�W�=�)M>�e)>��a>l�U�s
?Z��>M8X�־MH�G?���?
��?�?ZL^����$�������>ľ
��=_4B=7>-��g3>k���<���<\D�=6`�>+W�>�Ŧ>�h>`z>nx!>���T� ��̔��Έ��'(�[��z0�냖�x)ؾ:i8�%���@q�@������n��]�=� ͽn�����1����T>j��>�>=�>Ȳ�=��=/<����!���˾��+�� �
&�V��o�k�a,���v�.{ʾ��ȼ�YU�>=��t	>>}�>CP缍�>�,�>�" <l��=��>>n�=Apz=We>��E>N�=c�S> j&>T�C>C��=��v�9��L[-�h�z����b�3?��T��H��
�0����x���Z>���>^�:>�(�>������(�>�Lw����dA���<"ٗ>���>�S=6��<����^���u����=�p>@��=� ��L��a��`>���>g�ľ7�	>;9>Q�(?�_z?Bx.?�u�=w��>\�>{̕>T>|�u>�W>���>�?ݗ/?ߛ,?R��>��=�b���U<�=<�x��)�of��<˽h[O��[=���x�=��=B�����=��<�چ���<�s�=�n�>��M?5&�>��.?fh���H_�L<�3�ҽ#��=@�i=7�0?�,?*3
?ٖ4?�8�>�����4����r	�:z>9>�%�3I��G>�L�>���>]C5?fS?��">�e2�?R;$~n>P�S>�x�>J�=?�w�>v��>�y.�/���	׿G��%�K���i�ݼ���;��1�ڒ���:<��	�;ފ�:��=Z�k>,֝>Z�n>��A>ۑI>*�T>ߍ�>�ψ>��=�=6=��< g~�$	��V��)��1+��A齄V������,�	|�<���ue���,���,��.�?1�$?�½9*�<�������t�a��_�=�r���iw�?��=�Ѽ��ā�.`��F��t�>��?�B&?B/���>�) =�̦���x>���=(Pn=��=��3>>94�,{|>(9�>�6�>;Oi>��X�y�O�fo�c�	���>זO>��l�2�p?��S?B�,�P�=��@��Q�a�:/�M���`s�~"��Ձ'�m1��;F�N��w���B��r�X>���>�K�?�!��͑>$���*@����d��F�����=��L�k�>�^>~����1����)�ʿ$����6���T>�K����>�5)?��r>�e?�eA?7��>|�=��f?��2?!3�>B?ȜK?vG0?�H5?�P>uԫ�D���آ>��Ľ�N�-2���$p�����S��=���=3=�y>]A��z��͞�UË�������<V�}��p~=�3�=]k>�{?�W1?��!�t9�=b�U���:�I�?=��>�$>1E&=2bp����=3��>Ic?�s+? D�>��<�ܾ�a�� N��i�=C�$?*�
?=?��J>�OY>w󰾥�Y�8��=/+>�1�i����$��E;g�)>!��>��>��>o/?��"?-�{?%�.��~x���о(���Xu޽��&?]|�=����H��d	�I���~Q���o�c�ھ����|�=_�j=H2�>�V0>~ZG���T�@�>׼�`�
>��\>�k�=>�?�52?�?cjm>!�#=�S��;��H?�j�9sv���پ�2ؾ7� �1�>q!?�ž��7>�;�W����g��K��ģ>���?�;�?��f?f���,�T���W>T�?W��>�����x�;�&�=�j����x���;��@z��^��g�(��Xo>hX'>�S��J���8ߌ�g���l�ǿ��&��=R�aD�MU���h�i#����x��\��	��p���k��w�L<f�-�]�M���¾����vل?�eb?�_>өl;�Wξ�� �ٜ����`��څ��PS��X�������m��~/ξV辒)�A;�O�7��s�Ge;>�?s�v�v�ga���������KC�~�>�����ξy�>�����;ǈ�i�'��J�����k��b���B!B?C�b?1� �+;e�� ��
N�=�G!?!?���>��ң��r�>|�%?��>�s���`��#v�����>^��?�v�?'�??מI�(�@�z���b�?K?qw�>�����KӾ6��R	?��6?Ka�>8y�ss���f��j�>(\?d#M�Sd>���>0=�>
��RG��]�/��Ɛ�}�5���7>�"q��0���d�|�A�%��=(�>j�n>�Z��Ω��r�> Z�~��oq�����ͽPiľ�=0)���_����9�W�5W澸$��P{�q���f`?�I�?U�?��l?����ea��\�=�*O�x:/>���>.ov>c�H�l��=.��=��m��r��֟�t-?�K�?�n�?8�>?��R�+�ҿ�p���6ʾ�:ʾ7P=5[n=��!>$�C����= �%>gB�=��<(0P>��>��Y>�S;>H�<>{ i>Ǵ�>�p����.��ǌ����$��	�������;ھ� 	�J������Ǎ�{(�ֽ�"ǽm�E���=�X��Rĵ����=m��>ɠ8��?��$>+�`�]'������(����D�_�߾!���Ͼ�p��p����]����k�=�9�x�>� �>�?e��=��=��>�"ɽ��=��=�������7>��>��>��>��>���>�^>X���7yv��<�^pw�	��=��[?0����y>��:�[����=�?�9�>�'�|H���.��xg>�2��[)��;-Že��=瑴>�8>�� >�3Z=���93�*�j���>��&>�k>�_=�J����/���=~g?���ǻ��C�>��#?�Gn?�F%?<�@=9>��?>�!J>@�B>CH�<F�i>�E�>*�4?�-?��?��?.�=z<�?�Q=��=ӈ��i���<�}н�Y��ԋ�=��!����ɍ�<Z�=A�=��}=\2���4����o=]� ?��@?Qb�>�]�>{���J���Q�,�x)�р>C�>�3?��>d?�'E?~ݟ>8�ӽ�z޽s����vǕ>Z�=��+�LXH���<;a�>R�=�
K?��"?s��+�%=8��<�O>a��>݋�>n>.?���>LD'>P��<�D
�	z����*���Y�=&؃=zV�=���V�=>�g*>����8z�=15>d��>�5>�`�=7G>2`�=�{�=[��>iM>��_>;E7=�h=��#=,���>l��l��]�
�pm�9�_�<-��<mXC�ν�0@���<gfx��'����?<�?�_S�vv�=tf��T����<���%K�D�н��C>ܧ>i���iW���w��
��45?0�?�D?��{��=�(<`��z�>�i2>�G>�x���Y�<ť�Hc���D>U?)W�>V�Q�~�v�N�Z��`�����>�C�=~�����?�Z?���=:%�����;� c�����;g��;�=�����,�@l0���پ-��k4���=\�>4��?*�w�Ѡ>ؖ��E����E�3X	��Uh��[�8>�>y��>����N��j�3�E[�����3�H>c�L>)�z��N?x]E?��%?�s*?�L?���>]+Z>�h1?���>�?yi)?�9?.��>���>&�>�ꃾ�@��'b=H/����ꍽ_�H�v�2z����^�p�W��ܻD=���Iֽ�)��ŕ<��=��=
��=R�=�	>I�>��?��<>�Q�[ą��=�$�>j��>)E�+=�h = \T>�>?f��>���>ȶ=g+�������i��M�->��?�6:?	�?��?}b�>�x�u����S6����{6>�NŽ��$�޴�~�)�>��><W>8i�>��f?m�'?s�V?a�޾�oA���q����x=��(=Jg�>I>�	>�n{���~�z��[c�����̾3��&�=#�	>�P0�w�=�?�S�0�[>H>��9=��>�݂>*^=���>�R�>t�?R#>�(����/�n?.�S������׾�� ��҉�s��=��>�����m�>��P�a�܄��	
��I�<?I�?�;�?���>��>o���'�>�6�=k#>�����4�P�s>4�Z>��<>`�<'����!����W���+>��L=�JK�g�u�J�x=A ���k,��:@=��/�����þWy�,�W������,����G�3)�=I�/��s��|�I'�������� �q܉?��N?�C>��p��3�ښ �5iA��%>�:�˾�L�ィ�����=v�W����Ծ �@��
��v;����>���L��*v��9��3<�=F-?{��X?Ǿ��!�x��;/��=�q��Ͼ.[t����f �~�T?��;??���4�����[�'[�=s�?�k�>��z=�����*g�:�C>�>?�L:?WT�����*�����<@�?C�?b??D����!��{����`�Z`?�_'?y�>Q�о{ �UM�[��>��?��>6A+�{���j���'?ɨf?�f2��&>"�>O��>�W[�1z¾������xa>���>*��=�����_��x*��nZ>�>�x=,�Ͼ�����>���6�ό����B������6��𧿾�0��I������E��>e��J�^��E}?"G�?��,?��g?����h!�� ���<#s�>Bɱ=C{>𬑾0��=0�>�ླK\��� �Z`:?��?��?�W�?�S�I�ٿ'.��SS߾ܾ́�k=\�=8_�>a}�`��=�[>D?D�*����C>�O>@l�>�4�>�@>j{%>xL>�N��~E!�� ���Β��G7������7�H�^����%=�hþ�i��Q�ؾ��	�u��<�ţ=��]��P!�̴[�����B�6>��?a�>��>��8>��)>��s��⾔�X�\�������Ӿ�^��u�ž�ُ�;
q�\�x��S��@����W𾖽�>�|��>��>���<�>�b�>e��<ݕ�=�</>�� >�H\>�$(>�DK>9m$>��E>J��=���>���=
����}�̻�S���b��;fDi?�־�E��c�*�Y���)��
>�N)?_0�>M��D��>3���&>f�</G�����YY���Β>j��=p�>�J>MG�+���f����>݃>��V>�_
=�Y2�����9�7>�
?'!����@�>��*?�dQ?q+$?ў�=.Ȣ>��>��a>�(>��K>q�>���>6)?	�?�,?�^,?|n�=�*����=J�=|���HW���Q<s�������<y�w�d�����e>z�>�p�=Dj0�S����#��g��=�A?]W?U�>l�?T����y���l����=o>���\�G?�k?�ܯ>o�+?��H>^J�"9�=��'��:����>pY>0���O���>�w>�X�>u=?Th??mm�=G��;���=��=�C�>m{j>J�I?£�>�?�(7=W�	�\�Ŀ���^P'��k��&��3m��
{�F5���V>J�u=R#�<�W�=��>@R�>�T�>�c1>36�=��=��>L��>5˘>�=I>p��=�*��`:�D�<�D<O�<K�=T�=(h��G`<3鼽����Gc����ѽ7�Ľ�'?��!?w�<
đ=6}��sKľ�ʏ�\2�>�R�>�>�?CZ]=���ë5�QgT����@��>�u?=��>c _�|/�=��=_)�=���>��>}�:>/e=��Ľ��ڽp�輍>�>6�?��f>��YL�Bu����4�>�sL>n��=� [?�@_?��>�Oy&=� ��� I��^��>��sb��z]�����]�<�w�K���,��������U��=��>1 �?+���>T���6���S�$�����=��8?(��=�iJ����+<�	A��z�`�0u>#�#��s�>��P?�ɶ>��"?�?O?��S?���=;�??.��>�*�>b3?��I?d�>��'>cú�|e���>�#�4�Ͻ�cI��)�3L��L�=l�=c�>�~ �?��<@�<����f�=�<>�ʏc�J�=2�=/�=J�ʼ���=7�?-_ ?�ý��U����'���{<��>3�>LQ��)Q���T����=L?2�?�%�>�>z�.�־Ϋ�[/;��2?7?���>k��>@�F>Ep��?uV��fc=Y�>54��`�h�龺�����нxB>׫�>�YB>j�>�f?/�"?��X?��������k��C�i�5�b�s>�}�=���v�#��S@�mÕ�l�q��*U�Gp&=��c�Ǻ+=1c=�]�<Z߄>7��=ָE>��@>;�Q=�9|=����:��;Bv�>D��>�%?hC�>7�̫¾p�"��|`?jQ��X�9r���w��ሬ���˽&�{>���c.�<�Z־	���l�����1?���?H�?�1?�`)>��>�r=kE>��"?�X���|=W�j>���mAQ�*�5=\���iG̼!'R��� ��>];�$����Ҿ5��=���|�(�(�=����_=lM۾����ؾ�p ���a=B���h�[=+�">);:���\��e�_�l�� �KU ��ǆ?�Q?2l�=��M��tD����2���30���νz���j��Ҁ�� >�{�;U	� �Wp��)kӾ:T��t�>5ғ�`S����r�,��:� �B1#>4$?�齾#���%�P��=�J>׃<lվ9�{�󱗿i�����[?�<7?�a뾬��4Ե�u�>*�?;��>W�>r����$ǽđ>��)?�Z4?��C=T8����������ѷ?��?~`a?���[p����ݳ�L��>ܧ?u��>p7���3~�ٙ6����>�2#?`�"?�j�@�@�V(���>%,�?��2�y�>�|�>�!>�@��lӦ�\T�;)������=�=�¦� d��d����==Ȝ>9��>a����m��`�>����Uh��|(��>�>x��>�:?��B���>q��>�-3��x��Af�Xf���j=8\?W��?��\?h%K?w��0'�1g�idA>h�>�Y?�E=�`��#�>�v�>_q"��q�đ8�@8�>���?�U�?c?���	ٿ?)������]���M7>�|.<J�=��Ң>]ٷ=�0h<�8t=X.>멈>�X�=�*>:�>!�#>7�N>���� ��D���e��L�@�:.�+%��gG�E��C�q�<-�H����3�U�=�d&�I� �ŜN�g������G���>���>�RU>d��>�ƥ>�d�=/T��5P���
��(��H�پ��1�ܖ4���ȾQ���4b�=�<�g~�V�Q�L+�+�c?�iu��Fټ�z?��D�U�>� �>��>ӭ޼a��>�X�=@��>cGN>u'>F��>L�=*�`>���>[d�>	�k�4���g�J�����/���=G?�F�=>��-a����rԌ��Y?p�?>=Y�)������ߝ�7�>�pƽ]�g�����>씓>�?E{(>�I���Q>5޾W�Q�ء�����>L�>��=W,��W⽚<n� &�>���}�5>ڧE>t� ?��?�l+?�a�=�ϟ>�5><i>EW�=>�=�/>"�c>\?A�;?�-?�]�>���=��g���=iR�=Ϳg��X#�O���\	ؽT��:\�B%�oo���u=���<X�";���=V����)�L�<	?�2]?�Ց>�o�>��\�Z���m�_��y�>�b��(?�/?XX?ï?�O�>Jt9��Ҟ����'��b��>���>M�D�6Š�)�g�	��>�fl���>?v�d?b������CR=58L>��?�:?�>��>�J��E�H�	���ѿ��A�"�!��遾����b����<"�b>_���S!>c͉>�_�>d{>�\�=�ꋼٳ=��E��f��>�E>(. =�����l��W��=B|���?L�d<M[A���'<�ռ���2�����=�2q�� ��8���ܽ_N�>!@A?ب�x���G��_��\��� ��fn>r��=�2>�hj�e2� ���\25�{�y�0?�
i?��>8?X�1�=�#��|���>�Ɏ>����1��t��Dh;�-t>#�>,�G?dc�>�+�E_������*��H�>{bI=Ļ��5��?�b�?@���dp��w�����9�.������w �xAᾋl�3#���?��嘾gq�������K�="o�>�?;��2>'{�c)���k��f����=����><���r���p��iꮾjk���=#M>��>`7@>��=/5?��?�?�?��?R��>�]?���=6�?�bN?�D? .?/S?�n�<eP������ǽ�&��?��?����U��|1>��2>�(>����Z텽�;�;���=�<��x�t�����,@A�1�=i�=~d:>l>��#?BSK?8tѽ��@�f�:��L�UV<��u�>0��>��z>��Z�'=g��>��6?`sG?�>H�����+���@����n�����?K�C?8��>��"���=��w���z7��{E�E0�>���=�4T�H���Nћ��+�;V4">�L�>�ߠ>og>��w?�?}�c?ݚ-:�LC��X=�����-=A�m�.�>K��<q0E=`謾B=A���z��ua���$��<6>,5ƽ�L5��q�<��?	�*>!`��ҡ�>���=/�����*��g>n�<��>Æ�>H��>&�>�A۽Y��_��2&H?�W�mxI�����3�ҫ<��?L>�F���3:?9�b�K~��e붿sx�#(�>�C�?30�?eߒ?$$�>=t���.�>�g�>7��=�!X�5�Ӿ����S;=x��>���=sC����t���˼�.(�7.�>) ��h�оŗž�m��ꁿ��O��!r�O���6������辸K����H�N��^Ož��6�m�O� �½}?���y�ߏ���ݾ4žð�?�2�?N0�>�g�=��B��99�z�ԾD���*ྡw�������Vݾ��ƾ�	�������LF���1���;�A\>��T�����X���K���G�^�p=�P?�IվS����9����X�y�=Z�k�%�ځ�_Μ��$�ԾY?�"p?8��QW��ő�x�=%�;?	� ?���>P ���sM>玲>?Sd?�T�=	���g�ǂ'>
��?�g�?��??NO�ٝA��+��%�X+?H�?a�>_a��E�̾ "��6?m�9?��>����h��]7� x�>�@[?�^N��b>s��>�A�>.�h���DN$�����䇼<:>�+�����ph�uB>��q�=�>�cx>�\�
ˮ�z�=�2���w�7{�<�۾�^��	'>S�?�c���h">���>��=�e)��s��������%=��>?:j�?eRU?���?r2�i�Y��$��	�X>��,?��4?��J��e�����>y?f���о��wt��l�
?��?���?�K?n9��꿿���7~��m���O�=�3�<�q�=�d�ǡq=�9=nP=�j�%�>Zt>]�=y�>�J�=	�>�>s!��,�����v����H���(��C��xl�P���5������H������ڲ��Ǿr�!�_���mw���,=�b�Ha>\@b>#��>���>QY0>M��� �M�F��K�?tž�}?��4�����`Ul>Y8�>7�:��3�I��]x�Ξ?$߽zY>�M�>GZX���Q>�c�>L��=�%�=q
K>=!>��M=�?���=�J>��[=�=E��>LS�>��|�����$:��vH=LΒ��Z4?6�z�z����pA�Z��&����8�>��>��;=��<�y��nz����>F�w��E��~�<��!>m�,>���>��)>"�=�շ<�6оvY���Z;q�>/4�>
�=<I���c��t��@�>�C̾��=�v>%?yYt?�d-?�-p=Z!�>m+B>=6�>j��=�D;>[	M>�G�>��?vZ??t�1?XN�>Xj�=�_��=��.=�4���X�I���/=ż���7��<J)�	Od=3�R=�1K��32=<]$=����^�<[e�<I�?"�=?\�>��>�0���(>��c��q���>�=x��>lf�>�?=��>"�W>b�;,4��8ݾ��+��E�>���>��l�G��N���y'�>KRC>�zD?F�'?��;�G���Λ=�*�=:.�>���>
a?�z�>�48=�j����lӿ�$���!��悽�I��w�;U�<���M���7m�-�����Qb�<�\>��>��p>vE>��>:73>[Q�>�JG>EЄ=��=	G�;�;/ F��{M=���G<��P�Q��zTƼǡ�������I��>��K�aټ}��>�5?7�>�Wc;�a���̾*��X��=I�>Xhe>s�&>�H�<G���c�B�(�O�ۃ'�	�?��]?f��>i����мe�P��=8�m>=�*>�_w>!�=�WG��:>��>�??R<�>nOҽ(����Ξ���.��`�>浫�K�F���v?��`?���XM���v��m�v���sL=Α|�����}�A�4���M�S�۾o8۾������r>aW?��?�����;��Dǆ��߃��ި��f�>+:
>Y|�>�L�>w�8>�I�<"�پ�o�)�ɽo~9>�&�>�D�>��>�HA?�8?0:b?�#��TV�>���>�
?/]�><q�>��S?,*?��B?��?�1��w��GF:�H��G����g�ZK�=.FU=��=��=y��<����uF���=]=n�-fR<�͔<V=z>�A�<�C=��>$?قF?rk��y�A�4�s�6�ZM_=�#�>��>;�F=��达� >�n�>#�F?�]-?�H>�@��7�6yT��xپ�+"���?�vI?��>!!)���="؎�U{���Q��7�>�>p�ǾW���Zܕ��9��Z�>@8�>��<>��p>!�m?�34?	�"?u��X-���p�	���|G�x�H��x�>`1�>�F�=��Ǿ.*A�Ls��Tc�U�5�N�=��9���<:�x=;>1ll>h��=&[>�T�=���ѽ���<��0���>���>��>�uY>�z��/�޾>����1?�]��rt���I��q=>Ԍ?�Ӵ=d�z�-?}QS>Aҋ����c�^�O}?�H�?���?1�^?.3�=��t�8f ?0G�>�Ob>�01��ྺ2�a�<���=Q���!ݾ����:��9<�=�?肾5IȾ�;�!�Y9ĿH�b��K,�P�پª���,�ƶ�����F��cV8��(��S�����辇������"�R5���5���ᘾ��r?��5?>�&>˗�TsF�`�Ծр��Ѧ��[ �a��Zվ�r��>���3��۝�bZ¾G�����쮰�a�>��I�����{���-�S5��y"!>R/?����%�������U�=�
3>�׍<���2����������8]?e�9?���of �Z[���	>o�?�	�>�a+>v���s�	����>:�3?�
+?��%��o��3^���J߼��?p��?[[?�e<=*QD�[<������?廞>X*�>h㔽v��+l���2?�T?U��>��k�YIL���=��_?�&�˽�>!.�>](�=���;�@���>C���JU.���>����/x���K�����>�W�>��z>p;x�L�6��5�>5�	��D���M���?�N}�>}��>��G?�n&�O�>h!?�Am>6g�����������_=�KW?b��?\�U?hW?t�~gF��ؠ=�3>��%?�?9��;����7Q>|�?�͋� ���U%�LM?���?gh�?>�T?��T�$�ƿ�*���}�☰�N��=S�=I�B>����!�p�=SW�=�`�D��=ǽ�>���>��>�>�7$>8P]=" ���H ��1��R�8�L���ľ=ᖾ������t���]���+˾�?0��}Ž����;;���$��9��s�=��2>�$Z>v��>�l8?�f�>�=��1���@���J�����x������f��Z���`c�w>���=G�Ӿ�{=�#���?>0<y��>#�!�S;�=@�?�x�=�ϼ��`>m>�>>��0����>nP�>H�c=ܲ>���> ,�>Y i��������}h���<�F?�s<=x5��N��K���s�v*�>C�	?�r= ��ͤ�����>�>����)�=�x�]��ꃼD?�>e�>+i>Ȳ��I;_>o[�����x��C�>T#�>�^=D�>�.
��V������>��վ���=�|>q)?�w?��1?�w�=��>�rL>"'�>��=ښB>oF>�V�>N�?�O;?Ȫ0?i3�>��=�_���C=�SF=?�K��h0�B����C�?���m�<�uM���A=�U=! �Í2=w\[=�)�����:0�=?9?�;N?�_>>��>4���:�s��$�a?�?���>d2?�H?��?�]>��+�PȾ��Ҿ�s�=,��>�"z>c[3��ۘ�P����>��W�o��>��R?��=����0�C�M|�>J��>���>���>���>�=;�6��C�������H�p���O�<�×������H����l�h�>�b���f�=��=�
�=�?�>��=�==�̄=��K>��>2��>"GV=�P�=$1�=r0=��N��[Z=2�=I!���<V�=��w=��G��{3�t���/;�:�������=��>K�$?���>�W#�a�t�_͚��/�> �=w���ݵ�>wj��sd�Ggd�1d9�6��В�>��V?OO>Hu]�am�=� A����>���>��4>t�>�^H��4ξ�D��=W�>��	?W� ?��>�D��;�a�/[k���$��>�>��=�@*��ɏ?+�R?�iԾJ��=B(��$x�����%��yhO�A����"a+�z<��#Ѿx����>G�~��=v��>�E�?��a���[���̾�[��U����vVe<8	2>C�.>�������$��?Ǿ�%�����9��8!�>7��=��>Pp?�B?W��?���=Ae�>ix>~�?�6�>b�`=fx�>��"?��F?�J?tG=n-.;���zM��	�+����s�!=�f��*>bb>��A>&��=�?^��ـ<�L#>a2=W0�<'�=$z=���<��=�d�>,P8>�?��H?���;�aI�
��=IJ�=�c�^�����>
�*>�����о���>�2?�<?F�>��;Vn!��h3���پu@�i0?�M?h5�>V���v�.:̾+����S�;�my>�	�=~tѾ9������=aU�>y�>xU�>�͎>�hz?��!?�E?����+(�	+�-�5����E��> �|>��->K����6� �h�(fi��8,��*>����v�=��=�}%���k>Iݍ<-��=��5>M�=�Ey���f�J]>e+�>4�?��?��=����]5��X_?�?�Ĩ��Y5��@��O>�u?��>�d��-?�aO>�C~��CĿZ�r�P�>:��?g��?2�?�x����gW�>/�>�`�=UJk<GZ��K<����^=��<=kGf�p���Sݾ�!۽
�=���>-؏��C��Ċ�˙-�o����,D��F=D?�����M�������ս�9���N<�@��vy�[dN��Q�S<�����K����E�;yՋ?��p?��;>6l����1�����־�}z=Xq��[������S��ƾ��־H�;t��B3<�y��躾Ỳ>2�P�%|�X�|�}�6���
����=��4?Ǿ��m��	���LѼG�=�N��`�)d��
���~νF+e?RF\?��龃�E�\K@�K�����"?�(? A�>(z����=��>T�$?k�-?2}�<����A�c��l�=���?�J�?�B?��؃>����#���w�>�?��>��C�m;Ⱦ	�Q?�0C?G!�>�&�􎅿?a ����>uOO?�@�!�j>��>X��>�����p����3����L$�6�%>"�Ƚ<�K���v���)����=d|�>5��>�σ�{���҅>���0�o��.\�sE�v�/=�z��@?���;��>a?Nnv�����!��c�����'���+?�j�?IoA?g�q?����av��7�w=�?d_B?	�x>�]��>c�?�'����t�wv�����>	��?y�?��h?�@%�&Vٿ+���-���t���]>J*8>�{�>#�C���=�=�M}��&�}�>���>�]>�*3>PO!>�(	>�V->9����A$��X���,���.�\
�������J��R���f����n����Uc�S�[�5�o!�k���p�t�/�>���>w'?�"3?9��!��=�����^�F����a��������j��Z�K��c���]=ãľ��=�"�{L?i�=�=�=&!?�A��(����>a�>�=�9�>���>��>nB�|0�=2>=>*�Y>s>�>~V>�+}�"f����'�W� N�<�E?v�)��QR��>������f�TĚ>�:?&?>��2��j�������>V��(eQ��
;�Lu%�C<>{@�>_�=��˼ah����~�$��9�=�փ>+$�=�0<�ym����m�8�ȱ�>}+Ծ��=<�}>]�"?Vy?�,?�7=�M�>�&>3�>qH�=��%>��D>�4>�?G;?�R,?P��>-��=��d��y=�5t=��?�S�v�-���1�Q�
����<��[�o�J=^�=Tw�k�<�4(=I���:��<M�>-k+?�r�>�,�>������G�G����>�QJ���>cD>DҔ>xZ?�{�>'�b>>/=����!W�=|m�>˥�>�RD�	K��N;����>::-�E?�F?+��ӵ��k��A�=�X�>E��>��
?��L>E����(J=H���޿C��~���<c��#��=�༺�m�(9�=T�f�r��]�=���>v>�>�Y>�>��6>*>zT�>b�\>��/>�I�=�;��n��V��������$q�*�:q�=�<G�D3r����=���<�$	��D�=���͘?�~?B'<I_=�T=�	�� 6��Ќ>�9�>?�
>)��>a��+w˾C��qX�,�*�� ?�N?��>
	��T�=*������=%pz> �;���>��������T��Q?�>*��>�*??��>��q��Ut�NE��6��D�v>Y���HW��Ȍ?o�q?0�龜��v_��Z���L���F��ƽ%�c�񕧾�K"�}dB��[Ⱦg-���Q���>�f�>���?N�6��%>��/�Z�y��k����Wz>X�[>���>@D��E�����ٰ��E����<X��<G*?Q�>S��>~pA?�'?e&g?��=q��>9��J�'?(�[>��e>��F?P�B?��T?d�:?�!��x�h����H��ؗQ�Sw���Q=��=��=��K>=�<>�Ӣ;��뽶V���+>��<\Z���q=r�&>Ӆ=�ђ=�Kf>j[T>o? ,8?5¥��(<��"�<��i��֍4>_��>��=��^��}�>��>��?���>a��;I��Kg"���+��;���>I5?��
?�|Z�����*��ځ(���;�IK�>W�V>t�#�b���w�u��~�>�<�>x��z��>~ty?�=2?��? ���r:�o�`�"�+�&�S<nPU�ݿ>�D�>��>�����:��=t��N`� 1.�"��<��;�C;;=e��=\J
>��>�T�=~�o>��U�U��@�����t�L=���>M��>�?�o4>6O�<�t����ᾊ�:?X���rn�MĚ�_-���=�G?�*�>[WW�qp.?�u=pTq�bݮ�n[(��I'?!f�?�u�?R�m?P��=�h�Sݼ>I:�>
�>!�<�|;3�(���h=R>~�M�g��������=ҥY>��>T.B�@����9��5��h�ʿo^�X��=�͡�����
��B;۾���h���7�d��$���&��T��rj��7;�cs���˰�����ď��?%�?們?	�I>�=hg������-�#ԑ�m�}���Q�.@~�Y(�ٕپE44��\�+��'=�-!4�q�Ǿ��>��Y�둿_�|�b�(����E%;>��.?�0ƾ�a��=-��^=�$>+��<������Ŝ���$
�D^W?=4:?�C�H���2彝>�?�M�>#(>I���\���d�>��3?��-?��鼊ڎ��ȋ�!��}��?���?��W?3�8>_y�2]���n�$?��>�>2a�=�S���=�??=�c?��?q���[���{Y��l'�_a?EX?���>.�>:5�=R��=��۽:��=�&���K�n�>3�þ��r����0���_>���>�҂>�y����<��0�>K�ܾȘ5��h��8�a/���=p� ?Ոξ��>Ly�>�<������:����Ͻ�
9?\�?\K?Q�z?�,�t.f�M� �ȼ=�M ?f�F?�d�<^��D��>�#?�t۾�W|�������>~��?e��?�a?�C�hu̿�T������楾`��=0� >�8�>==������=��C>��~<��u>:��>;	�>CKG>��>��>��>�}����e����K���kK�>V*��N���/@� �%�\�a���4��zp��wN;񘓽�=���gڽ�d���}�޻>ȩ�>O��>qv�>ҽ�=l^�>�y�<2b׾O���0�����,�@����,��(������	!�Ԃ��e�����'��� ���:?�H�=�@�<��6?��e�Y~�>(��=_�=�$b>�2=�Q�=:�<Eѵ� 1������f_>'/�>E��=�傿<���/�D[[��(*<�A?�D�����&7���Ծu����X�>'F?��:>w2*�ꠕ�ȡy����>IK��{P��׹��!��T�>>�>�w�=a"�;�(������s���=�~>�v>�'��󈾒:�w�=WN�>
=ž5t>��l>�#?	�|?�K&?��<<Q�>�)>��>�:�=G>"{>�&z>iE?9s=?3�.?�(�>y�=5L�S��<��;4������`ȽD�}±�^�X=�Ò�6k�=��=����	=��(=%�d�ǂ<��<���>��;?�g�>
��>#�������mP� 4Ѿ��5>� ��xJ?dͧ>j��>�?��~>�k>0K���ߡ���P=�>Ϗ�>^NF�8������=�ۀ>6�>$�'?&b'?C��=Bsg�|MR�`��=��>V��>i�0?�1�>���=���JL��5ݿ��P��<@��G���+���>����x��n����v��s�<���=�G�>�Qo>2u>��L>�s>[�F>�>
6j>�Y>8�=4�=�~�=����/�r!S=�սK�W����<�P��!�2Z	�q��?=���<��<h��>��?Ϫ�=Ps>���◰��4��㱼o��>��>O=>X&a>�����P��xn�����y�?;pL?X�>8L����$�ͺ���>U��=���<u��>���>��g�n�x��o�>�j�>�fm?� J>H�ܽ��f�ꩉ�4A��� ?.;=Z�J�DΟ?-N�?�������r�n�y8�eya��n6��6m������ 	�S���Ͼ7֢���c�=A��>W��?N#Z���=���\�V�׀��x�)�-ɺ��%��Y��>���=c�Ͼd ̼
�Ͼd,׽�N�=���>�z�>H��=��>9�C?��?�I�?_�6>h��>���=+?p�>�J�>�.?wy7?�S7?��"? �����ٞ�X����0�vx����=�z�<Q
�=m"�=l�8>'t8=�f7���=)>?;=[0��ӵ=ҷ(>�B�="@>$o>�>`?<�"?\�:�*ƺ���[>������W=��p>�cG>rz-=�/�ŗ!;��r>#��>\�#?餁>&�� $��;��h�f>���>�,?(�!?������G�L՞�$k�r����ç>�{�=V�Ľ�����,�9��颀>�9�>8p#��)�>�dj?�?,)?��ｱ�!���N�IS���m#>�����>~�?��>Z4оg�H�MA���l��
����>Lt��E>&��GL���>wU�=�t>�'u=xv�=�s�&6�=�IL>d�>�X�>�J�>r}�=N�	���ھ����F�M?p|�N%�%���c5���>�ʱ>��=�ј���)?憴<����oڦ�I���t?QI�?F�?�L?�w��? �1|>2�(>�<>�j�y*Ǿ2���r=�Rn>G�=�������4Y=I;�>w�>
�m��ľ/���)Y�X���2�B����/uǾ�׉�����(��g��쉂�,���J���8%�����~��zս���.����銾<U���[�?�U�?7u>kÇ���W��D���(ݾe�>6�N�Z$�����Sb��y5ʾ@�Y���D�6Z7��!Ծh�����>�sT�����(Tz�͕)�Q2%�\�>r1.?�þBP����R=(�#>:.<�����&i��s���W?�??s�྅=�����=��=�?gd�>u�>>$��4敽}��>V,,?)&?�%a�v᏿r늿�����?�<�?��D?dW=�I7�͚%��;��x�>��?p�>/.�dr���1��?�PV? ��>�۾]���!K�9>��C?#?-�ñ>>{ж>�p;>�[�=B������% � �ν��v>VY���䇾�@(�9�8���>��>�Z�>�J���;4�&L�>p���������T8M�M˨��p ?��U?� i��t����&?�=�>�������2��.R�<�w?��?nA-?iW&?��������=?���u�;�=?��O��Zr���~>�i>��C��>��q���I�>���?7�?ob?TO�/5ʿ�����n���܉���L>[s\>ܪz>�~?=#5�=M�=ȷ��2���r>ڛ�>֒�>��>	K>�� >
ݥ=	b��:����\�x���wؾ<�*�"���ľ��u�k��3����ɾ*S����.��C�G���Ϳ��j�1=�lξ$*�=;�?r��>�ξ>�nG>��=8Ɉ��)��O�b�ƾ>�&��6�'�پ1�Ǿ^c����� C�� ���<^�о���>m ͽS��=�>�ν��>�4�>i�>�V>�>���>X�[>��>�F=��>ޭT>{J�>��z>�y�=�:���I|��R4�I>�^Ǉ;wwC?TJ����,�z�����K�>��?n^t>���ޓ�u8z����>��'�Q�h�A���b���>�3�>8�=/)^<l�L����|o
�2��=�ʆ>�\>�x������ǽꏪ=GO�>�����>�|g:��&?B��?�j9?j)����>Us�>�j>�^�=��2>��q>zS>�, ?�H(?w=)?���>,b�=tp��%�>J�D>8G�������=��:���'��= ~�:�q�>lā��
h>(P�> �ݽx�,��+=���l���>k�/?c�x>8�?��E@�R�7�W0n��>t笾�t�>�t�>�+?(9!?G?�Ǚ>T������6�-��>m9>E"]��8e�K�5��A�>ys�>{t`?0�$?��6��ꀽ/3p;�"��m�%=n)>U?��?�7>}�׽��Oǿͅ��s���'>A�h>؉_=~�g�cwb<eJ�� q�����\cD��q�d/>Lt>��<>m<�2>��>��>[>�=�H�=G��8�<S�۽"X�|	�5���R��)Ƚ�t��������Ԟ��@+�������j���?V�?��=��	��P�[�
��-\�N�>�_�>z/3?�	�>o�z=SM7���Z��U�೸=/h?���?�.?�Q'�u>F�=��E=�|?,R�>���!�(�"�b<{]��3^�x��=�?��>.g�V����V��8�kp�>�Z�=�KO�e4�?.%i?+3Ǿw������N�zK澺g�������3۪�\(Ͼ9� ����F�y&[�'��͌�>0��?h�־��=
@��a������1Yc�T2>F׸�ZŜ>s�>m��0��b�B����Ǖ¾ֽͧ 6�>�8�=r��>��?�"?1by?��/?��>�,���	?*�G>���>1fW>���>�	�>�Q�>a�>��v>���=�d;������>=y�!�>��o>�N>��<��O=���=Nm�=�8=�Oż�uX<�a=�
f=%A=8�Z=�sU>��	?u6?��#�
.>��>�<�;譽��x��>)Xs�O���Qƃ�k��>�l.?�+[?��
?��<�bf�7=����G=}��>T�?�?�e�=���=Ս�Z�0�4��>&y�<����
��dI1�C�7��%��_#�=
X�>8]>���>}�l?�%�>�c0?�
#���P�pj��(����t>>[��=��
�2H�>f��>��5>x/ؾ�����Xl�9�M�r�ཿܽ;Y˼����b->��'>�61>��D>���=(�K��Sؽd �=p���-i�>%�>�N??d�y>�y�<bZ̾�	+�ueP?ȇL��-�]���U�/��+���\�>¦�=�E��Ґ?�4=�3(�9���lD���>|>�?ȭ�?I.�?�}=����oS/>���>��>��?>���l����QL�>�g�>�ľ�
ʾJ`�;ϊ>��>Q���@j�����I�¿�{W��N��<���&�akt��I��o�	��3i���x\׾�E����������䜽���d�Ⱦ�Tɾ�N�ޣ�?��y?����	���B�$,��㾊�6>x����0=��7����$��b}�����;��[�������>��G�h��[Ä���jM��_�>=��_?����v�������ܨ=L��>�"���螎��ņ���w�}Z?�M?�2̾I�"���Ծ�_���Z�>8� ?/�?\쾢�k���?��N?[�N?�Q��R���ٔ�se>�f�?@�?.{=?C	N��nG��O��2��p�>�?��? ���~>ؾ�Y?�?�9C??j�>�
�l���ڇ��� ?�\?lO2�e�g>Y��>{+�>�,��錾C�+=�Ӗ��ʽ�A4>�}X<���Q�v�y!'�o�=�;�>�J�>�?�5t���z ?�i��'�{�6[�Dq[�3up�?T�>�E?F�w����� ?z?V� ����V���촇��D�?���?j5R?�:?D����˾A��=dDܽ=�:>��?�Qٽ,���%��>��>�ƴ����	�)�?�m�?WG�?��~?~k��ѿ�����N�ھ9I�=m�<RW>��;��>�����%>{@�=��9>���>���>Oܟ>��(>��J>�/>�k��?����������[�����Y�h<޽����ｘ	�*����켾ѝ����2H���f�X�߽u�3�v�̾.��=��?W�>U�>|l >�!J>�S��[#;HJn�aM����6����f��S\辸���\�Ȫ��'=+�r�8����>#!�Gr�=T��>�s==�#ý�I�>�<���P>�:�>�=J>�Š> ��>n�M<)=�==ߺ=�j=��}>7Ҍ=b��Ā�-~9��L���b;@�B?gi[�N*���*3�����w�>�z?��S>�~&�����evy��+�>ɫF�n_c�oν������>s{�>^�=��ܻ`�a�w�}X�y��=�ą>%�
>a�x�<��}��up�=���>�Y���ޡ>�u>;@Z?j�z?�6?-��<hh�>�s�>�k�>K��>��>nc�>��?�@)?q�?Gp?�h?�BF>� �[��>B��>�|��0��a�����V򽢦��t?&>���=i�=��C��ս�	h���ֻκ?�I?���>��?6�-�l��FL�d犾���=��|����>5��>�u4?���>:b?Y�U>�<��;��=��Y�>'��=���@=���R>�h?jW�>j�2?�!?gw�<�)�=A(�CHB>5i�> ��>�?��?�4�>ì�����JW���X��f��Q��3�0>��x>C��>XM>��A>�ݽx���-��6>�gh>�}�>����-ȭ=HB�=o��>9gp>"N�>��=�Ǡ=H��<�e�y�����ow=F� ����沥���%��1(5�����ཫA����>I	?"|�<��=�J����,�>�?�S	�>}>��?�+�>�y�٪@��Lm�ZrF��E���?Eg?�y?�ݾl >�=F�Y��S,?�`?��m=�H>���=[���j�_=�>I�,?c�>d���4;�.}��U,���>�w=�t�����?�1g?��Ͼ.���X�A~x��(����=Np��Gpֽx�Sﾜ�'�e���"�	�`�c 3>3J�>���?i��4r��y�ʾSӝ��֤��Z��?�>�-ۼ�8�>�H>g($<L$���`j�ٓC�e����4���>p1I>!5�>O�?8r?+��?9@D?T�?08<��?2��=�d�>x��>���>]?2�-?[�>`{>���=��2=pO�p]�����=���<X>�	�=H�>��A<(+<�������dBB=���=��b�E��I=هU>G?7>@� ??U=?�	��
	>�<>��=���R3=W_Y>�(��]v�����!�?��?�1?�Qc> +=��A)T��yؾ��=Œ?�?���>E���� >B�����vū��qN>{�='��U�7�-:�<mL�=�T���,�>���>C��>�͆?D�;?��>;�4�yk;��Ԟ�e�X����>q*��� ���?A�>�|�<1'�(mu�նT��s�����i��� (=�s�{½=Q�켒�.>O�>g��<m!����=�>��9b�>(x?3�?)q�><�s>�W��u-�&Z?�����y�J/��8���2�>q+>^����?�]�=�dI�������y���=���?��?#.�?�~��-c��np6>y��>���>Kk=ر��Gn��l��w۪>M�>t��k��M�.�&��>��E>��&�{����(�O�w�B乿��L�����¾%�}�z��(���N�C�\�7 l�}��&�����:�&�I&�I�T����o0�������?��t?Ѻ�=�|;�U0��q׾��Q��#��1�I�v�"�g����þ���j���������x�>��9�P
����e�!5����8�=��B?L�޾��ؾ@#۾V�]=�׈>��{�\��j��������P.�
�z?�O?�.�,��F¾K7�; ]?�?��>�x��Ŷ�ʨ�>r�G?�
]?޶�j��7��B؛�O0�?�t�?��??N���A��$����*�?�S?	��>�@����̾5���
?�!:?=�>f��@*�����X��>�[?<N�!vb>���>-�>�R�%{��I��m���
����:>'s��L�X�h��>�.�=+�>R+x>�~[�������>�S���"��Z�[���^�[u:��qw9��m?��I�ž�6?�wZ>��M��׫��4���_ ��|?�c�?�9^?5I?�{þ��?��:���7>6)�>
2�>�^>꾸����<��?L־�m�� �Bu�>L��?��?��?c'�
�׿[���]ݯ�����=�j�=Ko>>�AI=�C�=]�C�	����=.�>�
g>��[>B>��2>�N<>k	�=q7������;��H��i�3��s�7T�DV�����O�6o�>����;H��%���1ɽ�3�$;�n,��� Ǿ6�3>v�?|h�=�Jo>�f�<��>�ӏ�:e�����崾�pK��- ��7���ܾ��� ���� ��g
�j�=�)2���>����.�=(&�>��e=ǘ->���>�4��_���ɰ�>f�>LL�>���>Wo= �=<��>⥇>���>?� >[9��/>�� �@���;�l �W�*?�V����֬"����"B�����>��?�eD>�V%�b���{�����>����sd��)��p�ٻ�Zv>�J�>�=� ��z��Ѡ�헽� �=�Ah>��%>���;�(����!��}�=v�>���P_�>걄>��$?�m?>�I?Ow<-K�>��>`�
>&��=�;;>~>8/�>hk?��*?A�0?s�>�� >�Ȥ��`�:U^->�4e�����Խ�j��κ��ۉ�N�?�6
{=�i>xx>PL���+��m5�r��;�<H=Z�?rb?�i�>��[>SV�1(���Z�~%徘"�>�&�)<?6JH>�t�>�a?,ܑ>����D�4�����/��X�>�[t>�>q�1A|��VǾ0W�>�W>Z:?�^s?Nq�i�л��</#�>�>��;?�-5?k�>^H���O��$���ȿ�i%�E�0����<5:��%��<33�'甽Z�>�kT=-N��6��u>��>�>���=WV�=c��=���>�>��=k�$=��-=�Ҽ�s]��R��Bk= �{:ܑ&;}Y�mG���Y�]��H����E�߽J��= b?�� ?\X]���E��8���3��/оV�?g�$?�-?�\0>�F�>�=þ$�D� �j�w��7�%>��!?�\+?��j���f>Kv�iH��3�>_1?�s>L.o�����Y��P_�=�E�>@=9?��>��8��e8��r���"�!<�>��= v��x��?OI?����=�߾�����hܾ������T� am����(Ǿ�5)�� ����0/e�ap>q�?��?��վ�νg��☿����A_Q=�
�>h>���z>�k�>��s��"�n�O�3m+���о�:�Te?2�7=����A?�Z?\9�?�c�?��G?�_'=�>��>d�X>8�&=E�	?(�>_nb?nS
?Ե,>�A>�7�<�����f ��L��07�{�?��f=���=$�=������Z=au�<��0��b)�����v�=:=�X�=�+�=��$?M-U?k9t�g�m>�OӼI�s���B=�ڗ���>�־Z�
���==1�?^G/?��F?b30>�x��n�)��0]��?��3�T�0?��q?#xa?Ak�{ZC>{�㽭?ɾ���=`��=�\�x���w3�wދ�i���to>5��>���>�[y>H�?#�-?�+?��]<Q�W�\�W�"�:�J&�~��<z�?>�,>x;>�"�H(��*��N�O�?!<�/A����2�U��=J�Y>�r=�0N<N)a>9�d��]���-
>ݛ���U>�n�U��=���>z��>�|>�E�=�ge�4'$�y�Q?^N˾x�W>`�����S��M����>�.�>��>��=E0����Կ�������{��?���?��?<���<�Ht>�?@�>J�R�R����>����:F�>��?�r�����d��=��>��=,Ĕ�"���m*�ډW�"���h/$��>�y�����O�o;�zd��I�e��z�$���Z_���m��M�;��e�k���̾<ݾ�����?	Td?N�>���=�k�v
!�vc��8'=��˾�Ε��S\��>�aP��[E��(������(��m��%̾��>��&��;���t���.�ɇ�����=��,?���L������~�=w�='g�w��?���l	��az�b�[?|VE?��߾Bl���I��_=q?���>ڽL> [���̽S��>��4?Z�*?Q���;_��/S~��O�=���?���?�`?{�>�M���s�2����i�>B?�����>�B�=,O����/���p?żX?���>�iN������o�G����܁?�D����=j��>>^�>�ȥ�<d��|.>�DǾ](�} D>u���pNܾ�u�������>g�=a��>.x��oM4����>�ž���Rd�0�Y��G�\0Q=fH�>N�9��1N�v
?��>2�_�겿,%���[��-f?�¯? �f?��0?O�žD�?����>�:��¥�=D��>���ի��Zy�>C�>w��R���Y�3�~�?�t�?�N @��?𖂿`ݿ�P�������- �w7	>���=f�->'W���>^>�,=dP:;�	>u�>H�>�I�>�?7>j��=�>&����9Ӧ�1�����F�ѩ�}Jо|�y��堾�{v�3/�A���.#ľ�R\�Ã�<��4)9����v�S=��þj��=�?��>�?�'a>U��>������*������<�"���.��EV���&n��	m� �����Tjb��LT��?�9��ͧn>J��>���=��=EIK>�}��wc>u@�>�%W>.��>D��>��>�	�=}]d>�)<
0m>�l=������|���<�Z�g��h��w�??XXn�f ����(�م߾�N���x>U� ?�@>�g)�2̓�K-w�7��>��r�k���u�ڽ!8Y��M�>{Ż>m��=��<���B?v�ҧ��%��=�M�>��>I�-�������&�C �=�>!BƾFD�>�v���t�>g�?9[:?�f�>R`h>{�W���ɀz���>g(=)B ?��B?y�e?Me�?�*T?���<�JF�7��=�'�<sy�O��<��Μ ��챻D!R�<-�Iނ=���=�8==�:���˻h%��w(�=�7>��?L�`?,:�>�f�>�.�<,r׾~�C��6ܾ�S�>)"5>S��>�{�>ó�>)��>�Z�>G��=���<?����!�U�>�>��D��B�B��e��>��=�n-?��?�g�=��>bv=��4>�cg>�_?DG>?o�>�>Y=]��&�>ο=V��슿R�k�FB�=�r>�4�>�?��P���7��
�!1]>�f�>�,�>m7�>��=r�S>'<�>���>D>�=�6O=ƹ����=\�&=Y�>R骽H�"�
�u&�����=��3>׬�2!�]&��>�uj�D�>��?��	=��=�⑾���%���.`B>R�>�`�>+�F>�������k��sI���G����>�H?T��>�Ⱦ�z>���>+�o(?}�
?���>��=��_�]���V��p��>'�8?�3�>����!n�%_���@�[�>@A�y�����?�5F?vVؾ���zT�F�/���/���<<��������Қ˾ڑV�y�N��qM�|���A��=��
?�Q�?QR;/9���㾢	�����#����j�>J�>�V:?��?������J�Z�و��fȌ��D
�S�>�8>7Y�>�?�G4?C�?� ?41?yɕ=��>^@Z���#=��9<�=?7�<?��<?�A�>:_h>�1�=����2����t��y{
�Ӊz>G0��C$��:<>l}d>V��=�z�=�x=�R%�Ӕ>�C�̫=+�A>�8>�S�>J�/?MG?��D>�>��v�C*z�n�\��7��.�x=�φ=L
>�c&����>��>d�'?��>�O�<��!�	�[����=3��>�		?�*?��x=���>�}����Bm]��휽����{"��%t��2��C�<�f�=���>^�=�P�>�%a?�� ?Z��>��=Ծe�ȼ����1��ý)��>��?0V?s�=6`#��D(�{�p�OHV��O�𺇾�7�����=���<si�=���=��=�>h={2)�D:u��ɽ�����>�)=>G��>�3�=g,>`F�$���=l=?o"��F���,�P��\��lP>���=9J��c*0?�#8��'Y�qJ¿����T>��?^��?X_�?�h��]��Cx>��!?��>Fp��e�<�M��cӋ��/�>a�>w!�7���I>�>_Fd>dپ��^�L}B�:"������l�������!x+�L 7�B���}��=��ِ���+�����4� �6��=`Ľ5 Ⱦ(������=��Ձ�?�AA?��m>���>�Y⾌���m	�x�s��#�����/M��\ǐ����U��� �N?�x	/�Y�9�;=�u�i>[U���F��W�h�f�G�5������"?�Һ�C����{�=Q�>�v~��F3�8���F䘿��v��yk??C?� ���-7��nϾ��=|'?s�>�\�>����,zľ,��=2
@?N�+?�U�]ˎ��n��:=Yǲ?���?�??ԄM��5A����4���r?�
?�-�>����̾z�콑�?��9?ݍ�>#���d��a^��W�>�5[?��M��[a>X��>���>���m=���R��E��|ɐ�?9>����'���i��>� C�=�D�>�Px>��\������z ?�i��'�{�6[�Dq[�3up�?T�>�E?F�w����� ?z?V� ����V���촇��D�?���?j5R?�:?D����˾A��=dDܽ=�:>��?�Qٽ,���%��>��>�ƴ����	�)�?�m�?WG�?��~?~k��ѿ�����N�ھ9I�=m�<RW>��;��>�����%>{@�=��9>���>���>Oܟ>��(>��J>�/>�k��?����������[�����Y�h<޽����ｘ	�*����켾ѝ����2H���f�X�߽u�3�v�̾.��=��?W�>U�>|l >�!J>�S��[#;HJn�aM����6����f��S\辸���\�Ȫ��'=+�r�8����>#!�Gr�=T��>�s==�#ý�I�>�<���P>�:�>�=J>�Š> ��>n�M<)=�==ߺ=�j=��}>7Ҍ=b��Ā�-~9��L���b;@�B?gi[�N*���*3�����w�>�z?��S>�~&�����evy��+�>ɫF�n_c�oν������>s{�>^�=��ܻ`�a�w�}X�y��=�ą>%�
>a�x�<��}��up�=���>�Y���ޡ>�u>;@Z?j�z?�6?-��<hh�>�s�>�k�>K��>��>nc�>��?�@)?q�?Gp?�h?�BF>� �[��>B��>�|��0��a�����V򽢦��t?&>���=i�=��C��ս�	h���ֻκ?�I?���>��?6�-�l��FL�d犾���=��|����>5��>�u4?���>:b?Y�U>�<��;��=��Y�>'��=���@=���R>�h?jW�>j�2?�!?gw�<�)�=A(�CHB>5i�> ��>�?��?�4�>ì�����JW���X��f��Q��3�0>��x>C��>XM>��A>�ݽx���-��6>�gh>�}�>����-ȭ=HB�=o��>9gp>"N�>��=�Ǡ=H��<�e�y�����ow=F� ����沥���%��1(5�����ཫA����>I	?"|�<��=�J����,�>�?�S	�>}>��?�+�>�y�٪@��Lm�ZrF��E���?Eg?�y?�ݾl >�=F�Y��S,?�`?��m=�H>���=[���j�_=�>I�,?c�>d���4;�.}��U,���>�w=�t�����?�1g?��Ͼ.���X�A~x��(����=Np��Gpֽx�Sﾜ�'�e���"�	�`�c 3>3J�>���?i��4r��y�ʾSӝ��֤��Z��?�>�-ۼ�8�>�H>g($<L$���`j�ٓC�e����4���>p1I>!5�>O�?8r?+��?9@D?T�?08<��?2��=�d�>x��>���>]?2�-?[�>`{>���=��2=pO�p]�����=���<X>�	�=H�>��A<(+<�������dBB=���=��b�E��I=هU>G?7>@� ??U=?�	��
	>�<>��=���R3=W_Y>�(��]v�����!�?��?�1?�Qc> +=��A)T��yؾ��=Œ?�?���>E���� >B�����vū��qN>{�='��U�7�-:�<mL�=�T���,�>���>C��>�͆?D�;?��>;�4�yk;��Ԟ�e�X����>q*��� ���?A�>�|�<1'�(mu�նT��s�����i��� (=�s�{½=Q�켒�.>O�>g��<m!����=�>��9b�>(x?3�?)q�><�s>�W��u-�&Z?�����y�J/��8���2�>q+>^����?�]�=�dI�������y���=���?��?#.�?�~��-c��np6>y��>���>Kk=ر��Gn��l��w۪>M�>t��k��M�.�&��>��E>��&�{����(�O�w�B乿��L�����¾%�}�z��(���N�C�\�7 l�}��&�����:�&�I&�I�T����o0�������?��t?Ѻ�=�|;�U0��q׾��Q��#��1�I�v�"�g����þ���j���������x�>��9�P
����e�!5����8�=��B?L�޾��ؾ@#۾V�]=�׈>��{�\��j��������P.�
�z?�O?�.�,��F¾K7�; ]?�?��>�x��Ŷ�ʨ�>r�G?�
]?޶�j��7��B؛�O0�?�t�?��??N���A��$����*�?�S?	��>�@����̾5���
?�!:?=�>f��@*�����X��>�[?<N�!vb>���>-�>�R�%{��I��m���
����:>'s��L�X�h��>�.�=+�>R+x>�~[����C�>AC�s"����i��>���>�-s=�F	?�Ҿ˔�ƙ�>��>�+Ծ#���<���N���Q?�5�?zp?t�2?� ����#ؽ;]�=r~�>���>��3���Ͼס�>U�=>w���·��6��7*�>���?� @�6^?�����Kѿ���b��VÇ��<#>�= �f>o���2�=#*B�O;�m�!=3]V>�9�>��>��d>]hD>2`H>�>�D���2,�0#���א���;��!��5vf����DM��tD�����'Q��(�ս��潰㿽��X�:�#���D��d���+<I4�>rm�=)��>?	�>X��>������}-�\���>,�s���72��ܯ���� 곽�����4�:�d���i�>,�����=p��>�h=�d��?hN��9���3>$g9��]>L��=c>�=��g���=�fy>N��=Dz�����o�8���J�VE< C?0�]�
Μ��4����h���T�>s�?=�U>��&����J[y�C!�>-�?��a�N#ƽ�(�fX�> ��>
�=�{�9�	� `z��&� p�=+Z�>��
>o�a����#ћ=.��>�Ծ^�=��`>��(?��w?d�6?Ι=���>�2>���>$7�=�a9>��F>v��>t�?M�6?��,?�>M��=$rT��/8=dI�=�Q�uƊ��$ͽ��C�3|ʼt��<V�h��I=��x=f��<	�_=UjE=4y�|���X6=��>��8?���>I��>=�5��>�*�L�>V���>=���z�>���>��? �>\��>�2>J"j��þ����F�>&�>>��^��x�X���F{>��v>,?O?]�1?��g��c�=9��=b�>�=?�N)?:�>,�>J-������lӿi$�^�!��삽YI�^��;/�<��M�@��6Ȟ-�����:��<H�\>$�>N�p>�E>R�>�:3>\R�>�HG>:ӄ=�=Y�;>N;��E��M=?�OHG<��P�����$Ƽў��m���I���>��A�/ټE?�.?wJݼ�읽�Y��5쾦W�����>��>�c�>��>Ta=\[��(P�xt9���*�q
�>��e?S!�>�L��ݤ=X�ɼc�<�8�>���>�>s�սZ�u&��&��==J�>f#?���>�kL�i�]��}o�'���-�>,��;2����?;U?����?Â����+�C���Ⱦr�żu�+���O������S1��Iݾ��냲����<Z��>�j�?�gC��e�>m޾h���z��R ��$(�=��>^� ?��>��.�Y����%%�_�ꉾg½O{�>zmt��>\=??�10?٠�?���>(@A?�o<��h	?߸\=ۆ�>pZ?_�;?�
K?��8?ޓR������e��v����_l1���R<��LJ=��!>��9>����7Lk=\d�=����ɻ)�g>$��=Z�L=��<>��>�i�=�C����?H�?�oн��]��h��
�&.�<�>��/>��V�{|l����g�M>I ?T�.?��>S<�=� վ�,�9[����=o?X�-?�c�>���<��=:���Aj|���\=��_>�7��(}����F�����ꌀ>9��>p�=���=��?5�<?@8Y?�n�=�sv�^}�D!G���1>js�>)�"?Wq?��u=�����,6��~�YH��CV��A>:�5�&��d�>���=�R�>(t�=Etk=���=Tق��@$���F��L�<|	�>���>J�>5�+���ɼN�ӽ�����]x?����LC�+`��!���=D>�>@��>`"�M�>�D�i���Y᡿)!޾t�?��?��?�;�?%�R��-��T)>.? ��>^�>�<��u`轓��=ܝ�Ƌ�=\i��A��	ý���>�2�>%�*�	��K��^�"�� ̿Y�:�	>�4Ծ=�s��G��Ov߾��� ��<v�O�a�y�����������dT�A|����ھ���V��?��?�����P��C5D�
��NW�����=�U���1�;��Y��'h����~꾒 ��]��k0,�qG�>�k���=j.��ŉ�{d��@�0������^�v�(?��н������=�%�>Re��9z�9���ϭ��A���.y?B�h?��ӾiyO�C������	?�t�>{��>��x�$o!�Z	�>[??� $?����������g���<���?uE�?Y�??��O���A���=��W8?*�?N��>O݊���̾�S��?��9?��>���`���2�c�>:�[?�_N��pb>.��>5#�>���磓�]�%��E��7ȃ���9>�.	����Hh��3>�S��=��>�kx>_C]�\��C�>AC�s"����i��>���>�-s=�F	?�Ҿ˔�ƙ�>��>�+Ծ#���<���N���Q?�5�?zp?t�2?� ����#ؽ;]�=r~�>���>��3���Ͼס�>U�=>w���·��6��7*�>���?� @�6^?�����Kѿ���b��VÇ��<#>�= �f>o���2�=#*B�O;�m�!=3]V>�9�>��>��d>]hD>2`H>�>�D���2,�0#���א���;��!��5vf����DM��tD�����'Q��(�ս��潰㿽��X�:�#���D��d���+<I4�>rm�=)��>?	�>X��>������}-�\���>,�s���72��ܯ���� 곽�����4�:�d���i�>,�����=p��>�h=�d��?hN��9���3>$g9��]>L��=c>�=��g���=�fy>N��=Dz�����o�8���J�VE< C?0�]�
Μ��4����h���T�>s�?=�U>��&����J[y�C!�>-�?��a�N#ƽ�(�fX�> ��>
�=�{�9�	� `z��&� p�=+Z�>��
>o�a����#ћ=.��>�Ծ^�=��`>��(?��w?d�6?Ι=���>�2>���>$7�=�a9>��F>v��>t�?M�6?��,?�>M��=$rT��/8=dI�=�Q�uƊ��$ͽ��C�3|ʼt��<V�h��I=��x=f��<	�_=UjE=4y�|���X6=��>��8?���>I��>=�5��>�*�L�>V���>=���z�>���>��? �>\��>�2>J"j��þ����F�>&�>>��^��x�X���F{>��v>,?O?]�1?��g��c�=9��=b�>�=?�N)?:�>,�>J-������lӿi$�^�!��삽YI�^��;/�<��M�@��6Ȟ-�����:��<H�\>$�>N�p>�E>R�>�:3>\R�>�HG>:ӄ=�=Y�;>N;��E��M=?�OHG<��P�����$Ƽў��m���I���>��A�/ټE?�.?wJݼ�읽�Y��5쾦W�����>��>�c�>��>Ta=\[��(P�xt9���*�q
�>��e?S!�>�L��ݤ=X�ɼc�<�8�>���>�>s�սZ�u&��&��==J�>f#?���>�kL�i�]��}o�'���-�>,��;2����?;U?����?Â����+�C���Ⱦr�żu�+���O������S1��Iݾ��냲����<Z��>�j�?�gC��e�>m޾h���z��R ��$(�=��>^� ?��>��.�Y����%%�_�ꉾg½O{�>zmt��>\=??�10?٠�?���>(@A?�o<��h	?߸\=ۆ�>pZ?_�;?�
K?��8?ޓR������e��v����_l1���R<��LJ=��!>��9>����7Lk=\d�=����ɻ)�g>$��=Z�L=��<>��>�i�=�C����?H�?�oн��]��h��
�&.�<�>��/>��V�{|l����g�M>I ?T�.?��>S<�=� վ�,�9[����=o?X�-?�c�>���<��=:���Aj|���\=��_>�7��(}����F�����ꌀ>9��>p�=���=��?5�<?@8Y?�n�=�sv�^}�D!G���1>js�>)�"?Wq?��u=�����,6��~�YH��CV��A>:�5�&��d�>���=�R�>(t�=Etk=���=Tق��@$���F��L�<|	�>���>J�>5�+���ɼN�ӽ�����]x?����LC�+`��!���=D>�>@��>`"�M�>�D�i���Y᡿)!޾t�?��?��?�;�?%�R��-��T)>.? ��>^�>�<��u`轓��=ܝ�Ƌ�=\i��A��	ý���>�2�>%�*�	��K��^�"�� ̿Y�:�	>�4Ծ=�s��G��Ov߾��� ��<v�O�a�y�����������dT�A|����ھ���V��?��?�����P��C5D�
��NW�����=�U���1�;��Y��'h����~꾒 ��]��k0,�qG�>�k���=j.��ŉ�{d��@�0������^�v�(?��н������=�%�>Re��9z�9���ϭ��A���.y?B�h?��ӾiyO�C������	?�t�>{��>��x�$o!�Z	�>[??� $?����������g���<���?uE�?Y�??��O���A���=��W8?*�?N��>O݊���̾�S��?��9?��>���`���2�c�>:�[?�_N��pb>.��>5#�>���磓�]�%��E��7ȃ���9>�.	����Hh��3>�S��=��>�kx>_C]�\����
?�Ǿ�����pW�����	>��<���>�+ƾ�^�<�$�=m��>
�M�rH�`�����=��_?R�?7��?.�5?���k�X	ǻ���=�f�>�ݟ>vd�=�Tʾ���>Gs�>��"�@;����;��>(��?��@,��?�+��6Gӿ��������<��=3%�=�>>u�޽�ɭ=�K=:ɘ�)Y=�~�>���>?o>>;x>t�T>ޛ<>��.>l�����#��ʤ�2ْ��[B�� ���wg��{	��y�����ȴ���5�������RГ�m�G�Y��xT>�h�;��%9>U�?�.?J��>����k�5<,�����澏���X�0���	����{���=��G��G��;���\�&�۾���>�xټ�R>�??Ҍ<~�@;t?~>ّ�=CG{>��>@��=ϊ~>t8^>}��>��G>;L6>S��<#�x>t)�=�Մ��i���<���S�3Y�:�@?B�^�$ ��@�2���޾ǩ��ل>��?e�P>��'��I���x�gn�> d<��n�+⽵()�|��>^��>�I�=��R;4�������|�=�Ո>&�>Џh������jV�=�]�>߬Ⱦ;��=R5r>^0?y�i?Og??	�K>،�>C�>l�>���=v>Y>���>�
�>=��>+� ?�8?�#�>��=�\W�Ap���9���C��j�Ҏ���R�0s��R�˼G�Լ��=���=YI�=N��=��<N��l�<%3�=$�>A�O?�>�_�>M|��P5/�E�s�ɟ�%=c>�Mq�Ȥ�>n'?r�_?V�?���>Rǁ>N�{�}"�=r/���>6{>K)J��݈�}��Gk�>������"?Ưy?�s,>�[���5�Mv�=���>�@?/�?��>�E<>x>p� ����hG����g�=���=)�>��>pL��KL)�#�Ѿݗp��>�>��E>�>*`�<�s<���=��x=�V%?*�H>-=���>��=c��<�1^=�R6=Fn��N��!�y��#x=a���
��*�"���\���m��jb��\	?6�>��G=��B�,���F����?�y>��>���>z|^�'<��<s�'�=�s��c?��`?��\>�&�������=��=���>�2�>��>�~6����=�x��i�=��>���>� �>vX�� W��j��k���2>U��=���X[�?�V?=j�+�Ǿi����J�"��m�=8,��E��J�ґ-���>�Km� D˾��n��@�<���>Bء?X?��ac:>�O���ώ�[�b��I�p�&��> >P��>w�>E1(=gc�1t!�j�徭Æ�Y�H�#w�>��,>��%>�2?H-�>!`?�-?��Y?��>�u?��>���>r/?��>�\:?BU^?X =ĉ�<�Q>��<�wS�V����཰W�<�"��a�;4�R>\
>	7��.�ʽ����ֿ�<PU�;�R'=�ֆ�=ꦼ��<)�=f�=�?�H(?�����_��0�<�xί��3�C=���>k�=�*��7�<�fE>}?�7?�;�>o��=�=Ҿ����x
����<�?lz?���>��>�s>xƾ��s���*>��>=��������8@�h��mR>�7�>�<>�S�>�{?f�&?F;N?��e�ؔ���0`���p�������5>fN?��P>���={�5�RT7��Sn�(#:���H�JӒ�K*���6�1�=Dze>݁>�˼ts=\e<�n��2�f�_�%�����:?�>���>z�?��H>�=��ǚ����ʾ��[?t�`��q��M���)���=�3��ʳ>=�ᾞl�>����������}#��} ���?��?���?�$4��w ���>��?��]>H����^`<��>�<�H>6���k��l =X��a=#?M]�_��`����������d6�!�I�% վ� �;�	�g�;�S�������Bh{��eC�v̽����#�]�s�L���R���I��TA�?��?���=�!�S����$���!�6��F���&��p�g�\�����c3���۲�7z��R� ��3u���}�>�������秿�g�`�V>e8>�ʗ>��E<��O�\0��AA,>�h&>͂u>��5��Z������[	�9��?je?t ���S��v�W'�>�2#?�'�>5ݧ>�H<*bd��A�<�??%3?�X���p��"�E�=�´�?��?>W@?Z�B���L�Ʊ�D4"�C?y1?v��>�\�Ŀ޾�s%���?��5?U�>���̃� �&��{�>��s?�|8�waQ>7R�>DJ�>ZȰ�BB�����������1�� Y>��s=P�1"��ը6�*��=�>A�>��ѽ�S����?��þL�}��j���=���9 >��>��
? i�:Ͼ��=?�c�>�t�4�B�=����>l<UZ?.0�?\B?S�.?���-q����=��U>!p�>&��>Ó==�p�!�o>���>X�jb��+*����>��?M��?��[?l덿��f����������H�=��">"pG>=^ս��>���=�Qq���<^�>��>V?�>^k�>�'>1�>>��>����i'�#F��"Ϗ�!�A�_���m���8N�|���'x�A��}�����⾥���TS��=̱�1�8��*�#[=9[����=H�?ˋ�>I�>��> j�>�����ݾ8hE�*u+�
�
�?^�K����&/�/�G�ێW�(�u��~��Q�?J�5>��=�z?x.�=�?�)��>m��<[���Р�>S-T=?U�>qz�>��i>�">-=���F�{>�܇=� ���
���f:��VQ���;�C?�s]�kx����3�kt߾����M��>m�?u�S>�'�d����x����>��G�m�b�M�˽b2 �mi�>U��>�>�=�H»���a�w�V����=���>�
>#�l�e� G�bf�=��>��&���p%�>�rP?��?K��>Z�\>e)$?$�h>f��=7c{>�*`>�=�>��?mƮ>7�>�?J3�>�(Y>/.��fJ��C�<<������U��]����ܽ�q���(�9����<�ܛ��,3=�h��ե�!��<&+>�'�=�>C�D?!
?��>��'<��7��V��ӽ��{>	��<�G�=���>k=?s|?b7?�m>��	��.��*7�~۳>���>~=�$?��ݝ�=���>����K?z|D?��<�*��V��<���>��>�U�>��'?�`�>?�$>�������lӿ.$�&�!�����DJ���;��<��M��.7G�-�.���Q��<�\>��>g�p>_E>��>:;3>/R�>
IG>nӄ=��=�;�;<�E�=�M=��%[G<��P�mz��$&Ƽ������ەI�e�>�=�L7ټ�1?t�?'k�����颾�t
�Pӡ���$?��>\�>$m�>��+�e\��1Z�m�8�����J?�`?Q��>fpe��%]<��=�-�ph�>��>�>7�ͩ=��޾IҌ>��
?�|?��><7��,{g�ow�Z�!���>E7輵~k��o�?m�:?���a��9���a��! ����=.���*������z%��3:��x���yʾW����<R�>��?`Ɖ���>>��Z����؆����S�<og�>��?���>��=��龁��l��lVǾL�`�8��>���=��8>�/�>��?�?p�?�۟>�k9�7?��R>� �=��>��T?hT?h�8?���=GS�=�n�g�!����iq�ð	>�'��=>q�u>|^>��&�.�Ҏ�<�
�{�K<�~=�w�=��q=giؼ��k<c�y=X=b>H(	?	�$?M�����L��i�*���^;�2>NNc>�� ���y�A��9w>uJ?�.0?n��>�Do=,�ݾ>E��̤��P��=s�?�-?��>�V�<yڴ=Q�#�v��[�=8V>tl�:�~���ܾ�p��[�3�>��>���=Qci=8�?v=,?�@?3�A��ln��?`���J������$>s]�>��?�O�<}U��'�\�o�j�A�V�?;>[��*�=�4>�O=>H1~>x?<F�D>�a9>nm��w��b�;R��(�>^ո>X�?���=�脽�I�"���m?��¾�oH������^|�1?�>VR�>7�پ.�>�J�Q����q��W�W��>���?���?60�?�N���U���> ��>�A�>�'I�����j��!q>���
��>������\��Խ���>�'�f�ؾC���z �=��˿^�?�e<���Aߎ��ൾJ���i�ԙO�tX<<����J�Lq=�d
�.J+��D�K��K���b���?��?+E�=�b�Fg�������WQ�X� �MV�<i�X��5'�;�!����%����E3��C&�����gL;>x��^��Iی��I����d"<,��>R��+c�^H���l�=���=`�S=D��<��L͟��K���J�?:Mb?��žI��5Ǿ5�1>ڛ"?AT"?g��>n��`e���>�C?�?a�]>�`���(a��f�=d�?Cƫ?�A?��s�w�E�9��"���W?�?���>a�s��������?�7?��>2��J���G�����>��Y?�NL�!P^>���>빎>�����(�����X����g�X&>�n=4��*�z�=���=���>}2z>�R�����C�>AC�s"����i��>���>�-s=�F	?�Ҿ˔�ƙ�>��>�+Ծ#���<���N���Q?�5�?zp?t�2?� ����#ؽ;]�=r~�>���>��3���Ͼס�>U�=>w���·��6��7*�>���?� @�6^?�����Kѿ���b��VÇ��<#>�= �f>o���2�=#*B�O;�m�!=3]V>�9�>��>��d>]hD>2`H>�>�D���2,�0#���א���;��!��5vf����DM��tD�����'Q��(�ս��潰㿽��X�:�#���D��d���+<I4�>rm�=)��>?	�>X��>������}-�\���>,�s���72��ܯ���� 곽�����4�:�d���i�>,�����=p��>�h=�d��?hN��9���3>$g9��]>L��=c>�=��g���=�fy>N��=Dz�����o�8���J�VE< C?0�]�
Μ��4����h���T�>s�?=�U>��&����J[y�C!�>-�?��a�N#ƽ�(�fX�> ��>
�=�{�9�	� `z��&� p�=+Z�>��
>o�a����#ћ=.��>�Ծ^�=��`>��(?��w?d�6?Ι=���>�2>���>$7�=�a9>��F>v��>t�?M�6?��,?�>M��=$rT��/8=dI�=�Q�uƊ��$ͽ��C�3|ʼt��<V�h��I=��x=f��<	�_=UjE=4y�|���X6=��>��8?���>I��>=�5��>�*�L�>V���>=���z�>���>��? �>\��>�2>J"j��þ����F�>&�>>��^��x�X���F{>��v>,?O?]�1?��g��c�=9��=b�>�=?�N)?:�>,�>J-������lӿi$�^�!��삽YI�^��;/�<��M�@��6Ȟ-�����:��<H�\>$�>N�p>�E>R�>�:3>\R�>�HG>:ӄ=�=Y�;>N;��E��M=?�OHG<��P�����$Ƽў��m���I���>��A�/ټE?�.?wJݼ�읽�Y��5쾦W�����>��>�c�>��>Ta=\[��(P�xt9���*�q
�>��e?S!�>�L��ݤ=X�ɼc�<�8�>���>�>s�սZ�u&��&��==J�>f#?���>�kL�i�]��}o�'���-�>,��;2����?;U?����?Â����+�C���Ⱦr�żu�+���O������S1��Iݾ��냲����<Z��>�j�?�gC��e�>m޾h���z��R ��$(�=��>^� ?��>��.�Y����%%�_�ꉾg½O{�>zmt��>\=??�10?٠�?���>(@A?�o<��h	?߸\=ۆ�>pZ?_�;?�
K?��8?ޓR������e��v����_l1���R<��LJ=��!>��9>����7Lk=\d�=����ɻ)�g>$��=Z�L=��<>��>�i�=�C����?H�?�oн��]��h��
�&.�<�>��/>��V�{|l����g�M>I ?T�.?��>S<�=� վ�,�9[����=o?X�-?�c�>���<��=:���Aj|���\=��_>�7��(}����F�����ꌀ>9��>p�=���=��?5�<?@8Y?�n�=�sv�^}�D!G���1>js�>)�"?Wq?��u=�����,6��~�YH��CV��A>:�5�&��d�>���=�R�>(t�=Etk=���=Tق��@$���F��L�<|	�>���>J�>5�+���ɼN�ӽ�����]x?����LC�+`��!���=D>�>@��>`"�M�>�D�i���Y᡿)!޾t�?��?��?�;�?%�R��-��T)>.? ��>^�>�<��u`轓��=ܝ�Ƌ�=\i��A��	ý���>�2�>%�*�	��K��^�"�� ̿Y�:�	>�4Ծ=�s��G��Ov߾��� ��<v�O�a�y�����������dT�A|����ھ���V��?��?�����P��C5D�
��NW�����=�U���1�;��Y��'h����~꾒 ��]��k0,�qG�>�k���=j.��ŉ�{d��@�0������^�v�(?��н������=�%�>Re��9z�9���ϭ��A���.y?B�h?��ӾiyO�C������	?�t�>{��>��x�$o!�Z	�>[??� $?����������g���<���?uE�?Y�??��O���A���=��W8?*�?N��>O݊���̾�S��?��9?��>���`���2�c�>:�[?�_N��pb>.��>5#�>���磓�]�%��E��7ȃ���9>�.	����Hh��3>�S��=��>�kx>_C]�\���:�>`�ﾞ�J�G�q[��w���	=͒?>��W�	>$mz>@U>/�%�74��9O��r��7K?�V�?M!R?��7?a� �l��f����ϙ=���>���>9Q�=���3�>3�>-�2l���k�?���?� �?fX?)_k��ȿ�
��v��)7p�Ľ�>�	콎�>��1=��>���<�����h�=���;��>�Г>���>'W�>��>�D>1������h���}x�S�
�� 1�c��I�ʽQW.��{f�}t.�ρe�X܊��|+�?����>=�f/��K��Ծ�wu}��P>'y?��>�O�>]��= `�=�Jľ"@��e�e�����������&�ľ+�t���8���v��4������޾�?&瓽�Y�D��>��!���&>5z>BY�=WG2>��]>�>�D{>qv�>I5l>�	>d`+>�=�5�ҳ�=XA�<�O��u`�Zg��,��˻?�2�Wn��i�+�pE�_Ѿ9�>lZ$?��p>��/��{���w���X�>~Ԩ=A���gQ���ޜ�eҤ>"��>�B�=ݰy>���>\���UL��Y>f�$>&�=#e�=8����^�\�>$Q�>��5�뛃>�p>�>�?1Z�?-&�=���>���>I?���*pK>�A>Ǟr>�>�:?�VH?��>�7>n���1.=>�Uz>�>)�3ҽm�#�����RH�x`�����J]���b>'�d�'2F>�>c�|>)�;�?�<~�?eR??H?�>���>
�̽	�1�[�7����B6=T�,>��>p�	?�@�>,$%?�1?�̷>p& >�῾���ݰ>V\>p?�4�M�{�T>۟&>�z=�B?�m6?�A���=��fH>���=��>D�?�4??0�>�X�=�~ӽoO���̿��,�M�K�>�_�*���=i��P�6�h����6��@�=�?�>e��>�X�>���>���>�k'>qW�>��M>�G�=���<�x���^E>n�=*�ޤ��_���8��=����cq�}a��F���V��\�����=���=�?j\?�T)�"��E�f�4������h��>9��>���>K}�>7�=1U��U���A�7PH���>.gh?���>q�8���=��,�$��:���>�>��>�c�����F��2Ц<���>͝?a��>E��3G[��So���
�aϤ>���=�f�=��?P�d?	�����/�};~V�!�7�*��^Y�i��j޲�`Y �"�5�8(��>N��|b�qȨ=���>�5�?�Rx��t=�Pp�2��^����%���$>p�1>��>��q>��Ծ������#�E�����$��c8=��>��>O8??��9?φp?>�?Ź�>�ϡ��&?�l�>!�!?a4?�I?�K?�� ?G��>�"?^�=� 1��Eg�M�p�_�F��s�=j�=4�=_��=�vD>8��=xc�<2W�<lgK=qb�<H�G%8��,��e!>1{>iw^>�a?e�$?�2���� ����p���<���=�G>����FwT�!|�<�O[>�1?��2?��>G�=��ܾ��jq����==�?h�.?zy�>���;�=���*�h����=M�Z>	�9�"=��^��ʩ�P6߽0Q�>��>X��=��>�/�?��I?_?ț��˺!�;s`���d�y/���y=X�>��>�!�R�˾��'�`�P�WJ>�2d�?7t����ú�=�/>�缚B�[�=j��=5�=�f�;���ZZ�=�+>�C�>ƃ�>��?�x>U��:򆉾B���I?�C��"%�����_�ʾaf��.>&g=>���gW�>�����������7�;���>�d�?�0�?Hc?sl<�a��o|>��J>�<>���<�*I�KcP�˖��a�+> Ӷ=���z����2��ZW>ȱf>P�׽��о�6���S����W5�����'?��|J�������K����׾� 꾱=��x���x�����O�������	����v?��c?f7B>���;w=J�Ot��Z����4M��㉾f���o.����̻��Ӻ����D@���x�KW+���>+D�=���|;���|f��N>����4? ��=�j���9+����>e�� �(��d���V�����̋y?֐6?�Dپ��)�����Ib>&?`��=�I�>'�R�ܒ@��q>ld?nf*?=�:�=����l��$��]�?`��?X?h���H�7�i��=��y�?���>�$?1m�h��2ӽs�?�6?�*>�FW�t雿�Y0�I��>t�t?�S����=�?4 ?2�=�G��e�>OH��n���6>��>��p�/$Ӿ��T>}��=���>t��>��o��M��&�>ʓȾs>C��I���!��n��<٦?�j
��(=J�>cI�=X����'���¾v�37?���?��U?Z�?�p�	���[���p2>�һ>�T�>:�< �k�[>sx�>_�ܾ�n�����?��?`�?UP?�|���տ�ġ��4Ⱦe���+=﹉<yj8>#ç���1��g���>=��	=��=�P�>8AV>�u>��h>�Ai>���=�j��QJ�Ĝ��G��N;A�<N-�� ���{�ʾw���*0��վmJ�H�����Pڽ�d`��b�+?I�{����>�L?��>�a>E`>��G>ӎ�؝�������&��J��������	�p꾾�j��	E���Y�[��E�ܾ�a�>��>;`�>H��>z�^=%�n=�?���=Η>:t>�)�=3¨>��>E�?=#�>g'>�*<g�z>Up�=����ؑ:��1S�z�;�AC?	�^��=����3���߾�"��a�>�<?�
S>4�'�QҔ�}�x���>��E�l)c�b�˽����=�>�Z�>w��=�dǻ�z5x��Ϲ=��>�
>5zn�B*��[���o�=�@ ?^-߾����p�>��V?E	�?� e?�Y�>{�?��X>��>��_>l�B>�)?�L?>`?$T?BR?�:K>
�3>�ߠ�r��)�;i7��u�%���=�j<*9>�4x>��ν�ј<�`>�����=>Ö�=lI��9�i:lu=;�?A�*?�?�?3m��I��<�C�W�����>{r>E�>�I�>o8?.8
?��?�6�>ZB >g��6v"��`�>��p=��?�,�3��~C�� k>Ӿ�>�'[?e?[?�j����5� A�=9"�����>承>aV9?8�?|�D>��=��A�ٿ�P��m�fe/��Y�W��ʰ��,��3�=yoŽ�ؔ��MY�B>���=6 �=Q1.=�>��=Tz�>U�Z>�m>>�z̼�_<��g�
hO�3N��w�f>�2�;'���l߼�P�D�ݽ���R��q)���@=��?�@?�?.�l���xi�,��	���*��>�>
R�>~�>���=�����U�"(B��M�?��>�Sh?�G�>�g<�.
�=E*����;�X�>͟�>1R">�Ex�kl�;�����<���>��?��>�e�>�Z�fEn��L
���>�����q����?�8=?�D��%��0���K�3{ �4��=oJ���º���b,+�d-�u�Ⱦ�.����R`=j��>	\�?��+�&�����[���Z�r�J�̾J�k<Ru�/��>�=? c�� ��*�� D����&_4���=D��>��(>7.�>'�)?N&F?�??���I��>�=^?5��>5F�>\9?g],?ы?��?V�>9v�"����dL�¥�ga�=,�>�K>�h
=U`��&Iӽ���=���<��)=�tһ0w:�@�7>T	̽�J>�W>n�u=��
?`)?��T=�=w.׽j�����;A#�H�>��<E�����<�}S>�?�,?��>	/�=�e ���!��=,�>Z`)?Y��>ӹ�=�>Ru����u���.=��L>}�ͽb쥾��fs��X�J�jyY>	U�> �>&ؓ>ޚ?#hr?�>dI޾�}A�/�b��X��>f�pn'<��?���;ս���D������F�Bo��՜�a[��G��H�=��*>�J)>�?>/:n=@"�=!&��۪�j�&>�ڽ���>�?3h�>��t>>��=��0��,���I?���ώ�$�Qξ�K`>�c8>�E�I�?���N\|�;X���Y<��c�>FR�?W�?�\b?�9?�����{c>��R>��>�s�<UCK�+�"�׍��-->���=(�����j��7�U>�bs>_׫���ʾ���R�ޮ��S�5��$ =��x�;𳾄����޾���G���Zj�(�����)���}�O鶾�$Ǿ���r>ܾQ?����x?P(�?> ;޽�#�~(��O���M �d���c����9��(�|��6þ�~߾e��ʾ¾��D�?YX��e��Z>��d<8����n��*n6��� �U����%?�����Y��{��=�8�>�
�nxQ��]��wx����]�? �O?�Ѫ���_������=��q?4�k<X.?=�仉nT��]>�_t?#Ej?s(?�r0�/���L�Z=��?���?4�/?�;׻=a��qi�������>m���A�6?�*����NY澖	5?ҭD?�EJ��-�����7�0��J?Kߞ?"j���?>��D?�?�0ؽ������>�n �1������=)2*>�Ʒ��C���Ol>�^�[+3>�� ?[�,���)��:�>`�ﾞ�J�G�q[��w���	=͒?>��W�	>$mz>@U>/�%�74��9O��r��7K?�V�?M!R?��7?a� �l��f����ϙ=���>���>9Q�=���3�>3�>-�2l���k�?���?� �?fX?)_k��ȿ�
��v��)7p�Ľ�>�	콎�>��1=��>���<�����h�=���;��>�Г>���>'W�>��>�D>1������h���}x�S�
�� 1�c��I�ʽQW.��{f�}t.�ρe�X܊��|+�?����>=�f/��K��Ծ�wu}��P>'y?��>�O�>]��= `�=�Jľ"@��e�e�����������&�ľ+�t���8���v��4������޾�?&瓽�Y�D��>��!���&>5z>BY�=WG2>��]>�>�D{>qv�>I5l>�	>d`+>�=�5�ҳ�=XA�<�O��u`�Zg��,��˻?�2�Wn��i�+�pE�_Ѿ9�>lZ$?��p>��/��{���w���X�>~Ԩ=A���gQ���ޜ�eҤ>"��>�B�=ݰy>���>\���UL��Y>f�$>&�=#e�=8����^�\�>$Q�>��5�뛃>�p>�>�?1Z�?-&�=���>���>I?���*pK>�A>Ǟr>�>�:?�VH?��>�7>n���1.=>�Uz>�>)�3ҽm�#�����RH�x`�����J]���b>'�d�'2F>�>c�|>)�;�?�<~�?eR??H?�>���>
�̽	�1�[�7����B6=T�,>��>p�	?�@�>,$%?�1?�̷>p& >�῾���ݰ>V\>p?�4�M�{�T>۟&>�z=�B?�m6?�A���=��fH>���=��>D�?�4??0�>�X�=�~ӽoO���̿��,�M�K�>�_�*���=i��P�6�h����6��@�=�?�>e��>�X�>���>���>�k'>qW�>��M>�G�=���<�x���^E>n�=*�ޤ��_���8��=����cq�}a��F���V��\�����=���=�?j\?�T)�"��E�f�4������h��>9��>���>K}�>7�=1U��U���A�7PH���>.gh?���>q�8���=��,�$��:���>�>��>�c�����F��2Ц<���>͝?a��>E��3G[��So���
�aϤ>���=�f�=��?P�d?	�����/�};~V�!�7�*��^Y�i��j޲�`Y �"�5�8(��>N��|b�qȨ=���>�5�?�Rx��t=�Pp�2��^����%���$>p�1>��>��q>��Ծ������#�E�����$��c8=��>��>O8??��9?φp?>�?Ź�>�ϡ��&?�l�>!�!?a4?�I?�K?�� ?G��>�"?^�=� 1��Eg�M�p�_�F��s�=j�=4�=_��=�vD>8��=xc�<2W�<lgK=qb�<H�G%8��,��e!>1{>iw^>�a?e�$?�2���� ����p���<���=�G>����FwT�!|�<�O[>�1?��2?��>G�=��ܾ��jq����==�?h�.?zy�>���;�=���*�h����=M�Z>	�9�"=��^��ʩ�P6߽0Q�>��>X��=��>�/�?��I?_?ț��˺!�;s`���d�y/���y=X�>��>�!�R�˾��'�`�P�WJ>�2d�?7t����ú�=�/>�缚B�[�=j��=5�=�f�;���ZZ�=�+>�C�>ƃ�>��?�x>U��:򆉾B���I?�C��"%�����_�ʾaf��.>&g=>���gW�>�����������7�;���>�d�?�0�?Hc?sl<�a��o|>��J>�<>���<�*I�KcP�˖��a�+> Ӷ=���z����2��ZW>ȱf>P�׽��о�6���S����W5�����'?��|J�������K����׾� 꾱=��x���x�����O�������	����v?��c?f7B>���;w=J�Ot��Z����4M��㉾f���o.����̻��Ӻ����D@���x�KW+���>+D�=���|;���|f��N>����4? ��=�j���9+����>e�� �(��d���V�����̋y?֐6?�Dپ��)�����Ib>&?`��=�I�>'�R�ܒ@��q>ld?nf*?=�:�=����l��$��]�?`��?X?h���H�7�i��=��y�?���>�$?1m�h��2ӽs�?�6?�*>�FW�t雿�Y0�I��>t�t?�S����=�?4 ?2�=�G��e�>OH��n���6>��>��p�/$Ӿ��T>}��=���>t��>��o��M��>B�\&�J���>�����G�=~��>M��iog>�̈>(��<����#���`��*�f��/?KQ�?��_?�3?ʩ3�jr��1IV=,V��r	3>�ׄ>3�B���X���>�	I>���m�V��T��@C?
�?Ϲ�?\KE?��V�oJ������D �����N�b�T��RD>ɼ[=<��>[s%>S��v =��5>��>t[�>]��>�G>fC>�L�=�������}l���:��3;�������Խ��e2��EiA�0�&2~��ʽq�����#���=�l�@�F�������=J?ĵ�>���>��>��K>��g�gL�X�/���e�/�&I���ݾM'�r����L�K�8����+��������?fj=��<Oݾ>f�
>��h=6;�>c��=�>�p�=U�b>���>�5>�0>ʧR>�:�>��=Ĭ{>BT�=�'��A��t:�^�Q�%1�;l�C?<�]�g^����3�Fd߾�������>��?��S>��'����a�x����>XG�3�b�t�˽M��iO�>���>��="z˻74���w��6�Q:�=Ⰵ>�!>��m�����f>����=� ?wY��h �&��>�TV?�Pi?Ϥq?/i�>҉�>�T׽�Z=?�؀�j޺=ߑ?+&�>ӗ2?l�w?	�x?->=�>��	���ͽ,HV�q��J���&���xD=�}�<(���4l����X+0<��=�>�՚=�&��`�>�����g�>��"?xl�>�Q?֗9��I��%� Bv��m>���=���>\��>�1?�?��>�A�>T�3=�ɾ� ����>�,>�V>�mL��5>��>H3�>Y�c?�?�� ��gڽg�½�% >��>s�?��?@]!?��m>�kK�^:
�3dȿߏX���7���Ě�@�=�2w>��0=�,�c\v�1���U��7x�=�b�>�E�>yy7>ȠD���!=^f�>N>d>�n>���=��< �k�뤫;T��:f%+�t�=,ޔ=�l���5[��|
�a�׽�4Ž��=�.=����=��?4k?��*�0吽�?d��H�������>���>Z��>}a�>���=���pU�n�A�z�J�� �>ߥg?C��>Y�8��J�=��-���:Œ�>�;�>��>a?\��X�����Ĳ�<m��><�?���>����~[�@�n��s	��2�>Ij ����=��?~A?!�=
��H�Op��u��Ǫ�R���Ư�j�<V:�75��h��������},�ſ?
 �?ZQ�h`��w�Ƃ]��B��W ��[�s2�>��=@~R>֏��B?��WeO�
��􏩾��*�`�p>@�8>�S>]�?T�2?��]?�08?�:�>r`Q�F?}�Z>"�?��?�[�>��?i�?�e�>*'�>%e�=BY2��Қ��5A��\��m���q�<!�>qg>���pc�=w'>Rj�> g�=�5���H��W�=��>��'=���=�{*>\?��?N��=� > 8�<V2R�6���~�=�KZ>��C�:"�=Um�>1�"?P�?N��>}�=��)��Ҿ�r��z_�>k�5?��?b6@>�Ϳ<�Dƾ����9��Iq>
	�=y���.�W�ɾ�8ֽ���>��>�y[>H&�>x#{?`�7?�>h���F<�
nq��B������=1J=�B>��=7�ʾ��ʺK��@���?�Nͪ���~�����>h�>.�>��>�C#>���>xDʼ-1�=�|���=�~��?�h,?�8�>���>-/=+0Z�<5�>M?����J�����7���˼s�>>0\>GA���y�>Gԯ��r��v��/���>���?oj�?��g?�J�A���5X>$!d>�>j�<F%6�Ɯb�T{��4�A>���=��r��?��z�3<U�x>Ȕ>'̴��7̾���A��8��W8���-<l��R`�i5�k��t�8�|���i/�����MɾP��&�3���l��ē�7¾L���DŌ?^��?�s�>��<	�=���6�������T���v�*�
���l&=�~ݾ/#վ�<��< ��&K�w]b�]�	�I�>ef�=+E��s����IO����<IQ�(!�>�v�3ܽ+<<��ks>o����ꮾ��I������8���O2��2g?��C?�p�@~E�;+��б>��'?�� >"<?g�#d���>ą@?\/K?)��o�Z����%:Ὃ�?�[�?P*4?+Μ<�TY�w7g��^���>��v=��	?��ľ�^������Q=A?5�?|���>������M��Z�>��?�:9��:>4�?��>+ߥ��@���-��E�Bf�=J�^>�a���9������A]��(3>��>^j�>�=��_���>B�\&�J���>�����G�=~��>M��iog>�̈>(��<����#���`��*�f��/?KQ�?��_?�3?ʩ3�jr��1IV=,V��r	3>�ׄ>3�B���X���>�	I>���m�V��T��@C?
�?Ϲ�?\KE?��V�oJ������D �����N�b�T��RD>ɼ[=<��>[s%>S��v =��5>��>t[�>]��>�G>fC>�L�=�������}l���:��3;�������Խ��e2��EiA�0�&2~��ʽq�����#���=�l�@�F�������=J?ĵ�>���>��>��K>��g�gL�X�/���e�/�&I���ݾM'�r����L�K�8����+��������?fj=��<Oݾ>f�
>��h=6;�>c��=�>�p�=U�b>���>�5>�0>ʧR>�:�>��=Ĭ{>BT�=�'��A��t:�^�Q�%1�;l�C?<�]�g^����3�Fd߾�������>��?��S>��'����a�x����>XG�3�b�t�˽M��iO�>���>��="z˻74���w��6�Q:�=Ⰵ>�!>��m�����f>����=� ?wY��h �&��>�TV?�Pi?Ϥq?/i�>҉�>�T׽�Z=?�؀�j޺=ߑ?+&�>ӗ2?l�w?	�x?->=�>��	���ͽ,HV�q��J���&���xD=�}�<(���4l����X+0<��=�>�՚=�&��`�>�����g�>��"?xl�>�Q?֗9��I��%� Bv��m>���=���>\��>�1?�?��>�A�>T�3=�ɾ� ����>�,>�V>�mL��5>��>H3�>Y�c?�?�� ��gڽg�½�% >��>s�?��?@]!?��m>�kK�^:
�3dȿߏX���7���Ě�@�=�2w>��0=�,�c\v�1���U��7x�=�b�>�E�>yy7>ȠD���!=^f�>N>d>�n>���=��< �k�뤫;T��:f%+�t�=,ޔ=�l���5[��|
�a�׽�4Ž��=�.=����=��?4k?��*�0吽�?d��H�������>���>Z��>}a�>���=���pU�n�A�z�J�� �>ߥg?C��>Y�8��J�=��-���:Œ�>�;�>��>a?\��X�����Ĳ�<m��><�?���>����~[�@�n��s	��2�>Ij ����=��?~A?!�=
��H�Op��u��Ǫ�R���Ư�j�<V:�75��h��������},�ſ?
 �?ZQ�h`��w�Ƃ]��B��W ��[�s2�>��=@~R>֏��B?��WeO�
��􏩾��*�`�p>@�8>�S>]�?T�2?��]?�08?�:�>r`Q�F?}�Z>"�?��?�[�>��?i�?�e�>*'�>%e�=BY2��Қ��5A��\��m���q�<!�>qg>���pc�=w'>Rj�> g�=�5���H��W�=��>��'=���=�{*>\?��?N��=� > 8�<V2R�6���~�=�KZ>��C�:"�=Um�>1�"?P�?N��>}�=��)��Ҿ�r��z_�>k�5?��?b6@>�Ϳ<�Dƾ����9��Iq>
	�=y���.�W�ɾ�8ֽ���>��>�y[>H&�>x#{?`�7?�>h���F<�
nq��B������=1J=�B>��=7�ʾ��ʺK��@���?�Nͪ���~�����>h�>.�>��>�C#>���>xDʼ-1�=�|���=�~��?�h,?�8�>���>-/=+0Z�<5�>M?����J�����7���˼s�>>0\>GA���y�>Gԯ��r��v��/���>���?oj�?��g?�J�A���5X>$!d>�>j�<F%6�Ɯb�T{��4�A>���=��r��?��z�3<U�x>Ȕ>'̴��7̾���A��8��W8���-<l��R`�i5�k��t�8�|���i/�����MɾP��&�3���l��ē�7¾L���DŌ?^��?�s�>��<	�=���6�������T���v�*�
���l&=�~ݾ/#վ�<��< ��&K�w]b�]�	�I�>ef�=+E��s����IO����<IQ�(!�>�v�3ܽ+<<��ks>o����ꮾ��I������8���O2��2g?��C?�p�@~E�;+��б>��'?�� >"<?g�#d���>ą@?\/K?)��o�Z����%:Ὃ�?�[�?P*4?+Μ<�TY�w7g��^���>��v=��	?��ľ�^������Q=A?5�?|���>������M��Z�>��?�:9��:>4�?��>+ߥ��@���-��E�Bf�=J�^>�a���9������A]��(3>��>^j�>�=��_�����>�ܾ8$�����n �� ��,�8=���>��$���g>�e>�,%=Ә+�Zˆ�y���=��}L? ��?��L?9�>?�7�����g�T�.=��u>P�q>Ju->�`ٽn>w��>����p���3?��?�e�?�ma?�'��Svɿ��������!v�^�0>�F�=��_>�J�$��3Z>`�T�`��b>��>k7>���=�?>�=t0�=P���'����C�x���.����i�ﾜí��4,�+ݒ���$����{������8Y���׽�F��#�'��5˽�`���@�=O�?�?��><ȼ��.>�Ҭ�V�8��/�����$%�n����P���!پQ;[!پҐҽ��;�u���?� R�R�>���>���=H��< ,>��>�B>��4>8�>�xO>F� >��F>c�>�3�>>́>}�?Y���s��<���վ��<�8�>z#�?���}T=^8���6�elt�]�?�R<?/>�3�.�S�:�6��F�>jޅ��/�����T->J�>��>��<��>tz�>yƼ2垾���>��>�1>	���E��X����=��>��B��v�=$j?��|?=f^?l�>��>$��>5��>Ь����>i��>[��>��?@s
?w�+?:��>/�=v�߽w->N�u=B7L��BP�#6��3i(����S�C,��*����A*>��=��<=7:=IVڽ7��Z�<� ?��;?�'�>1�>o�)�9��EZ���߽Sp�=Ɂ�� ?��>Ac�>9�>)�\>!�@>+N	>\+ӾMe@����>�5>����ɩ}���K� ��>ꏬ>ZrR?�&e?E����T���*j>W�w>��?�-?��1?w�?�`>>lڽ	��ٿ5h��t���m<��#=�zw<�.�a�� -���w�3�/��j7=��=i��=�|�=�~>�	����N<� �>ge>]j>W����n��њ_<<=�� U>ں
>И?<eT�= hT>L�f���Q�Գ=�l=u����K�*�;;�/	?�?�+ʼ������U������-�7>�v�>Z�ν1??�(�>��/��1�g{��m �ep??	��?��<?����>�yp=�ͼ/�c>���='�=��=��h=�T��b.�>��?�>��=_�h�����o|u���RG,>��ͽv��*��?�=�?\����4��{�x���c�B/�>Z�ƾԘ���̾��)�;�a�#����.�����2�=��>:/s?�:����G>�񡾌�S�q��3����J+�<�$=+�>��Q<f�������E��$���0
�<���>���>eh���5?-�+?F<�>��?�D'?��[>,H��{�%?�[E��?Fg)?��5?�n"��v�>��^>�B�����>�z��:����|���z;�W���ɉ=�^M>���=�2�{�<��M>&׼��9�2<$��;=�A�9�ԝ� ���o��=���=��?�,?I��O���>-ͽ��6�x[���v>�b�>�>�߁����K>��>�m�>?"��>�P>��z�Y�)�q�3U�>��?Kl?���>����a=&������S1���
>��=�p��Kܾ��l��;m=TyQ>�}t>���>\�>7[y?ٯO?
=?Yu=��WR��ce�Q���1 >�����>���>��3��0�7eC�9��V1_����d�!��%����=9�%>{�'>5�R>$��=ҝ��2=Bݓ�+�h�$< ;���3�>�ِ>�H?��>�HԻ����D�E�N?Ы������~��[�����VG>�2>.x��˳>�P���`k�b'�����K3�>��?�O�?�SM?�P'>� ��9A�>J��i2�T�=-�=�xd�*�=�>N�:}���=��{�Bn*�('�h�<�_{�bև���<>���.�B���*�UX�����#�	�O��<������kp����Ⱦ֦M�?/.���r.�"/A�����*��Z�����?� �?,K�=Sw�>��:���M�"(Ѿ?��%#��Y��0�-���?�8������gt��7��7y�.����>��Z��0���}�j%(�_����?>Ǐ/?��ž�����@�VgX=�x">�7�<��s#���l����vV?ƒ9?*��p1��G�޽�2>�?1�>�w$>h���6�0��>��3?�-?5�Ѽ�O���ҋ�� ���̻?�r�?�ZL?j4��k�L�e��8(�K��>N�/?4?�B��}�a��
���ҋ>��M?tw?��M��:����>��9?��C��J�>��>�w>��T�8Sܾ�h'�HGS�n���-">#픽�~������V/�j7�=�x�>���>��-�dh�Mg>Y��ǣ��U<�p8�;f̾�B>b�?(��C�>e\;>C�B�& ��&|�$A���*��?4ح?o�8?�!w??_9��EY��������ٵ�>�?���O�.<��>�v�>e���"8�@��ԕ? k�?��?˦|?�1~�z�ҿ�A��P諭W��]S�=B}�=��V>S�ս��=��z=��<��=;�->��>��N>%�_>=e)>
.F>�M>�)����)��ˠ��f����A����g��	�w��O
�R�/������|l;�Ƚ�����˽�l��\6���X�����=�T)?&�>!�g>7U�:?=>�Î���%G����:�g����$�龧�˾S	t�t�kS�<���ѓ��hO�>�d��}��=�8�>��=Ք>	��=hn�/$>|�[=��>� 4>x﬽
'��>jl=�F�>��N>��>���)$j�����C�*�!3s�=Ά=�b?DtK���\�$�6��E�������>�?��s>����s����w��щ>Ɓ�<�����������:>\¨>Ǳ��7�9�|3i�Xj�������>��O>�n�=�ѽ''��F�7���=s��>�XѾz�=a�h>f�'?��y?�;?�p$=��>�^>�.�>���=�}^>�B_>C4>
�
?��2?7u2?��>ns�=Ō{����<ׄ�<i�P��Wü]q����V�5��J�;�3H�=/0=��ݨ@=b�f=�V��Ws�;V��<av�>�yI?Қm>�.�>�{Q�����w�y�s�V�KTy>~H����
?1�?v~�>b �>%C6>�N�=�,���׾���!�>���>+5^� p��2Z>��>��=u�(?��I?(����ӊ���>Q�>sX�>n��>!1?��>&3>�;;���lEп�%�	�+�����C���:;B��J��������ϽA ʽ̯a=]�>?�h>��Y>J�>~)N>�VG>%��>t�N><}=f`=�-��_8��L�Ϫ=GZ+�Tf��%���w<d�M=�C��n����%��b9��u��?�2?x�5=�>��S�5�Ⱦ4���=�>� v>D0�>�>~B=� �=�P�y�!���7���?�AP?4�>Joo��S�=�d�<�Z�=I��>�|>wU�>⋄������J��q+����>�_?/��> ���M�^�ANn��>��^�>2=ſ<<��?�(d?�I �xd�	/��/M������0�-������7����:ݾ�� ����հ����_>ƌ�>P}�?#��o��>�0��-��q�����,�=Ό�:
"?zh�>ľ��u��;������v�=_X�>��<��>���>���>�z?=);?��?C���w~7?<Q=>(?h�?�vA?Mu�>�l�>~a�c��<�Vq>��=����!;�5輐�н����Pxs>(�b>j��=��<~],�j��Vb���a�p�1�"��=�)�=Q�-<�s=㼯=(v�>a��>�������=��=(Խ+��O��V?>��z��.��x�=����Ԅ?�m)?���>�>�!h��,ھYk����>��"?�� ?���>�\(=�n�=Ο���;��+�=L٭=��= �����)��ؖ�F�~���>S߉>�W>(XF>&0�?��"?�D?��=����+w�m�'�B>=0m����>�6�>S�>�{���4�k�o�Sg��=�[�_=v�Z����=_"�=J>mku>2:r=���=�;=СB<x�W�n1�=	�=��>�>��>U9>8�8��)���5���?Q�>�k�y�����H̾���>���>L�>��Y��V?Q0�=q	��a\����ؾk�7?���?.p�?߯d?�3��ν��>o�{>x�.>���<�7���3_��ޞ<9>>����Cw��>)E�f�����$?��>q9�F�4�.�2֨���ÿ��+��V<�����$��9^)�d����~�O/��m3=pȾV[�bc���o��ېK�'�{��$Ծ��li?���{?^�`?��>ze'>h�
��2��Ι�bZ>ˆ���S�=4޾zd���>��G빾� ;T����	�ĶF�i������>��Z�9���?Lz���'�_���B>�G/?��ʾ�*��fR��Y=B�$>E�Y<m����%���b��!Z?��9?�����{��K>��	?e�>:0%>���~��ϐ>J�1?�&+?'��D���7��)�ͧ�?7��?B�;?�uj�7�M��v�筙��
?7W�>3�>�����׾ؖ���(?u�@?�E�>���%����I�͸�>�3?�~h�z�W>�W�>�E{>\����ݳ�6������=��y>&�����N�<�d�>z6�>(ͅ>���я�����>�3�Rb5�+�D���4��n<�@�>���>� 9�w�>[��>q�(��]8�q���������:}Y?b�?<A3?�Fd?FcξE�O�_���.Cf�&\�<�}?쉯>5>�� ?��><B����u���۾7�e?V @�1�?��F?�4�~�׿t������w޾	.>�V�= w >�f{�>3�<X�=!��;cR�=�xL>��>o7<>�Z)>#=5>jD>f�'>�����,�(6���%����:����*���y�����#�_�w���]l�����4Ţ���y�h������9^�;]�w�de�=���>�l ?7q->��>��h>r#��1�0��혾r����S��cϾ�,4�m5� ݾ�v�s�ξ�־�B>���ۓ>o%���J=
K?�[h<9�W=�B>E��}h'>g�8>A_�ݴy=��Ͻ��;�B(>Q/�>���>�>n?	>T䁿�1����J��R���
���R?�=����-����󑎾N��>�&�>e�0>�}4�E0��*XN�Tۚ>Ԙ�<����b5�!9�=N�>�a>|!3�b\�=� =l�׾)*����=�>�;>.W�=���ƼT�n@����>�0���t\>��>��(?��?��)?D	�����>7��>@��>�X9>���>b�P>�Ǉ>��>x�?��2?%�>��=B9нv�=��<����2�fH��6������=�Ԋ=}�~>���>m�<�;<���<�6<
��<��=�r?E\7?�q>�w�>�;�D��>V��.��M�>�6H���?ٱ?S_�>�:�>s8�=�D����m�}��셽�f�>��'>l"w�]��d׈����>�I��bd?�Fd?�����G�����=@>�U�>,�)?M\Q?�zl>��([�����n� {�f�k=G#=Jp�!y���;཈\�=�!��lӤ���=>�Q�>��e>�w>\�'> �x>�}>
d�>Yc�>^�=���<�Z�A��K ��0=c���*\��E������ c콷V���ͤ��u��Ę�/������S�?W�?\����>������3������=f->�:�=&ˈ>��=�7�Ԇ[�qsP������g?xHM?�:?ow��؁=z�����>-��>E?>m�~>�~<>�!{�L�����>��>"�U?�/�>�R�.o��ڈ��r���m=���=��Ҽ��?��h?�� �)���[���64������_�-ã���l���Ѿl>"�K!+�_���	aо\B���>&��>`��?,��*��<���r����iB�$o>%>���>XM�>_8��9h�K����ɔ�*�N=N�U=��>.z�=�i?ӜL?�Ϸ>���?&�#?yڨ>�'���(K?���>ۍ0?�tB?�W?z"�>a?��^={9��ZU�>X<�=@Ž'��8rD=5�.<z>�< 9>H�>5�����0����=�M���޽�M��of���mh;Bӈ<}YK=�1>!\�=��?�"?�S��C>��8-���k��\�����>W��>4������M��=7�>�r�>�.�>[*�>��/=w�� <���=
�j*>5�7??�>?�?�z����>�N߾���z�=�jB>E���sl��G��%�m��V,�URT>��>�G
>ic>�_�?��9?Q�,?��K�(�(�r�֍�U�c=�<���9�>�o�>���=���[Y'�[�h���\���(�A��a�Q�d=�G->�>�}�>���=N�>!'#=+��������<:K�<݆�>�6�>�U?��L>�{�Z<��$��Pe?v�߾|�y��A��)�͒�Ҵ�>�x?+Ʊ���?��^�(����0��!\+��CX?���?=�?�;?�p��-
�s>�Ģ>$��=�Y>lʽ�P���?>�ǈ>��!�O�-�Ν���Ƒ<Ӧ�>H0�=Ls8���ʽǶ�0A<����j�9�H>����ى��.�ߩ�����sO;�����	1w���Q<]8{�Pk�`Į��2���n쾍>L���~?�Q�?�u�>ĥ�>�-��{#�ܘ��XN=;˾X��	0��E����'���о����u¾{%��	8��Q��z�>�eS�®��3&f� �&��A;X�_>J�?�پ]l��a�,�ﲱ��2!>��L�#.��݊�io���Y�I�7?ҷ??����
����� >�!?�	�>+>\����,��x|>݄6?n�?����5��#�����H=;�?Z#�?%f@?-H���B���	���Y�?�?fd�>�+��eiϾP5��M?9?�&�>]�أ��S��ad�>�Z?^�N�Y�e>���>��>"�z��]�6�qГ�!�;��/=>�b�N���d�>>�v��=���>ʺ~>7X��n��b�>�}�k�߾,�H�LCA������I>��8?X�1���=9r�>IVK��F�v���!g����.���T?���?��?�x�?�1޾Gp@�,M��%wϽ5G�>2?"ON=5w>"*+?��>�h����*����kn?��?���?64?FE�Rܿ|Z���֫�����:F�=7�;=��(>.!?�ڞ<_��<�����<Po!>vl�>v0R>suW>��@>�y>��M>ك�� ������ ����E���v	�k~o�������/����� ୾@Kɽ�&�g[o���4��� ��*I��� ��5���
8?��%?Bd;�����Ds;�3x���2�F��	�P?�x����zB�z1̾���m�&�}q$�L'�=Ũ��B�>�ȷ�2g�y�>
J>��>	�H>���1��<�=�{'>u��=�|\�^I�=B��v�/>(�S>���>�=L�c��=�}����3d&�A��>(9w?�t.�4�Խg=�1� �4��?Q�+?~E�>ܝ��ה��Y-�m6�=U����==�Ag���ݽЌ�;���>�R�>Ė���oe���q^���>�?j>���<<?�N����O��X^���>�F��g=O7t=W7c?Y{?�?�����>#�g>��A>�m|>�?�\>�!Y>���>�f?wu(?N��>�V">�P��k��=�͗��M��>q\>��`ٽ�B��|�=�շ=�4�.y������(�=�˛=lQ=��9p�=+R?�>?j-t>H�>��Z�Y$���KA��Kֻ*7�>�Y��u�>�?o?i��>j">0��=ri��д	�ၘ��?u�>��l�E/�����[Ġ>��=�+?5�y?8�>��|��S�="�>Y�?���>>�/?[",?�(�=7���(��0����þ�0#� �ٽ�[_��	{�z۾����7K.�	����N�(�!=�k=�]>�z_>�O>��>WZT>���>>�x;>���=�u�=O�1��g��"z�<�k�[K=Pɽ]�Q��5�f����G�=��=��<�<��׽B��>��,?U9�G�x�s4-��c��$��G>�=�>O�s<y��>ٴu>q���I��y��HѽZ�M?�q?�;�>�ղ����=Y�<t��>gRQ>�%�=V�@>z-�=<4���T����>R��>E\?dj�p䦽%����Cw��+���@>s�t�Cy����?v9[?Sh��%ľ���	*�����<��lv ��ܜ�x���ȁ0���E�ք�I],��p������9��>���?�w�����mzо�h���7^���6��'s�	�Z�?8�>�>}>bV�d����j�%Q��v�����=҉�>R�=�X?�	?$9D?�eg?Z�>���>(��NK?�˟>r�<?�uJ?mvN?�<�>Wb?��}�)e��MM�>�qN�k�:��iƾb{N���<��t�l-�=K�w>�ɨ�DD���a,�@�i<����U=E�=��l���\<�?;�� >�A>��?�� ?L����v�����<�?��z==�o>���>db��J� �!>��Y����>�
?=d	?ݺ�>)����"{>���^�>'�>-,?`�?r�<��W���=�(�����칀=��J>�r�����u�����|]D>��>��U=.,>nY�?tl0?6<?~շ=(�	���k�q���:=�/w>W��>��H����|�E�ꃿ� ^�ӽ��CFH��8����S=B݀>~�=N�Q>�����wG>_�>վ�=���1ӽۼڽ�ß>Z��>T�?��>t骾�M۾���3"k?��b��������
�>o0�><T�>X�μ�
'?�B�=����Y���}}�<ި1?��?N��?t��>Ӿ=4ߴ�>Fj>~�w��Vd>�K�>�;������W`V�Nf�>*=��H��.�ʽ�!��k�>a�>F~���]Q�)�ؾ����`�ſ�B4�Gq�>�3��2��Or/�,���*����� ��=>�u����w�7�����g�F�96��Ac����+�T0�?�6?5�f>MY>�5����7M�:'Y>�A��i[�=<K�+3��5�-�!���]l���s!���B�nu+�cF>^���jd��7_�N�<�k	ֽ�]N>J�(?M4��̴��	����X�/>�1�Q���~��~���V:��v2?�;?�����������>�?#��>'A�>�־�4A��%�>eL$?j�(?F���҉��\����=���?x�?��@?�Uk�vj<������j�?w	?2��>�zc�Ҵ����:	?B?]��>s����6���4�p�>�KU?�\C��	F>���>�]�> ���]��*z�܂��7>���/>�.=�2�T�����A��=���>i=u>�$O�2���b�>�}�k�߾,�H�LCA������I>��8?X�1���=9r�>IVK��F�v���!g����.���T?���?��?�x�?�1޾Gp@�,M��%wϽ5G�>2?"ON=5w>"*+?��>�h����*����kn?��?���?64?FE�Rܿ|Z���֫�����:F�=7�;=��(>.!?�ڞ<_��<�����<Po!>vl�>v0R>suW>��@>�y>��M>ك�� ������ ����E���v	�k~o�������/����� ୾@Kɽ�&�g[o���4��� ��*I��� ��5���
8?��%?Bd;�����Ds;�3x���2�F��	�P?�x����zB�z1̾���m�&�}q$�L'�=Ũ��B�>�ȷ�2g�y�>
J>��>	�H>���1��<�=�{'>u��=�|\�^I�=B��v�/>(�S>���>�=L�c��=�}����3d&�A��>(9w?�t.�4�Խg=�1� �4��?Q�+?~E�>ܝ��ה��Y-�m6�=U����==�Ag���ݽЌ�;���>�R�>Ė���oe���q^���>�?j>���<<?�N����O��X^���>�F��g=O7t=W7c?Y{?�?�����>#�g>��A>�m|>�?�\>�!Y>���>�f?wu(?N��>�V">�P��k��=�͗��M��>q\>��`ٽ�B��|�=�շ=�4�.y������(�=�˛=lQ=��9p�=+R?�>?j-t>H�>��Z�Y$���KA��Kֻ*7�>�Y��u�>�?o?i��>j">0��=ri��д	�ၘ��?u�>��l�E/�����[Ġ>��=�+?5�y?8�>��|��S�="�>Y�?���>>�/?[",?�(�=7���(��0����þ�0#� �ٽ�[_��	{�z۾����7K.�	����N�(�!=�k=�]>�z_>�O>��>WZT>���>>�x;>���=�u�=O�1��g��"z�<�k�[K=Pɽ]�Q��5�f����G�=��=��<�<��׽B��>��,?U9�G�x�s4-��c��$��G>�=�>O�s<y��>ٴu>q���I��y��HѽZ�M?�q?�;�>�ղ����=Y�<t��>gRQ>�%�=V�@>z-�=<4���T����>R��>E\?dj�p䦽%����Cw��+���@>s�t�Cy����?v9[?Sh��%ľ���	*�����<��lv ��ܜ�x���ȁ0���E�ք�I],��p������9��>���?�w�����mzо�h���7^���6��'s�	�Z�?8�>�>}>bV�d����j�%Q��v�����=҉�>R�=�X?�	?$9D?�eg?Z�>���>(��NK?�˟>r�<?�uJ?mvN?�<�>Wb?��}�)e��MM�>�qN�k�:��iƾb{N���<��t�l-�=K�w>�ɨ�DD���a,�@�i<����U=E�=��l���\<�?;�� >�A>��?�� ?L����v�����<�?��z==�o>���>db��J� �!>��Y����>�
?=d	?ݺ�>)����"{>���^�>'�>-,?`�?r�<��W���=�(�����칀=��J>�r�����u�����|]D>��>��U=.,>nY�?tl0?6<?~շ=(�	���k�q���:=�/w>W��>��H����|�E�ꃿ� ^�ӽ��CFH��8����S=B݀>~�=N�Q>�����wG>_�>վ�=���1ӽۼڽ�ß>Z��>T�?��>t骾�M۾���3"k?��b��������
�>o0�><T�>X�μ�
'?�B�=����Y���}}�<ި1?��?N��?t��>Ӿ=4ߴ�>Fj>~�w��Vd>�K�>�;������W`V�Nf�>*=��H��.�ʽ�!��k�>a�>F~���]Q�)�ؾ����`�ſ�B4�Gq�>�3��2��Or/�,���*����� ��=>�u����w�7�����g�F�96��Ac����+�T0�?�6?5�f>MY>�5����7M�:'Y>�A��i[�=<K�+3��5�-�!���]l���s!���B�nu+�cF>^���jd��7_�N�<�k	ֽ�]N>J�(?M4��̴��	����X�/>�1�Q���~��~���V:��v2?�;?�����������>�?#��>'A�>�־�4A��%�>eL$?j�(?F���҉��\����=���?x�?��@?�Uk�vj<������j�?w	?2��>�zc�Ҵ����:	?B?]��>s����6���4�p�>�KU?�\C��	F>���>�]�> ���]��*z�܂��7>���/>�.=�2�T�����A��=���>i=u>�$O�2���
`  �   =2y>����p�;����F��յ���'���/?,�ʾ����jI>M>p �T�o���|��V��.�L?��?;�?sGU?`������+�s<���>9�e>p��>d�E>�Qr���>�T�>0�3��t1�K��g�>\��?���?ug?d�]��|�B�x��e;��XX�=<��R[�<�q��=��=J�7>�
�;�6�Yi����I>��>ؼ2>���=b�">J@>0ֆ��C$�����$Ƀ��N����;�*��������D��x��T����8��&f��B�W������}��&
�� ����� ?�?��>Y�>�0d=v8 >sо�} ����=&�r����Xf	�1z�.����#�	�5�Z��_�ML���T�-��>�]#�@B��|��>���=l�`�>l�>ϭq>� >P�<ı>�{z>�vZ>�>�>�T��#>D�G=��x����1����̇��+W?p���o����<�c¾�⾾l�>fw?i�>x_�k�y��'*��?�����;��wM'�M��)�>���>���<Y����Z'����	���>y��>\?�>-V�<>��������=��?�z����=˲>�*�> ��?��?G��=�1�=`��>���>���>��?0AG����L?EsU?��=&=>��p=%��Q;>�G�=�P���d�=$@x==�ʽ�ګ=�G�#�o�v���Đ=8>$y�=e�i��pd��M>߯t=��?��>b��>��>S5��2
q��6��Z�~��М�w�?��>ܣ?y!?=C�>Ne��kL>�W\�0���\�>�D�=PS-�3ō��=�OI�>��>n�?<?�[�~þB��9Y='�>�D=>O�?��>_�0=e5�<����qǿ �%���'�D��c�,��������^|�=O�%>)BJ�Kh��0�����>)�>\�> 5*>o��=�O@>��>�ZU>�����Ъ�m߄=�I��R���\>�އ=C���"���=D�y��;�B�÷��f&�C��<i�e�?�/?aƘ;�R4��qA��Ծ�k���7�>���>m)�>�k�>���=�Q��ysU�T�H��NF��?��^?���>�@7�c�=�i�Ƕ�;���>�g�>��2>��#���+�J/��2xX����>]�?03�>��Z�S�l��5���>�Z�=^|T�<�?��[?_⾶�n�c���R�~V�L��;�/a<�c��Oˌ�Gg��&��?��UvӾ[䥾�$�=�>[�?��M�ҷ�<� о���������Ǧ�)�y=�o�<�7�>m2�=D���TL]����]f���A�ڌ?>��5>�:|�2?w�M?��>��P?��>ػ�>�3L��)�>��?׌_>$��=��D;��>��[>��>X��5�<'?ǽ�e�ao}��>��	=�v��ˠ�=�ҟ=������>I�=������$�B�=��<�����ئ<Y=tP�>�� ?��?;�0������-���?>mC��/ �>Ճ��4�׾�&��f�=��?��4?A��>`�
��E��)�=����g(�>�@�>I�?5I�>���Fdl�ct��@L���>ӝ�=��i����8߾����yнL�=��>�H�=��9>V��?.2E?��"?�=>�~�h��a�ivݽ����M�>	�e>�@��`羳\E���g��1P��w
��@��F�W����=���{>2�?>:>:0�=l���{A�ʸ���<�ˎ=]ܢ>�>�:�>�l>�£=T��"���G?U!�l-��WH�F�������/>��=��?�^�=��χ�^L��ݐ>R&�?�m�?`�?�������/��>2�f>۪D>�饽�V%��]a�b�	�^�O>AF>c_L�$9���?�(�>B�l>���N�ʾ)�ƾ͜�<G�Ϳ��7�ﴸ��K
�6Ii���!��?	����=.���0��\׾4YK��[۾�Em��U��nQ��۾�߹���/�b�? O�?�ڂ=�������=�����P2>����U���מ�/��mW��덬�X�Ѿ�n��2��_����x>�_������#���S��Bн�	>��/?�����[��
.�Xr�=��>}q9>⿇���g���'�"r??��S?��B��x!�F�=oYR=��E?���>�6��N������?�O?���?[��� ���l������=��?Y�Z?#�<?h�پ�Z �7�:��y��%?�=?D��>cZ>A�v6�rJ>�o	?��?�f$>A�p����Qa'?,?����>z�>v?��t>�뾾��	��=�9����y=��?>��>�B��a�J^�>ne�>T;F�ZXV��T�;�'>��վ�
����n���ܾ�j!�
�3�m{K?�Ͼ v2=h3�>�1>^�9��@���Kq�{�;��c?'��?`}/?��[?x�����`��		#�OE8>�R�>�<K�&�=>)ef>����v�6X�9$(?)�?��?��B?��M�Gӿ�
�����������=-$�=��>>��޽.ȭ=��K=࿘��c=���>o��>o>�:x>@�T>؛<>�.>M���d�#�yʤ�ْ��[B�� �פ�swg��{	�5y�����ȴ���ԗ��I���Г���G����V>�8ݾ�f�>^��>{�?*�?v'���)�<���Z������/ͼ�G#�c*���G���V��X����=�������q����A߾{�>"�=)m#���>[v�<��=?�>9������=1~k>�_<�(�=5�A>vdL>0>>n>jP=>'��>����Z�I�N���tC����=O~=%�9?� >{�'��5���� �]��;��D?O�$?7X�����N�Ҿ8��>g��~V��½Ӿ=v�t>�TT>7>7��=�|	�����ϟ����>�O�=¥>!7�< wʾ�{s����=���>��پN�<>S{Z>(�>Qy?�s;?��<���>4$>�QN>u=��[>R�>ԣ>Q��>��
?!#?���>Ņ�=9��}wH���=�-_�������U��`����D�p��=|`=]�]��+�=$����-�<�a�=sx(<6�����=a��>ٖ?�Χ>�ھ>�嗾��A�N0"�p������=[���e�>�f�>���>]�?Pj�>���>��5�>X������U?�2>o4&�/�~�%��zx>���>N�?�q(?�n,����H2=z��<�A�>�9?k#?lc��>�tW>�
�a��`>��Y����J�̽J��������b��=�=����ʽ�F��	�κ	Z">3{>[O>�@=��^=]U ?�jM>��{����M<]�s=��<x|�=\���k<=>�<�`=�
�<�"��5RG�(/'��k�F;]6<3a�>v1?B�ۼ��N����&b*���m�>�,}>pi?
E�>��\�� ��D��y"�z^q�� �>�jt?/!?N�ܾ�!�>r�=SP���}$?ș�=��!�8ؽM��k8��z>~m>A�	?�2�>���؀w��y,�ȼz���T>4��=FȽ�?�W?�������u�r�G�r��NHQ���0�l�'�%밾5���I��彾^��dP�,>xE�>�ʦ?�����
>2Yf�Z0����*��*���$� �?��;>i?	��w����?�ؾ��U��V�=7'�>z��.>? -?��(?�]?�X�>�0>����x�Q>
g�>�<"?���=U+�>�7�>���=CnͽW|>��2>q�=K��mO�rS9��������=��=�4K=aZ�S唽�xP>X����ku<�;�=;�i<�$�8{0�=���=���>a>Z�?+�h>��=���<A���8��>/z�>$�����2?�X	>�>��n�<>[���ĽP�B?�@?9Ѕ��V����=�+�I/�>��*>�)�>�x>�Y��d=^J��
�A��Z>>��F>�^������Vʾ�̾Y�ٽ�>{>ë=���=���?�Y?��>��>�<`���������pz���P>:�	?�Ԁ���"����;��f��L�5澊:��o��+_ٻ"�=��>�k;>7�	�!�%�#6>;b�=���������;��[>���>���>�m>�����
Ҿ4	,�,[E?@���6J��8��߯�A��<B�>+�K>���9D?4L.�� y��'���g?����>r2�?���?�0?`ý�!½;bX>:�>ќ�=�ō=hH�*��:�:�̣>�ւ=��I����z%<.>�с>CBv�8����� ��V�Կ�gG��޾�Ҿ�����r=���^>�bD=��5�L��9���s�S�F�+:A��� �ha���R��ᗙ�]�?*�C?/�����
����վ�a�U�?/� ��t��拎�	�k��&��`�o���Z����_����Ͼ�þbz�>�z��8'���`g�,;� R��{;�=��]?y��L��� (��/Q>zM7>�q�>�y��V�j��a��aB>�r'?�,\?�8u��z��U�J>�Z�=��#?�?b�=_�þ���N�=A�{?�F�?:�>����'l���p%��|�?enF?T'=?�NB�������ge��V�>Jx
?G>>���$	����kLg?'�?�(Q?�5ؾ�`���Q�1��>B�n�OF��C>���>�j>��Ja�=j�G>䕹��I�>��> �,��-��`���|픾g����z�>�}>>8Q����a���\<�Ҿ �c�u:��$Ww�_�ƾ%B����>�G�$��=2au>;��=�F:��5���Ճ�ò�1JX?Rդ?2,!?&D?xXվj�'񆾮[�=Nl�>���>R�>��=u��>��>ߧ��<�P�t꨾�?a�?F��?"a0?U�o�%ƿ��q��Zݾ1곾R>�*;ڇ�=�(�X��<��=�dC=�}0=�~�<>;�=��w=��?>�n>�*B��t>�����Z���Ŀu-��6��r$?�$��4����+�K@���r��������E;�#ݏ���Z�~Ɛ�sB�B O>z0�����>sB�>���>De�>����Nj�>	���� �\Z�;2^����S��#��2�Ⱦ,%6��RN�+)��Mپ* #��V�Z��>4���ݽ��>,v�=?Gͽ�+�>�[���Z>č>�j->��}>�<%4~>���>���>//=��>/ļ�n�����>��1�`�eT��x�A?㕭=�g��x!��߾�۾>>�?G3?�5ξG���4�Z��E?����|��Q@�K�A��U�> M�>ib0=�A��D"���%Ǿ�JڽqNN>S�?-4�>��E�����NK�R�>C1?����b-?>Li��?g�?�P�Ԃ ?��?A����%>Y��<��>�	?I��>�> C�>��>�1+>�t_��Q��zq�=�|%=%t���� ��;@�=�����es>������=�����o}=w8>R�^=��T�/�&=\'�>�:?�I�>��?Nwƾ
8��(/��oȾ��>>�_��-�>�^'>4}�>�%.?Y	�>b�?�� ������2�?#m�=��cK�%;���?rM�>�p�?�D;?.��̠��zu�=�l�(,^>�2$?��??�.�,>�>`�����F��rQ��8�=F��<^J���K��-h�*%ܽ�VȽ�����)�L�זƺ��V=E��=��M=͟>�W�>�O�=U<>�=6�<�[3< g�K?Լ��=l3�<�)�����|����
��
�_U�}ߑ<rO�=���)ؽ>�g?Z�+>*:= OX>�q��VǾ��?��=��>��?B�쾾����g��N!��Rҽ��?]��?]J*?�bo��x>�+��l�=��>���>�у<|�3=C,�/�E�g0Y;q��>!�>V=:>��j�"�E�d�Q�y�վ�+>�M>�ǭ�Wv�?]�H?�����z�fs��GV3��	�~|�<�����0���|ž~��b��ʦ���b`���->�I�>�>�?�Z��\7K> �4��)��� ��1��0��5;�N�>?q/=�u���оSb���"V�؍>ı>�8=y~�>�D?D?Z?M?��!?f��>�zֽ�4�>Qg=0?;��>�+�>�x�>蕠>��5=�n>���;(��Mn������Q=���<�~>�/>��A=���P�=�S�=��=�y�SX���ʡ=�k)=��=��=�܇=5h>��?�@�>�+>�LN>�	�_1l<���>�->~b�>ld�=�(;��=�z��̟�>�$F?��?�g�$ˑ��-��d�>�3?�/�>�>kɯ��|�=��������?�j�<(T�=����H���CվW�|�2�>��h>j�=�y�=Fz�?��/?�:(?X̻=�!��p�}�����H���c=XR�>�S�<�������Z�'��!`��e��N�����x�:?���=��D>��>�e"=ԧ�=?��A!ͽ�̓�qr�R�h�i�>K�1>Y��>Wm->�q����
��W"�/>A?���|���;��4A����C�
�>AJ>o{ý0� ?��׽ͻ{�뢢��[:��$�>1��?į�?�d?��l` ��̓>�*>�-�=R�=��U��Ͻ�%߼���=l	e=
!F��w����q���Q>h�s>^ݺ��Ʈ�Zz��oj�<�Qѿ�-��1�_N�%�?���G�R���|����������)Ԝ��ha����q߾ ־�Ԙ�>���/��߼�Q?Z�&?�G>� Ƚ�ؾ�xž����8�2������^ ��V/�=�i��L����_�{�پ5���l���f�>�7��c���p(��2�b&=pO�=#�?�i��4�ʾ�j��Ri>pU�>t@�H�a��9�����fx.?��A?��?���d�e�&> ��=�8?`��>
�(=]-Ⱦb���>~�L?IƓ?�ee>;����my1��۬?�l�?�x??��6�$о�f���`/>��#?J1>�7�>�"�S�þ���="`?��?�38?���q��8�|>.��>�-p��G��m>N�g>���>h#���A���=���">R�>�$��Q��)��������=���>�$=�7X�4��=2y>����p�;����F��յ���'���/?,�ʾ����jI>M>p �T�o���|��V��.�L?��?;�?sGU?`������+�s<���>9�e>p��>d�E>�Qr���>�T�>0�3��t1�K��g�>\��?���?ug?d�]��|�B�x��e;��XX�=<��R[�<�q��=��=J�7>�
�;�6�Yi����I>��>ؼ2>���=b�">J@>0ֆ��C$�����$Ƀ��N����;�*��������D��x��T����8��&f��B�W������}��&
�� ����� ?�?��>Y�>�0d=v8 >sо�} ����=&�r����Xf	�1z�.����#�	�5�Z��_�ML���T�-��>�]#�@B��|��>���=l�`�>l�>ϭq>� >P�<ı>�{z>�vZ>�>�>�T��#>D�G=��x����1����̇��+W?p���o����<�c¾�⾾l�>fw?i�>x_�k�y��'*��?�����;��wM'�M��)�>���>���<Y����Z'����	���>y��>\?�>-V�<>��������=��?�z����=˲>�*�> ��?��?G��=�1�=`��>���>���>��?0AG����L?EsU?��=&=>��p=%��Q;>�G�=�P���d�=$@x==�ʽ�ګ=�G�#�o�v���Đ=8>$y�=e�i��pd��M>߯t=��?��>b��>��>S5��2
q��6��Z�~��М�w�?��>ܣ?y!?=C�>Ne��kL>�W\�0���\�>�D�=PS-�3ō��=�OI�>��>n�?<?�[�~þB��9Y='�>�D=>O�?��>_�0=e5�<����qǿ �%���'�D��c�,��������^|�=O�%>)BJ�Kh��0�����>)�>\�> 5*>o��=�O@>��>�ZU>�����Ъ�m߄=�I��R���\>�އ=C���"���=D�y��;�B�÷��f&�C��<i�e�?�/?aƘ;�R4��qA��Ծ�k���7�>���>m)�>�k�>���=�Q��ysU�T�H��NF��?��^?���>�@7�c�=�i�Ƕ�;���>�g�>��2>��#���+�J/��2xX����>]�?03�>��Z�S�l��5���>�Z�=^|T�<�?��[?_⾶�n�c���R�~V�L��;�/a<�c��Oˌ�Gg��&��?��UvӾ[䥾�$�=�>[�?��M�ҷ�<� о���������Ǧ�)�y=�o�<�7�>m2�=D���TL]����]f���A�ڌ?>��5>�:|�2?w�M?��>��P?��>ػ�>�3L��)�>��?׌_>$��=��D;��>��[>��>X��5�<'?ǽ�e�ao}��>��	=�v��ˠ�=�ҟ=������>I�=������$�B�=��<�����ئ<Y=tP�>�� ?��?;�0������-���?>mC��/ �>Ճ��4�׾�&��f�=��?��4?A��>`�
��E��)�=����g(�>�@�>I�?5I�>���Fdl�ct��@L���>ӝ�=��i����8߾����yнL�=��>�H�=��9>V��?.2E?��"?�=>�~�h��a�ivݽ����M�>	�e>�@��`羳\E���g��1P��w
��@��F�W����=���{>2�?>:>:0�=l���{A�ʸ���<�ˎ=]ܢ>�>�:�>�l>�£=T��"���G?U!�l-��WH�F�������/>��=��?�^�=��χ�^L��ݐ>R&�?�m�?`�?�������/��>2�f>۪D>�饽�V%��]a�b�	�^�O>AF>c_L�$9���?�(�>B�l>���N�ʾ)�ƾ͜�<G�Ϳ��7�ﴸ��K
�6Ii���!��?	����=.���0��\׾4YK��[۾�Em��U��nQ��۾�߹���/�b�? O�?�ڂ=�������=�����P2>����U���מ�/��mW��덬�X�Ѿ�n��2��_����x>�_������#���S��Bн�	>��/?�����[��
.�Xr�=��>}q9>⿇���g���'�"r??��S?��B��x!�F�=oYR=��E?���>�6��N������?�O?���?[��� ���l������=��?Y�Z?#�<?h�پ�Z �7�:��y��%?�=?D��>cZ>A�v6�rJ>�o	?��?�f$>A�p����Qa'?,?����>z�>v?��t>�뾾��	��=�9����y=��?>��>�B��a�J^�>ne�>T;F�ZXV��T�;=2y>����p�;����F��յ���'���/?,�ʾ����jI>M>p �T�o���|��V��.�L?��?;�?sGU?`������+�s<���>9�e>p��>d�E>�Qr���>�T�>0�3��t1�K��g�>\��?���?ug?d�]��|�B�x��e;��XX�=<��R[�<�q��=��=J�7>�
�;�6�Yi����I>��>ؼ2>���=b�">J@>0ֆ��C$�����$Ƀ��N����;�*��������D��x��T����8��&f��B�W������}��&
�� ����� ?�?��>Y�>�0d=v8 >sо�} ����=&�r����Xf	�1z�.����#�	�5�Z��_�ML���T�-��>�]#�@B��|��>���=l�`�>l�>ϭq>� >P�<ı>�{z>�vZ>�>�>�T��#>D�G=��x����1����̇��+W?p���o����<�c¾�⾾l�>fw?i�>x_�k�y��'*��?�����;��wM'�M��)�>���>���<Y����Z'����	���>y��>\?�>-V�<>��������=��?�z����=˲>�*�> ��?��?G��=�1�=`��>���>���>��?0AG����L?EsU?��=&=>��p=%��Q;>�G�=�P���d�=$@x==�ʽ�ګ=�G�#�o�v���Đ=8>$y�=e�i��pd��M>߯t=��?��>b��>��>S5��2
q��6��Z�~��М�w�?��>ܣ?y!?=C�>Ne��kL>�W\�0���\�>�D�=PS-�3ō��=�OI�>��>n�?<?�[�~þB��9Y='�>�D=>O�?��>_�0=e5�<����qǿ �%���'�D��c�,��������^|�=O�%>)BJ�Kh��0�����>)�>\�> 5*>o��=�O@>��>�ZU>�����Ъ�m߄=�I��R���\>�އ=C���"���=D�y��;�B�÷��f&�C��<i�e�?�/?aƘ;�R4��qA��Ծ�k���7�>���>m)�>�k�>���=�Q��ysU�T�H��NF��?��^?���>�@7�c�=�i�Ƕ�;���>�g�>��2>��#���+�J/��2xX����>]�?03�>��Z�S�l��5���>�Z�=^|T�<�?��[?_⾶�n�c���R�~V�L��;�/a<�c��Oˌ�Gg��&��?��UvӾ[䥾�$�=�>[�?��M�ҷ�<� о���������Ǧ�)�y=�o�<�7�>m2�=D���TL]����]f���A�ڌ?>��5>�:|�2?w�M?��>��P?��>ػ�>�3L��)�>��?׌_>$��=��D;��>��[>��>X��5�<'?ǽ�e�ao}��>��	=�v��ˠ�=�ҟ=������>I�=������$�B�=��<�����ئ<Y=tP�>�� ?��?;�0������-���?>mC��/ �>Ճ��4�׾�&��f�=��?��4?A��>`�
��E��)�=����g(�>�@�>I�?5I�>���Fdl�ct��@L���>ӝ�=��i����8߾����yнL�=��>�H�=��9>V��?.2E?��"?�=>�~�h��a�ivݽ����M�>	�e>�@��`羳\E���g��1P��w
��@��F�W����=���{>2�?>:>:0�=l���{A�ʸ���<�ˎ=]ܢ>�>�:�>�l>�£=T��"���G?U!�l-��WH�F�������/>��=��?�^�=��χ�^L��ݐ>R&�?�m�?`�?�������/��>2�f>۪D>�饽�V%��]a�b�	�^�O>AF>c_L�$9���?�(�>B�l>���N�ʾ)�ƾ͜�<G�Ϳ��7�ﴸ��K
�6Ii���!��?	����=.���0��\׾4YK��[۾�Em��U��nQ��۾�߹���/�b�? O�?�ڂ=�������=�����P2>����U���מ�/��mW��덬�X�Ѿ�n��2��_����x>�_������#���S��Bн�	>��/?�����[��
.�Xr�=��>}q9>⿇���g���'�"r??��S?��B��x!�F�=oYR=��E?���>�6��N������?�O?���?[��� ���l������=��?Y�Z?#�<?h�پ�Z �7�:��y��%?�=?D��>cZ>A�v6�rJ>�o	?��?�f$>A�p����Qa'?,?����>z�>v?��t>�뾾��	��=�9����y=��?>��>�B��a�J^�>ne�>T;F�ZXV��T�;Y�>�K�i�y�\���ɾ�����>��?���#,>+�O>)C�>�]��爿�8��yMX��4?_?�?Md?ȗ!?)�־�r��%m���eA>�S�>�`��ս8V�>J ?�e��gZ�N!�a=�>���?|��?�@?�c��8տ�Ԧ�8����І�-�>�n>;CC>`��J�=�����=g���e,>�:�>� r>�F�>r��>�h�>O�B>���}'�s������}6;���p���F��?"�ۨ߾
�S5������a�3�D
=Uݼ��=ߧ�g�-;y����F ><�>O�>(��>DAI>��%>�h�����i!��]t��d���k���ܾ#섾��8�Q�M���c��У�ڈ��:?#���Օ=�Q�>�f��z>}�>*c�=�Y>�JH>r��=�>'$>Y�=>B�>�4L>��=�>�3��ˆ�z
���db�M6�8z�<�9Q?�|�bV��t`\�8%����1�*��>ZX?/��=N�D�ӣ���㡿cx?��=5i��-���t�mA
?�	�>"tf>>�q���=����X�Z�4�>�������=��=�ؾ4����}>�R�>����Q=��>�o4?bVr?��8?��u=\�>K8
>*�>��7�l>if>�>?�?&�.? '?���>��=�cz�?��=�̮;�<��˼�{���ƻ[r ��ʼ�3A���=7�1=������L=�Ԍ<�� �=��<O��>/p@?��>�$?9����5��������>�ی>J�#?EX�>�39?�U+?�l�>n�j>k��>bV�)��:�>��S>�S��.Z���M��/J>ޠ>Z�R?+GD?���j*��}��]'=0V�>!�!?k�A?���>]Z>�������%ݿ�:�_����b�ʼe�ռ�٘��jM�A&���|-�*�@�G�
=���>�>��>^O�>�^F>�W	>7��>9"�>�Jt>�
��1콽�Z?�1�];Y>w��7Im>����O�=�G�r���{�����xe�,x ��E�&Z?r? �����)}�_*��\ɽ�-n>���>�e?���>�q>j���k#^�j�X�	����>4?g?�?�����QN>����yw>m�?M�>���ŗ���j#���l9����>!y?�6�>� s���S�@�x�!*�@t>�v�=��h��L�?�yL?�پ���� ��Y������I��Y���Y��ذ��O��;R��+�����J��B>o��>�h�?Q�<���=>�\������~���b���=8�<8�H>[��=�;��6�`�-��S��t�1w� D`>?,>�%�>�$?yX^?`l3?��?;D?��h��4Y?cI����?he����>�>?o?�?I�?K�н��Ҽ����_��zݠ=��%>I�_> @>�r>�2	���=#5�����<��ѻ�Nf�lW�<Ž����d�>��">�	�=�u	?H^6?��<�P�=�������a�=�L/=_��>����%Ѽ�]���>_��>�/>?E�!?��w>������^����Ew���?�x-?���>i�"=0>RL�n@�ՆN:�>����n�|���?��.<�3��>�ֆ>D�=��>؊?�Hh?���>ż>��ݾ�᡿ͯ{�g~�� �> 	<^�)>!������o��\���G�)<4�x)�<`�b󭽫��=a �>Yf��K�<�2=R�=�x���>�U�>W��>�e ?0+�>X%5?,�>��>�S�����;�I?ƌ��������äо����>��<>�D���?�����}��勵x]=��1�>�r�?e��?�Wd?�3C�L��~,]>�]V>�}>e�)<V?����톽�;4>��=�by���"�;��\>�y>i�ɽp�ʾą侅iH�}���.lX����=¾�ǜC� �3�$����>�J[��a�JSi<�}�n�=f�>�vʽ�4��ߦ�������?��k?��=�^N�x����F�Ӯ����=��>m��R ���0=��̾�|8��k��D��[��y	���+���>w5 �j#��[q������>�>�?da�ϧ���,��
�>flx���@=Ө����k�����=��Q?�6B?̾A(K��B1����>z:L?٩�>2X*>���q�����>��#?,U?^��=�Ț����"�=7��?� �?LS/?0�+�f�|������=�t?�h?!�>ǂþ(l�W�=%�>h�I?�~����5�V�{�����?7?�<s?L�P��e�=��?�Q�>�$����x�ϛ���Q ��89=A�>p)u�7ӕ�A�S�j���,�p��>�AM>;h����*C?*˾�[Z��Q��,���@U�="ͣ>��K?A�OY����@>��?����4��Q5��lĂ<��&?#�?ǘ�?7�0?���#]�h=��(=�>�S?K*�<ݩG��}f>v�7?{������h:��?�p�?<2 @��x?�FW�ŭ�����
��& �旬=��/>��A>�Z7�'>V��=�Q<���;�Ep>���>��l>���>:�A>�8�=Kt�>Fe��nL(�p���2J����D��p�y*"��!@��y��k���b����|@�����/w�F�缐��;�}��~F���=��'�|rN>�ɩ>|��>;|�>p��>�.>�]��]���"���A.9�D�������@�;gy������ �I��"��m�Ľ�!ľ��>{o�=餻=ϟ�>9D����=H�>�Y=	�C>˳;>+�z=,t>!Zp>־W>nh>��=�/v=3��=�4�tuQ�ߤr��\�������EI��D?��4�񐺾�l_���O��Ş���>Z?��.>��$�~��������x�>3=f=�1W��`i��W��"w>�P�>^#�>�J<9:k,���:��c=)�g>p�=�����Ĝ�Z���~T�=�f�>o��d�B���>I0?P>a?��2??��=Lh�>��h>x��>7=�/>>=�>�q >��>�1?9p(?ی�>��=5qb��	>F��=9�,�4���ky��}��B����=�p�FI=��B�����f=��;���"�rw�=1��>�;7?���>.?EA��o ��^�)���	}>_�$>P?�>��>� ?�6?�*?�x>�Hq=u�޾���7Z�>��>@2b�D�����ܠϼ�>�o?ǭb?�m���h��>���=f ?�)�>��P?폵>�D�>=�=m�����ؿ��T��-�w��H
�<l"=�-���я=.=�3 �Gc���8t=̛�>�>Z��>^�>��A=��<>p��>�`�>�S>�
 �l�=�1�%���K+�;��+�F 6=���ꀽ5C̽RM�1��	���6�B���l��_]�3f?��>�6G�x�^�[G�l�Ⱦ')ʽ���>��=k^B?J�?�i��߾��K���d����6]�>�Ku?�O?�[����a>9��>j>?W?V��>W��}�J��hz�����f�*��*>��?�U�>y���5�`�STR�N�.�-�1>5t�=�� =`�?�/F?׃��q*��5D��Z�M�)���,���:�ꇾ#��mu+��XM�{��b�	�M7R��@>���>m�?�<�XF�DQ������!��02žX�<>��:P�]>�E�=�V}�U�e�`�,�*�žU�ﳽ�>�ٹ=t	�>�L\?��`?Ud?�O&?*�$?*�����w?�j�>#?�>�X�=�}?14?�b?�z�>�� ?�8�/�=��:��)&>�=��	>�e+>t�f>xAڽ��>�iI>���==<�<�G��8�=�Iǽ�B=�vR=�e=�V�=��?%>B?l��;�u�8����pѪ���U��t�>B��>��S��9��B�(=���>�x?�oC?�g?H�d>�殾���� �ug=�w?}�J?P�?ۘ>��}>�O��<��.�]=�:>�%���=^�V��������g�4�q>��+>���=`�>�v�?��`?xM�>�s��;Wg���`��+u�k��=���=zI+��M��%����4�+��V��jF0�u;e<"��@�
�N{Z=W�>�<2��5>�@>�@&>Y����mC���v���޽y�? c>{�_?��H>�i}>Π��D��jd?����R#��n�辞����T�>�g�>0C��]��>R�y=ch/�ǫ����p�g�9>���?r��?�?y����s$�Y>=��>�m�>X�J�7�����%��ѵs>pe�>�z���H	�;�$�>�C=h������}��Bdý�ۤ�q�K����;�t=�_I��Ǿi_"=ǰ�%#J���-��z=GH���;|=�γ�2��������
���/��x�?T�q?y��=��k�rl�~b����Gdg>��u�ֲ��=ľ���� y��d���qPX��\׾�O0��M����ࢽ>�Yν�9{�%#���� �r2�}�>��X?��ݾ%��!�K��U�=�=��`����{5��$���/üX�*?�5^?aC��-C��dv�UA>��N?��>��>&��̽�y>1V?�P?����^���m�u�˶��H��?\��?w:?���T�M����kGa��?!W?׵�>h���Ҿ�"����>_5?h�>� �Hs��؁��>��E?�u�K�t>���>0q�>����G���~Ǽ39_���%<�=8��=e��,S�z /���=���>^#�>7���b�����>,%��rQ�����3�'?#��/!��c?O�;���
��˪=8�?�1@�����T3��l�>��H?��?w�5?�U?�M�[`<�����b�>v�?�?�0>Dz��<�? �R?s�Ѿ���t�;UD?�=�?���?$�?�]�°��Q��m�]�� ��3�'>�h�&�r>t3<ʠ�<�=P�@����=�n�=���>�ȗ>�y�>��>��>��=���|j#��%��uϓ�/�0�|_����Lń=@G:������W(��I�����/+��K=����׽�t���Y.����Ͼ~x�=�d�=��>,�=�A>y<�A�������:��E'0�A��n��a����k�QB=��/�UIϾy�oTľ�?�{���>
!�>�Q4��BV>��>��n��1Q>��>rj�=
��>�M]>���=�>�*y><�>�m>�9c=>-��B���{8�v[��?.<rRD?��`������N4���پ������>�	?@S>��'������y�!�>�OH��e�j�ν����Y�>���>'��=��W����qx�����!�=�h�>�>7������@�SC�=� �>c׾���=;�~>�$?pTu?��4?+;�=ƻ�>KmY>ܑ>1��=	M>�YV>���>��?
�8?/?�F�>��=��_�2y%=��;=��=�5�H��ܱ����_C�<�V��2=BeV=o��;�Nm=�!4={ż������<���>��E?š�>�%�>�����##� ")��@z�!�
>ci˽���>�g?��+?mR	?+B?��>�W��g�Ծ�5ؾ�U�> ��>��Z�����F������>8�=�/3?q�"?Uf�;�W�[Ȅ��>���>6k�>\�,?�J�>�>�:��U^��ο4)�v�	��ڽ}�M��-&���	�c
��׽��9���!��r�@>�C>��>74a>��/>�>�B�>�*!>� >�=&��<���<ƹ���<r=S�_=F	>�<�8���a����tu��q]ڽ�mr����2��(?]�>�~%��d<��o��d��ބ����>n��>��?���>Fu=��N�X�Q�_�&��b�>�aY?eʲ>���~�5>��S��>�Ǹ>��>D�<^-���؎��:��ȴ��iS>?� ?�	�>�/M�0�a�!lx��.�tw>ƕ;���2B�?gRT?s 	���Z���,�e�D��+��C*���&j�@��DlԾK�
�)"C�����*���B��)Nm>?��>)��?:��<����򗏿;}��Z���Ü��Z>�ڪ>/a�=#�q�=*����jf��(�ʾ��1��>+LB>{��>m�?��-?��M?W�P?CG,?�h��!	e?�=�>7A�>��Z=DD?j�b?�'F?.��>&<->��U��yY>�ǁ��_v�i�C=G�>�Q?>.��=߉>� Q�ͽ�=�v��gm�=����#�lg==�UP=1�h�p��=!�+>�?t&?r.Ž~�@�}'\��k��%Z�<�O�=0�Q>j�,���d�jj:v��>F)?5e0?���>���=nb�$���\��G5�=9�?E�,?ؑ�>`�*=��=gi꾳�q���=`�F>c�������bҾ����H��穇>���>	J�=6$?>��?�_V?�7�>�Cɽ� ���1���/�W{=���=E���X��Wi�=�����a�2w�����F��6�>�]��#޽©6<&�\><�<���=DfW>R�,>�$A�_�F<���<7�>
�	?�>6b?=�=��=i���O�%���?g����b�uo����ľ�����>0��>j���J?��>[#��4��T�Y�(jt>��?�]�?�O�?����Գ8�,э>�1w>�u�>BfI�=ľ�������>�6�>r���& ��E~�>�Ő>^ܽk�������=��Gν�	ʿd�z��݉��8Ӿ�B�<\�E�EX�~�f>6ϟ�$ �����%=�=r$߾�����Z#�?ꮾ��ʾ�肾� �.�n?��p?�>�O���`��[��$�<���_�<��B��̥�W!4��	���B�$�;�&���`�o�Ye!>�燾�{�/W��Ŵ2�CNo���t=��<?Cپ����+>��>���=��ҽ���v��+���������=?�6M?�㽾�۾Ա�����Ȍ'?�r�>.�>�0��UP��sH>#;?2�"?{{���Z����X����=z�?���?��??��O�m�A�Q�����1?��?���>Y�����̾}L�%?B�9?���>�!��h��d6���> [?GN��mb>���>M=�>��䯓�9&�L7��������9>%�	���xRh�6+>���=��>K~x>8*]�����b�>M�S�M�T���/$���W<'�=�(?��p~�=�wE>�J�>b�8�f-��ٕ���5a��O=?���?	=>?�OL?��&�/���D�=׊>���>�e�>?�(>�p��>��&?a9�������6 ?ϔ�?@-�?rpk�$6���僿�����{��J��=���=J)N>�<�Rx�=4
�<�h�?v=���=���>,t>�Ey>��+>�e>�l�=��~��^�	����d���0C��;�K>�-9���
�R|o�d�8�ҙF�zɾ7�A��ϼ¡�㤕�8�i���a��ܟ�T8�=*��>T1�>�[�>�<�f~=�E�zH)������γ�Y�`����������&�'�����\i��P����m����1?����K�C>Ȕ�>�恾�\�=�>i۟�$�5=�3�=U��;>�?�>���<Uǒ�(�+>��>EuҼ�躙؊�{��&'�<T��_����C?�<%%i�F����S���>�?�Q�>ϻ�}��8��k��>�?}��[7��u���:>
i->~�>�'=K��<8�h<���H���G?>k��>�J>��S���;]�K�꽃��=Ub�>����<�<.>o?j�?��P?��$<$��>��c>	�>u��=��I>�!�>晇>k�?!|<?ӎ ?���>�I>�<�!s�`�<��� gq��Uս�ִ<A��2ō<�=����=�G�<-*��4<S��<��#��Ӭ�=s*?�$?0E�>l?�Y�;ݾv�����H�=�	o<K�?o��>�0?(�?F�B?8��=�<�K̾ �߾�?4F�>z����ֈ� �
���e>	q>T?,B]?�y�&�"��f�>+i�=���>�z�>�]H?�>�>�T>��=�	�8�ͿJ)�D ���<>�q���:�����9�<됗�3��ԙ�=E$�=���>;o>p��>��=
"=�0ʼc��>"��=�/>��=C,=vP��N��<̱�BQ�e���=���F�������q�ٯ�W����o<�k���?��?����c��e|���
�f�����l>7��>�q#?�&�>�8�<aO���T���[����G'?1�P?a��>գ���ve>�ҽ���=%l�>Ol�>B7�=�7k���������ئ�L6>J?�B�>�x��^�	���3�+��&�>uq+=��bH�?W[?<����[D�x����B�����@�<����ח�������$��'����<���K�{��i�=��>�s�?��k���=sݭ�tN���چ��+����=><=u��>8:T>8b;��a�E��u׭�l�?��M=��>�4�=Ф
?��0?��1?*e?0-&?,0?�����Y?�ᓾ���>���>Z�2?<;J?��?2��>��>~C����=8�;��:���lF>7�= �>Z�6;~�>�h�=(�%=y�=BX�<;
U��獽P�=ä.��l�B��<x�=w7>�?��E?Ym�rf8=�􁾺�F>��=�`-���>L�e��5�?�,>�Y	?�!?m�Q?�� ?�m�=�OԾ�=V�����=��?bv1?%�(?��=��{>ʘ�o��կ<�-[>����Ps�4b��U>�?ڥ���>��#>8U=�`u>�L?��u?�L/?�j�q�k�(�p��7���=��AX<>����礽��=���^*��ȉ�|�����U�>����~��)>��>��2���=�`>��8>�V� ��=�"�={ �����>��7>�3B?���+�1=�)��~�"���f?�� �>D3�湳�.Ͼ�����>��>�=��A?羀>ca_�H$���wG�]�G>/$�?/�?ME�?q r�-�J�Mٹ>�ܐ>^8�>\R��J�쾿��O���sx�>z8�>o����kS�`�>b�>�]Ľ�f�������:����^���џ_�s�W�D��n���)���߾H��=ĽG���m�Α!>��F��ܥ����qsG�iؾ�U���	���e?rH?��=�%~��W>��ھ�@پ�^M>>���=Sཌ�޾�]������ ��x��@�	�7?-�73������:J>��{�P+|�:l��3$�Uܽ�` >�Q2?����LVǾ�g(���>n80>
���^�t���uǞ�ڨ�c�F?r�T?���'�������ޥI=Q#3?�~�>�>>��پ����q�>�%?u�?��v�v����i�����<H|�?���?��??�hN�/�A����y	�;V?�?���>���� ;���,?d:?���>z���8������>à[?�pN��Vb>��>b�>3���뒾.1 ���L3��,f9>�h
�3����g��>�˦=�֠>�ex>�]��߮��� ?v"��nI��䆿����4��z$=�I{?��1?��K��>��=�c&��Ǎ�Wo�R P?}v�?m�P?MS?�L���P��5�_x�>6�>ز?t�$���!�H ?��?�w)����ѝ��I�,?���?��	@Z��?�{�@�ٿ�0������񁚾�� >��=t�>�����e=�| =]�:옼��2>C��>9~�>��>?>e��>�(�>�؆���.��{���ȋ�!�����{I��N���3.�~胾���Y�o����O��佈�`<Ǹ�q��C�<ўD�
o9>>��U>6�>���=Gj�Y*�~4��#��^־g�����}���b�\%s�y�$��QB� �澗-s�᪾��>�싽=(>�-?�ڦ���=��>�FN>�/T>�>��>�~�=z>�U$=f��=�6>�� >$��=�]���3J�_E��U�N��I�p�X�v_9?�)ھ[L��@�J���=��a�W<�t�>
�=�*8�Ą��@���q��>�g�;��L�>���^�+>�D.>��>��=��I=4�n=��e���X�g��M>f��<����w�?w����=+��>�Ѿ���=��>�	!?��v?2�@?��Z=���>'U>쬨>��=�*a>瑅>���>b?�2?�+?l*�>.�=�NU� �=��D=�d�Q�p�Dɐ�W�X������<\=G�Wc�<���=�Xg��̖<�$\=��c�5=��C=~� ?��o?z�>̹�>�S���3Q�Z.N��֊��ԛ>�x���i?`�<?�T6?�#�>Z�q>�I3>a0�������*����>ۣ]>�Yj����A<�=w/�>�H>�._?i4F?ӑ�����?X�>�?�U(?<�>�<?�?1[>��(�^G��R�\B�2�� *��	=w���˾������S.���h��=��p>�&�>D�>�>�<�>B��>Ba�>�̡>�|�=i����J�t��;�X�<��N>*����D���X�����)����������=�0@q���:��u�2?�)?SѦ=8��A8���+��1�g�>U���RƇ>� =��彻c��P��k��6��؏>t9?t��>�H��O>|z̼f���撊>ڢ�>/K���¼�|o�]
�����=+��>�(?���>W`ɽ�V��kl�L���9e�>���=�0ݼ�܌?��8?����O=�F"�Cx�L��*�9=�և��U���վ�\%1��GL��Q��C�L^_�D`�=���>�5�?��׽n#>��֔��}�1���:�<b]k�=6z>���>��ν(�� �>|�bw������x�>5�=X�>�Y=?0�W?ӰR>g�_?�rg?���?�P?�J�&�O?r >(�"?�$j?LR?�<>"����)�>��� ��B�H�[F_�:�]7���=.�1>�I< ����	>d�=(�-�T6��6�<�=��<͊�=9x>,��=�v	?�%Z?��߽@ܠ�R����Y�On�<�B`?೰�-�n�>=u>+C#?)�)?1�?ѡ�>O=������;% ��D#���;?�́?"??��I>y�f>�<���_����=ճ�>�D��E�����Jh�����"�=�-o>Ic�>��>g �?c(?T/P?�.��z2�f�w��l�r�L�x��\N=�R��
�=��	�Z���䡿Qf��\UZ�88>E�R�hE�=%z%>랊>)��=�CS�84X>�e��ƹ�>���_ί>�^j=���>���>�?�>Jq�>~�=���;.�	�c?l�[����]�1�>���w�x>��>`�c�;y�?��Ž�̐��u���Z��׀=/*�?Px�?�?�?:�m\w���!>��>I��>CX'���Z����w��8��=c�	I����X��=�\>�KW=؏��L�v�&�^s��j��MM�Ag��bb��&��������l0�=��ྕ��:@����Ҫ��{t���!�?�y��Q��g��q���2�?��?�� >�D�󳾝D��^&���R>X%˾�Yw��i;��<Nª�_������d߾�4�<XB�Ʈ&���>X�8�V�r�.���Q�f��[�HW?����N�9�>�{�_>���<��ݻ$��2���֕��5,�R<?-�>?񊆾浾�^�!V߽��,?���>��>�,R�N\�>&)>#y5?<�/?��t��o����e����=���?�.�?\�>?�@�V�>��{����'�?��?�T�>P��j�ξ"���	?I�6?K�>dZ������Yr�>�>\?KM���^>J��>*C�>XZ�((��
�;��������;�.>R)[��e���d�sA�1ַ=��>'	m>�i�/W����>���K�=6�,��\\#�7�˼'��>K
���%=K!&>���=7!,�a�y�uٽv�L?���?:!J?�N5?%�ɾ+��=�F�E�<dh>��>A�<��>���>���>�����w��;���?��?!��?��[?��l��տ�����ξsY��fa�<�&�l]�=Ľ�"d�!�����^��	>���>���>���>��m>��h>Ou	>�b��-�%�U���鄿>6��_��0�W"վ�J����Vl#�	���3�����=�A�=�H�=�{���!�s��%A��<v� ?�s�>��>�[��<�1�yl����-����H����<5��*��q>�zu>u1>�T�T3���޾��?�����A�>�D�>��=���=�!�>r��>ؘK>7��>���=8g�=� >�>�j&=�R�=�Iw=н�>@��>3���>���aǾ/����$�h?��>���<��,�ߚ��������=�Z>/�=|�9�ɡ���c���?D�=��ȷ��ǔ�)�>��?"N�>��Y�MS
���O<Cz��)?(��W5>�e�>��������m���9���>V�U�>���>)*+?�u?��)?3�Z�Y�?>CF�>�I>f��<�@��lc�#I>c�>c�%?�?�?���=�9ݽ�
A���/>�긻p6�c�U��@��u�Q�j�R?/=�ȑ=��ν��O= /�(�/�V=k��=�� ?�GJ?��? ��>�_%>+�־��"��ST��e�>6��>��>���>�V?2P?�P:�C�o�&o-��N۾*3�޸�>1�>Z7]��=z�̎��?�V
?��?��0?IEo��閾uH�������2H>0ŷ>ń;?;��>��>��C>���V�ٿ� d��T��7"/����,Pپ0~�<��+�y�;��=�뢽C��H?�>X7?Xe?d�y>��>n�1?��>�PR=E�<<>�v�ji�=mnB�{N�=U֊=2�K���/<��;�(Ƽ.��E�!�'����+���q��b�=8�?ٔ?�$v�D_�9JO�T�Z�����>���>�<�>�_�> d�=%��7�Y�/)<�~�B��5�>@�e?@{�>�u.���=G�-��B��B��>�j�>�D>��K� ��?ё�P�b<���>{�?@e�>�|�k�R��Zj�}���͠>�1�=��轗܀?�L\?�ꟾ�J��I:����yyٽ���\x
:K8�
�4��1B��龑�[����`/�g�>/м?(*���>�r¾=u��q:���K��<��A�F�>'Q�=���=~å�x�#��x��~���,}���<yH�>A�>�N,?�q�>u?�X?�O?7��=@T?B�>i?I�>���>���>G��>���=�x�>ؿ="�'�r&ӽ�����i=�9>`P>=����(�=4�����L�4>�*>l�w=#��'��/1O�%^ǽA�=c>�=r�'>��?��?~<��ɪ��5��{�==R�x>I�M>�4k>�W�=��&��M�=��T>y�>��?Dն>��$�>�/4Ͼ*"߾q��<�[�>+�*?WM"?�J{=O��;�b ��l{��@>��v>N���f���n�S��E�@�v>ޟV>�����>��?��W?�C ?Ip���I�����Tid��2�h�_>�&?��6?	?;��s�6�{)i�S`c����S���/%��'>�]P>�+f>q�!>��=z@���d۽�%_=�J>��>�#J=,^�>	B?�
?vΐ=r�>�Vf�I�+�?�������h�ܞ���(x��;̻�D\�<Ѿ;6;>�t������F��[�D��+�>l��?f��? �q?E)����R�>��>�2���Ⱥ�����=��l�a�d>0�!>��%��>)(=��k>���>����xβ�f義����F���{<�4Z��NϾ� L������������h�6�+�G� �B��l��!�3�����ث���8~�K����!�?�m�?W>B�-����B�۾o�վ;#<��o�) 2��ͽ�x
����E�����D����%�w2��A�!1H�Ӌ?\�#<U��������3`�td�=76�>��?�+!��M侤�ž0'>���lO>���/q���~ɿ��d�͓?�#?H���Ӱ���nO>=����	>��?$$�=^���.8��ס�>C�N?�<?��=lA�����[h�q��?�ݿ?l�B?��r=��<��x��H�A�>�l<?��?_�3=�b龹8	=�0?ǡ/?D0�>+Tf������:c�e\6>�0?��pH>�;?���>$\U>du���	�0�оf- �E��>�ս����	>�6�RA>N $?�P4?t��(#����>>���N���H�W����ݗ�<��?=��~2>�i>L>t�(�l���ω�`4���L?���?�S?k8?/\�����֫���=]��>Ӭ>���=�����>���>Xa辽ur��ۘ?I�?���?�XZ?��m��Ͽh���V��^�Ͼ�14<�o=��[>M��=;��<9��=I�=�\=�]>���>'Í>�Q�>�ǋ> W�=�@b>H���p2(�ѭ��>󠿇�W��Ӿr$#��t���������ܾ���;�?s=āv�b
>A���Ս�#��Q7N���<o�?��>���=��>�p>��j=G���g���!��ŢZ���s8�H�%��پ�31�E���y�O��58���"���>N�=�Y>й?\I����W>F>b�9>��u>���>�B=��@=a�G>5&+=ۄ>O��>f�>v��>��>����^`���;�J�������?qu-=�Q̾쟃�y����)� �*�4�������g]���W�F������> ڍ=�4`��h���Ⱦ	�{>]?\y"���l�㽾�:<=�^��.c�S�>�11=}u��Ӿ������C?�0s���>��>nE? AO?b�+?�q��q5�>���>B�[>I1<!ӝ=�%�=�-�>S��>��;?HOR?�
?G�=�b���#<�����=��{����K��<�_=��>��Q���=]S>� �7��=�:1=e�%>��<���?��9?]�4?H?W���B���.M�<��h�Ȯ�����>b�?�c?�:E?|t�>�Ӹ=���U6�.�Ҿ��>�8=�J�VsT��0#=��?��?��?�$?�(��� վ�N�{��=��V>�F�>�-?i~�>a�>�6>Z����6ѿ��r��:������<>\~��D>�M������$���l&�P�3�V+�>�?�!?�'>\U�>���>�m�>M�l>��=y��<c��<���gm�<�B�/̓<�`Z���2��[�=��@����}�R�{��0�;p}�<��;�??�;�<[�<���� @۾U�6�_J�>��>�.#?�`�>�Yl=���~�U����_B��' ?�lm?\\?�#.��a=��`���<�P�>K7�>Qy> �P<H����`�����;�?%*?۰�>�6p�nOa�ٟt�y<�@6�>��=����?a�Z?��"4��3w
�VWF�?��q=�r���R�����B���S��sF�Y��7=R��>�w�?i���>2Ծj���%��ۍ����䦗�~?suy>�xѽ��o���� Ǿ�v����|>Ɛ>1��>��,?��@?t~T?��G?i
?�BU��|?�K�!~�>M�>N��>0?��>�H�>AŞ>�[�=U5�=+r.�M����&��Q�;��>;M�
�=�¸�q�J=C�>!�=�r��d����=B�9=��P=�%>�J�>�p�=��?G?��'=ދ=�	���7��Q�u=�ѐ<x�<>y$�i.��d��Zމ>��	?b}?���>�B��z�����Ҿ'��Q��;%�>�%J?�?�.X=�|�=�H˾8���S�:>I݌>�%��Í��J�'�y�r¼<���>�Ɲ>.G�>�\�>�.r?Z�P?	�/?Y̓�!*7�qEr�Q���܀k������2�>l$�>7��>h�U�aX꾒^�F�x�0i��f���*�8�&>|�>��<}7�>�A�=u��K�f�e�𐽳�q>k��>��>�??��>z5�=4@=a��S龊�I? ?��������޲̾N��=�>�;>�C���?O@�f�}�[r��і=����>��?�(�?4e?�=��?�[bZ>�)U>	>R�M<�B@��'��X}���3>$��=e�x�8%��|F�;��Z>_�p>Duν�rǾsP�bH5��=���>�˜��������z����5�:>s�>�vx>�.�=4�Z��g"��C���*zO�<���̾,��
��?��{?�)�=�B=�;�;%�+�,���n���D��.};����E���^*�9ၾ����]��~O8�6@�L�d�T�>�==��(���g���$���O���>!%.?���,?���<#��b=Ӊ >�������h����t���C?z�8?���9��
���=�n?�:�>�V>���(�*o�>?�)?1�?��	��b���N���ڼv�?���?��H?s}=�R�B������F!>&O�>��B?��?���e ��Cu�<��U?��!?ݡ?����m��4��*?�b?���J7�=Z��>1١>^���{��u彡�|����;��>�:=�ۊ��P�t,���><�>�->�̝��3޽���>l���N�X�H����#��h�<�h?Q\�>ai>%U>ܶ(��	��>ŉ�J����L?|�?:pS?�38?;I�����夦�9��=�^�>O��>�Ů=v��'�>%��>ڪ辏fr�_(���?�:�?���?�Z?хm�O�̿Q���Q����Ӳ��H�=?r�;��>|�	�O'={7�=����c�t$>��>X�x>�AH>=�7>��U>Mg)>r݊�;�%��Ȧ�*��}�>�(�&��U�2f��$[�6be�������o���e���e
:���=;W�rd��������X�>�d�>$��>.8>|�>�T�>`Jr�
Ծ�@"�b�׽��,��#�������M-��t�K�{������YQ��-��h�>��׽^;>>�	�>u'���	�=���=�>�]N>l��=| >��>̑�>� f>a�'>*O0>Y>���=��<>������i�!�u�P�L��a��?���+��_\�C�����Ĺ<:?>�>p"j��.�����`1�>A���M��e�a�	F��iZ>cM�>�n�>�H���ⷾ�@>�>��ٽ���>L��>-z�=B =�Q��=�2\=B��>zۅ��z9>@� ?�?�`?~G:?G�x���>��>��>�:B>=F>���=��&�rzE?�L?TNP?E�!?փ���G�en�h�;t� B2�\V��@���<���W�J�a�v=�r�H�սd`f�PrY=x��v	;<��d='�?�:5?��?L?^�ƼX(�� L�!�þ����.={]�>[?fM?��9?7��>��>���F�ݾ�"��l/?>��>�.��)����;<��>��?�]Z?�RN?�����Ft�L�I�H���}.>\� ?׫�>|�?�=�>��<>c���˿"�m��zQ���=2�`�B'�K}�;D�*�͢1��C꾾Sc��Y���9�=��>z�9>��p>�F�>߸�>���>St>�N�=P��4 M>�K�<� 6�VL�=,���F�S�򽨠.��!5�X�����a���)�o� �U;4���?d *?'=z�=a(K��˾� �E�>\��>�
�>^��>�tļ���7�b��5G�e����>8(K?"y?Zʽ�]�=\��{��=��>��>���=����$fJ�Y�3�=~ܮ>9�>�"�>r�;���a�!3�(m�ː�=��=wE��6�?�R?˦����8�,8��4��#e���=m��=*i�=׾f�"� �>�"�B�B�	��~t��� ���>���?s}�<^ܒ>�V�m��aĤ�ŝ��h���V��;��>�E>�u>	۽�.D�zi����G���O����.�>��?�"?�?��.?��?O�?�����?q+Y>��>`L<%��>�w�>��?}��>!�>�3>��>6	4��a��wy�^=��#i�=��O>�>��=���<5�v=0��=<���I��GҸ��8]=�h�>�/>��4>K2�>���>��"?��%�V���8B��=�	>��N=��{>ҫ^�;�彀а�9m�=e?�>ǩ$?�"�>A=ټO�žl_��}3���N=��?��5?t�?��s>8	=���l,־'K�>��L>g9^��'��N��W���k�+��>%a�=��Z>uj�>N�6?��f?��?lx���Z����U���߾���=U��>\��>�?t���w:��@l�L��\�⦾R��Yy>o,�tN;��V7>���;P��=X\�t��;6W½i�9=g�<,��>DJ�>9?��{>?��<b䢾�Ѿ-�I?����=�������ϾH#!�l�>_=>{��T?fg�п}��ǥ���=�9��>~W�?��?�d?��A����Q^>�W>�L>�k)<�,>��F����K�2>��=��y�<C��84C;��Z>��w>�0˽��ʾ~X��I� &��\g��¾�R(�e������¾z�=Z�s<Yм�?��2��Bف�����ON��@�U�������C��B����?�3?�E�=�ۦ��� ��\Ծf������=cG�q�(�㾹���g�Y��q��0����=���B���U��7��7�>���f���#>��2X�q��� d>��?�<���V���߾��>�n콵O�>��������<��E⿽�> �?}`ܾ:���U��=�F��>���>��P=�ֿ�9�޽6�>��:?��Q?c�S>�c���c;>>��?=��? o=?J��'D�4��־�+�>#�
?��?1���+�<
ٽҔ?:&?>6?<�s&����5��2�>q>:?����Y�W>J�?V��>Q�E��~"�Lz��I��c��>1蟽����.�R���L��<Ho�>H�>����{=Z��~�>�+쾋�N��`H�����o"���<4�?�%��>�Yi>��>d'�97��/艿N��LL?T"�?��R?�8?L7�� �㠽�M�=f��>�2�>��=�D	��P�>Ą�>H��0Sr��_�6�?��?���?yEZ?p�m���ʿ�[��bQݾ�fƾ\}�<U��%�>W�����j\<�ڽ�&>V��>Y��>y��=`��=(IO>��0>U�>����g'�������H
Q��0D�)�(�b$�����վ�w
��{�wV���t=%%��yy��;=7�K�-����l���B�/=R�>�g>خ>G~�>n�,> �����?w����c��\!��վ�����˾?43��]`���E�� ��<�L�,?�>\�>��>�J��[�C��>��>���=g�>b�==)�=�.>�T�>�ŧ>�B�>[�,���=�"�=����fj����sl���w��X? X>*������jϾ�����
>�'�>3�;��G����3����
?�M=ןǾ�^J�.���W>��?|՝>'�=�-���m��\��TɾH��>�+�>�Ť��6� ��s��=��?��HO�>j6�>À
?�jW?!:?��V��D�>�
?Մ�>!�<�>�c2��>SZ>?X�H?��.?"�3?gL=�}��!�ܽ����b�m���Z��=J��=!�Ľ Wi�����y�=$�">f�8�ُ׽Wٝ;�����J3=&�=�?#M9?�,?or+?�J���5�y�K����/����Q>���>���>S�?�
4?X�'?�s<*
}�m�곾=��>�h�,3^�O� ����<�os>'x�>m�^?B)?����nQ����d��Wx=�ؿ>��(?:�??>��=Q����Nӿ1�?��)�ܔ:��P��Զ[��o������s�}�������\���s=��D�o�߽�٦>[��>ȋ�>).=���>q�e>Y�=_EU={kq>�	�=�}"�g�º���<�ra>�w��5�5E{��z��0����;P���=bذ��\=#?n?����w��_��[���~��Q��>i�>��>���>rT�=W�4MU� �@�D���>�h?���>S�9�&q�=2�0���;h�>���>��>�yV�@c�+љ��<8�>n?zԞ>H��iZ�X�m�E��4l�>){�=�����?=nj?帾�������N������C|;2⢽����iȾ��'��[0�����[̾�9K��2>OZ�>�ߦ?_��]S�<w�Ǿ>��pl��Tʍ�J�<ZG���>/��>����qJF��V����_�r�� ����==�>Z��>�&?:*?�S?�i;?ƣ,?n�`���?`��>D��>b�F>ّ�>���>2?��>�o�>�o�>ʕz>�����s��x2=0潞��;��>o�=3���t�=���=�-�����&��FO��j�����<�Pz=�2=!">��?�u&?gH��	
>^ؽQ ˽�m>*��=!�6>cs�p{���~-<���=���>�:?��>�$��P� ]�����>(4�>+d$?�%?7�,>F�q�hX��l����h>'-�=��>�]i��,v�=S��
p���`�>w�>�`;>��{> �?�vk?pq:?�[K��&��%����i�[XA���h<c$?�t?0-�=w5����2lw���G�QE��4;��B�i�k>t}�>݈�=Bp>1JZ=#s����8_�-.>�qz= �M���>HM?��3?�J'>y�F������J�s�I?�L������� Ͼۇ��J>�=>9-�Y�?*,
�W2}�د��� =�mb�>p�?�r�?Qc?'NB�v�][]>^9T>�w>u�J<�;�E���F��Ӄ3>�k�=Z�x��j��
�X;�cY>�V}>�ývV˾��@	@�j�����K���������G�D���R�9������S����Ӿ궽���Gī��þm-K��U6�����i��y�z?��q?V��=������X�9���->�ͱ�dI��7���̕��Ȁ��,��Z<��咾��/���A�0�E�n>d�����6����R��̵�)5�>[s?�R1=�TM�Q�2k�=T�:���>�������d���Ľ���>��>N5����d=�eϾM�'>�J?�\>��A���>��7?\�?�ji?��P>8���a�X��c2�,�?V��?T�>?��н>�1�c9��� ��s�>V�$?�Z?�����N�v��]��>��?k)?^�M�����A�oY�>�V?�����f>��?�?�޽� ������
��L����>iT��z0�G�D����w�@=���>_5�> ���Ѥ/�;�>/����N���L���վ��(���[�o�?h�ʾ�$>1w>��=z�%��1��(݋�`�H��=W?ӯ?�yN?�"3?H"ﾰ���鮽`z�=�>�4�>�=�Vܽ&\�>_=�>�WѾV�R��&྽	?/��?���?�5S?OZY�|7���9������&��f�l��zC>+�>�H_��qj��~�=�1ǽF��<��=4I�=��_=V+>�;>�U>��_>�s��ͯ$������aQ��M
����}d��S���䔾��4�i�ɾq嶾�~�WUž[�5�Q�B��}m��w�T��7~�����>́>즥>z �=��>�� ���龺�P�ξĎ
����)��U��@T۾S��*ؽ��9�gF1��\�����>�x��?��>�f�>d�5����>�w�>��B>e��='~�>8է>#@>��`>��#>���>�G�>u؞>F��>!k�>�g��Ϻ���Z2�B���Z���.��?��>�[�yK�?���*��M�>0p�>B�?��y��ڝ��������>�u=�]�s�V��稾�XH>�03?�ը<ޫ�r�þɧ��+q��S��=�x�>��^������ ���+N���x�{?�U�[z�=�ˮ>x5�>�ay?TF?Ϯ�=&CB>'(�>��?���=�>�+;",:>���>�X=?�YG?�?�C>.���)ʼe�>1������O��i��>��=���=w(�=��>�bH�P��<�}�=���1��%}=�D�� ?
e?��.?��?ש���?�Ũ0��n���4�=��<�?��?��B?��%?�	?��7>X���*��c���Xc�>c|>�G��}L�%���g@>6u�>=i?0-6?K���[���J���)�:[�>d�>~8&?9]�>�[�>d6~�v3���п����on����4��q<�Ƅ��FD�_=��[Y��k���������=�� >�q�=.�#>�H�>��C>]1>[����B>}1�#����}=H�=Y��=i!�=0~ݽ�3�����>�!�:������=k�����?��?^��dH��8���_S߾d<����>M;�>;?6A?���<
���S��1>�=G�}@?^�v?c?�^+��x�=���<�{L=�q�>:��>��G>�d�����J0~��ݏ��B�> �?�$�>���
^[���n��o��j�>���=�6=���?	;�?C���R;�����
V����&�9�<b:>f��M����f�#�v�A&F��0@= ��>N��?�e�;��=��;���`�!}��&4�#!��Dm�=�u\>�4>"�=�K�y+���'�׾�S�����=?�%>�P�>=F?}�?�K?7)?�8�>*�jy>��>x��>���>�>�6 ?��6?��>	�m>�o}=W��='��F�r�:����;Xz>��V>��J>�FX=Ϯ�=�L�=�p�=��B<WcܽK�(����=!?3>YTR>�&4>���>�%?N�-?y����L�m�G���X��.>_K>�i�=��L�9�q��!���L>�?�l?�>�`H;U�����/��:=��?(%7?I�?ȾI>O�<8��l^�N��>g��>��s>��Y��>�H���.н��>�!w>xT�>�f>F��?�Id?��!?�N<E�%�$j����i�{5��c1>m�?#��>���>Y����� ��'��J	_�JtL������t��.m=:��=�+�=��=����T>�C!>�#�<k����F�=�����S�>��>�9?'G�>z�>sϬ�e���J?ܚ� �����x�˾?͂��4>�?>t��(?fӽ��y�TU���-:�z��>S��?b8�?�k?4������Q>J>���=eO����$���ϼ��~��FA>*��=��S�>����~��1>�qm>�?�P����̾�ޛ��Y����`��x��_���5�Fy�-��l�<Q�5���<	�$�Ô[���)Qͽ����^���w��y���:���$v?V��?3Ȼ��R�E�5����k�
�&)>d n��v[��x��>o9�����
�b�����(���)]�-�_�) 3�3�>��/�?���M�|��jI�S���$H^>�/?[n��7�T�����"�>� �=*.
�����퍞��,�<"?)#?�Ͼ���W��8�=�'�>�]�>eSk=�S��I���>��>?��7?�5~��݈��?���=���?`g�?E.??oF��2@����X4�~?<t?w�>����z�Ծ�'����?�7?TA�>����]��c�}2�>'>T?��S���c>�&�>�>������9
�t����弅(L>��9zs���Y�VUI�W9�=P6�>��>��a�􁠾8P)?9�A�y���W���G��j�>R(�>)>;�پ`9��g�/>`�>Ě�h��J7��ԡ�sMf?6��?c��?��?�������t�<M+>�s>\�>�^㼒����
�>��%?5X�~ R�`�c�'�>6��?�s�?م_?�u��ܿpޡ�����Z��"�>>�_>���=h<E���	>ŨM;<[<8��=�=��>-�F>D�O>Z�*>�(>	��=�w��r%�N҅�o�%�������}����펚��{��$�Z����o�������O��E8�����*�}�W�T׿==��>玆>��x>�Ф>�L�>�А��L-�vls�R��+C�DX׾���&�f�Y�VQ!;i�ټ�$��ω�,['��QU?�*K=���= 5�>���=��Ew=h �<�d�=�=�>�f�>�g�>�8�>|y�>@��=tW
>��=��Ͻ�̧=]�N�V�f��_C��_D�!��Bє?�˾�����p�z�¾g���ή>	��>����Xa��I��Tyn�	��>��ɽFpP���>�F�=�ȇ>�X�>�N���K�=�W���0�gmԽ��=�V='��'g=
����q&�+*�PP�>�y޾�N)>�F> 04?D�{?�V:?�8��V�>p��>"t>S_3=�>�S�>���>�'?J9?i�(?o��>�C�=\O7��"�=�Ō=�o;�4eo�P����bӼ Ŏ�'U��W�ʽLv+��4=�ji���|m��Վ��C�=���<c�?�R?��>��?q�3�8��(h���;�c��=��J� ��>�g�>{� ?ET*?r��>ݜ/>����
��G=��]�>d����(��]y�eb>ī�>ご>/C?�b?}��yܾ/ꌽ�O��u��>v�?��?��q>8��<ƞD����FY忄��;��;�1<?w���4��CF�����<�ڂ��2u;�a�=ݖ>R��>�`>�5?>7�>Qw>n��>��T>�wټ�\��w��E������="À>U�޽d,�=��t�?����<;C��M��=�-��s=�(��/>�?�i?Z�ѽ�$��"Υ�]����u�ļ�>�m�>UC?B��>^S����_��`��z�� ���i�>a_?���>!+W��3.>R�ǽ�����?'t>���L(�<���le��i�>�I�>�?Q��>����5T�Z�k�Ӧ��Im>��>��!����?��A?xY�J�V�9����/�:X���<�>O���~��ލ���5�F�㜴���������M>��>�c�?� [��[�>�n�Z���ޤ�n��W�?Ўv>m�(?9^J>�_�H���Ц�	\����Ș��O�>�^��>> K?�?�l�?s��>Z!"?[��ʘd?�����Q�>�x`>Ω>c�?6"+?��?5>w�)�?����z�@�ܲ�=���*�9=0�&>�_~>T�|�.>�Y>��4�jF���H�=H	>eh���q=�ٟ=��=[d6>e�?*$+?������>G�y>�r���ӛ��Z�=h��=��g��f��(>RK�>.�.?�wW?���>Ք�ut��	����?�{��?��?�-�>g��<��b< �Ҿh�K��H�<V�>�)=Ѝ���t$�ZS5�o�5�HА>0j�>pA&>��>Ӕ�?2dP?�?L�(��&�<���&�ջ��F>��J?�h�>@��>����T<��ܐ^���_�s���ن<LS��9�=z>��>�>�b=S�=裔�={��'�����=rߡ=l��>OZ�>u�?�Ox>T��=����<��%X?\R��?;2��ޑ��a)�PP�ٶz>E)G>!���-2?6�ٝ��n��V�v�Z`��?Y��?Ϩ�?�5?�4���	�>���>M�>��<�q������Bx>�S&>�L������@���==ݥ�����Pj�K���N��qſ R�D^t�H�$��E¾<>����$ݙ>��پz�(�)�+.��HV��M	��:C=o�}�Ӈ\�0,þd�D����?14�?o�v;W;q�]m��3M��/��>�,�.I��.Ӆ���s�t�ؾ>�þ������VI�ţb��.�<}>��p ��@_�r?��p���P=��r?��sp�|D����=p>ּu�u��D��ہ��n�O��0�?`]?�8���?.�r1�\�^��V?���>:�K;�����9�;�<`>��9?W�"?�V��֡��ힿ ��=Z��?��?�@?�2Q���A��W����Ћ?��?8�>�����k;~W�I?�9?��>�E��O��e��L��>֧[?N��db>���>
^�>"D�䭓��&��Ò�K����;>��������Th��D=�9��=H-�>�py>c\��}E?�_2���o��dy�̂-�a$]>`�>H�M>��ھ�����^>�E?Xg��������������R?���?�jt?��?#A��H�f�f_�=aTo����s7>Q�A>�0+�o?�[?6"�T����$�&z#?x��?ē�?9�?����EӿB��D���}��w��=�=e�>>��޽�ʭ=�K=�6��3p=��>S��>$o>�>x>~�T>|�<>4�.>ؤ��v�#��Ǥ��ؒ�ZZB�^��L���ng��x	�Zy����ʴ��������֓�^�G�Ѝ��6>�9{u���<>Tq?Vz
?�v�>Ț�>��>�y漓�E��
̾�㾟�޾�ƾ����	��*}�vƽ�vD<�k5�pf	���>�k�8?�d�<��u>�}�>��?�-9>��>���=Z>�=�i>�>�Ѭ>!7Y>�}�>�s�=���=0SP=�x3>�w�=��l��,z�r��A��G]���6P?h}Ծj��|J��PѾ����g&�>:?�@>.�g�!Y������,I?� �J;;�>���_Wt>7��>r�5>+*>��f��A͹=�!>g��=e*�<�uq>�m��׬����׽�X�>�־%�=<Ny>R7)?<�v?�$6?^,�=sE�>��^>��>:��=��M>�QR>�>��?�9?�[1?�!�>;��=8�b�g�=��4=^t@���_�7���������(�>�<�
.�ʁB=��s=�<�e=�MG=�t��db�;��=�?\�2? ��>��>�n����c�0� �4=�I�=�@W>�?�C�>!y	?zx�>�f�>�nE=�|����ɾ����3��>�3�>S�=�#V|��9ѽ#�>}	?3�M?Q!?����ֺ�؂߻��?�?n\M?��v?��=L�@��ܾ_Z�x-�6L�6�2����"��b=��G�೽�'�<�����J�=��>�9q>n\>��)>��=�)�=���>:8j>�z,��U������u�=�Væ���{>(��5>��Y=�C�(������$߽:=�F��@���QB=G(?���>�V���I�=������Q^�L��>��>��??e"?�1->��-���f�G�h��վb��>Y�2?�!?q����G�>w�x�es �A�>��>B�%>t���H^�i>�\y���w�>:�?���>m��`uy�y���.1���e>��'> ����+�?�k?V�]|��~�%�I0%��%��U�>�΃�j����w�FL5� T��ɯ�܍Ѿ����X<>U	?d��?C!���=�4�_9��#�v����>�>�N�>�?s�G=Z���&��N��[�׾�ѐ��`��d�>]��1F�>��k?�$?���?ڏ?�?��FN?������+>�yA>��&?�\?�u$?�-�>P�'?� �=gs���"��۳��[z=֐$=�{�<R��=�L="���%��;�Fj�&�=���=���q�(�����w=��=��.=)��=�-�>�!W?��z�퍄=e�<��>%>8�>�X�>E��Xm��>��C�>s6?�&]?EC?h��=�� ��^H��SN���=Z��>�c�>�?��м
�;���{��w��\Y�=X�B>�����ϧ�������@�����>�r�>bɇ>�}�>~UN?���>�o?�� �g>-��䓿���}��MU�>�?�C���le�*���衿P]Y��M�f.y>�D��J�m<Iq�>\��>�>>�Q�:{.X>$�k��Q7=�A�=H����#>��3>�8,?�aK>;I>E�<�`#ܾ+�W?�־�u�qO��/��QϽ��V>�_>>��0��?"#=c�n�&ͫ�9�b���Y>�?��?��?��Ža��˳�>��>���>��<kmo���!��x=x�C<E�Q>�b��H
̾ˌR�H-4>� >ъ���� ��ѽ8Iǿ�`��a���/������"�֜ �H=���Q�x>��F˾�~ʾ��(�W�N�<�Bќ��,��8��2�?�s�?��=Qt�F�?/��s�$0>`hྲ�ǽ��ྌi���ƾ��پ\��!G	���?��K�����M�>>���*��E
��x�:�r{2=��	=?"�׾մ��7����>C�q>7���}�]p��m����U@��KW?��L?
3�H���w��Q���}i?x3A?�-G��Z������f>IFD?h�C?Z��J�����V>���?֥�?�D?	w���J�]��<�@� �?�S?�o�>�Ɓ��޾�6̽��?,�1?^�>s��D��7G����>��i?�!L�?�S>���>I�>�S½��|�#�ļ$��D(���F>�ZB<Z���抾;0�7��=�ߤ>軘>���g���/�?5j ��-n��|���V �ݓ>��/>
� ?Ga�J�;�`�>/�>�X�����Tl���b�<��|?fܵ?��u?�!?u�Ѿ<+���+�̽��)�>k']>���H����>��>��'��E��8�	�m?hn�?��?�ۃ?x~��wTϿY☿�씾$iѾ��>���=��>��Q�:a�=�>�l<�'����t>�>�o�> �>&�>�3>��>����-�𧩿�����A>�?��}�-���J���Dq�����ۍ��跶�����"(��cH׽�*]�y�:��j���5��OK>�ێ>���>���>���>J$����ҽmBG�����wxO���C�W=ɾ�c�
b�����3:f\�=�����Y�Ƶ��,B?:.��6nO=Lʵ>��<=0�+>i��>�=	�>"��>�~>;��>_ɭ>t�>]�/>l�>6��=L�>�>|�D8u��92� �x���P���H?�6i��6��my'��d�T��q��>c�?;�Y>�D2�����A���͐�>��˽L����N����;��>�p�>��=��6����kF`�(���9�>�{�>7�=���<�A�:�޽�ƻ<���>�AӾ�,�=Ϥs>['? #v?  5?s�=���>�~Y>��>+�=R_G>~zJ>^Շ>��?� 8?-�1?�5�>@0�=��i�-�O=��=X�F�X����p��h�μy@!�F��<�O��
x=��[=5;�F^=��==t�����q�$=��?\ja?�&�>��>ŚC��)>�,�^�@+o�V�*<��=m8�>1��>В�>>��>��?Γ�<q���o��5'��>5@>�S��6`u�ayǼs|>UI�>>=�?0t?Hξ��E����
�(>x6(?�%?:Ab?��>��=�w�� t��Qٿ	���^f��$4�I�_�4z*��=�vA>�5�=��������!���E�">A��>q�>�>�C�:���<8��>i�#>1	��l�>d�<w,y�-�=�݁>�ey�J`�< �[�簜=(�<��=}I.���B��i"�/��;1�;%�"?�6�>Co�aJ#>����$��s��?�>D�n>�n�>v��>B�/=MG���V�q���(���_\�>��,?���>_�V���>h�9��==9�>�>Ä =O������QU�E`ͽ���>e�L?[i�>����y��R�t�b�7�s�s>9x>���7�?@�8?6��ԥ��	��Z���&��ϲ=�����P��5�3��8B��3׾���
e
����=��>-&�?�~˾�Z=>�������!
y�z~�@"�>f�v>��.?鶋><)�836���C�6w�oa��QRg�|�>��%�S��>I�c?�#?��j?5"?��V?%���MXU?���<��>#]�=?IBK?&�
?�i�>w�r==���{+>'`5�����:h^>�Z=�a����=z�E>ou%�C��=��<�aĽ�d���<ޠ��q��<�	=�Q>���=��>@�?�D?q��Ro>�[�>O�X��PR�
n�<P��<�`0��[�<��E=P�>�2;?B4?�>�>u(�Q~��D���.}����>'"?,:!?,3>[9>L��������>>�o>���=|N������덿�!Z�*ֹ>��>�|�>���>?;B?�!?RR���5������c���:�1?�H�>��?uR�>;�l�I�`�J������u��nt=��m�F�p>�4M>�9�==*�>���=>����{�/p��2Ԏ�_Q�w�;�ά�=�ڪ=�b?e�E>8�ҽ*˘�E���od?����J+���оy�9�]�(�qa->b�B;w����s�>����c���Ŀ������=oj�?��?3Ú?UlV�Ȑl�q�>��L>t�?�������}c��g�S=��>��w8�,ݽ�E}=>ؕ<�����8���5���I�ө���Ob��E��8�̾�d��,j:��M����>F<�v��]�T�9������:���?�<������Ǡ����/�?��o?M�꽷u��� ܾH�߾8���r3���z�j�0x��[�Ƚ��k�1e
���uu���Q޾1�������>eh|��ᙿ����-!F�0�=���>�?:��K׾ ���Ԥ>h�>vl���.��z��p\�G�=�t]?�l?L� �F�پ��ݽZ��4�L?�R?�L>�������t�?��W?�\?>2<�b�����ی�E,�?m�?��G?	�m�PPJ�e����D�+?fw?c��>O�������Ղ��}!?�E?���>�E��삿g����>05n?7�5���>C��>Xx>M���R�W�qˠ���N�S߹�.�=[E�=��!�tK�����>��>�ډ>�E�Gb��2��>�mᾫJ�t�F����
�4�Q���@�?z�,4>?H]>�k�=�f(��R��ƽ��و)��_@?�?�[?[L.?���E�Ծ�צ�0��=%��>��>/Ͼ=���&��>���>�7��:t����Q�?�3�?f��?SGN?|o�/�ٿsh���rP�A�ɾ}��=U����2>���︲=��<)���"x=EX�>p�>؋q>�^q>NQ(>��V>O��>B����M*�2♿�m��6�I��'�+��{s�#�����M �!��&Х�Q������Kt��)þ��-��Ӽ�?�rj6>��>���>�O�>�?��>�8I>X�i�va��� ��2=�m6Y�?��\��������=i�>�ɽх���|��8�>�Q$=�5>'��>�u=��s�> ��=ͼ>��>�v]>�R>xl�>Н>�7�=u>7��=�>m�\>�!���^��>sJ���|�F�����I?ACo�d��huP�����ꅾnDV>C�?\��>Q$K�a����U���K?���/�ԾK��'�ɽ���>��>]p�>�M'=kjݽ�����,���->}�>��3>��5=`��ܲ
��]p�4#�>#sr�el�=&�>�d4?}�m?��9?��^<�6^>��t>:�j>���=|���Im�>�`�>*�#?z<?��?B�>���:��8�!>Q�1���e��򣽑?���
�=g}~=B*�����DU=�F�I�	=���;��<��=2���t�=��?�V?YD�>�b�>4�[���5�C�I�5�k��JJ>�q�=�m�>_>�9?'��>Yo�>�$>�%�y�쾭#�~h�>Ag>��W�z����ׯ�j2�>�l
?c�p?g} ?�G��x־�k�j�>�V?k;?�J~?���>�FԽ1���9b�
�ݿ��Ѿ�%j��vQ�qս��~��&a>*5x�SgE�;��>�f�>c>?��>G/>P�>j%>LE�>d� ?.i>!����
�<����0>]���>d�W=,*
���ǽ�=�w���$��Y�=�Ӽ[T%>�6�[=��$?�?�#��x�~	�3�M��9�>�&�>��'?�?O�4<R�5�~������о�
�>e,X?�I*?URk�_X�>�Ja�(yQ<j��>j�&?/JY>wޫ���L���	�Ip�=�0�>{g�>Ar'?{1�wC���4�ͣ8�̉E>ہ)>�X��ʙ?C@6?��B���i���m�&�I�)�\��>�*|��վ������j���V�q�ܾ4�|��<X/D>֝?��?/ݗ�,�V$�\���D�|�>����>��>uA,?���>\���2;��G���X��� =�|`=8�b>�q�o�=�P?�'d?'Hc?�="?�J-?z��""?�9��u?]�>�O>g�?�T&?�!?2�D?P��=t	;��ѽ��`q=��=���<�1=j��=��oZ>���j��=�<¬�=g���=�V�oV >���=���=��?�NJ?tw����C;�;&>$_�=�=hڽ�5���M�=�(���ʲ���m>��?7�.?��)?�fF=%_о��L����������e�>��>?0A?�S>� ��,���ؾ��=}*8>��=�۾��CAܾ@r<��_�>�M�>���>E��>:0�?��9? ��>�2�+�i����|�P�����c?�>ai1?5	�>��Q>7j9�د�j΂���q�R����>��@���=�
>L>�s�>H��:�Ž�Q�Q��R-M������h@���Q>F��=�R?	�/>�V��eUC��)���I?�꠾�V�����s о> �^�>
�<>�u�ڠ?�7��}�����0=��2�>�V�?��?"&d?ҽC����[>�V>c�><�>�I��-��G&4>]��=y�B^��Y��;W^>�w>)�˽]`ʾ��J*D�ç��=�8󨾫��X-��}���5	�s�=����ԏ�,��P���ਾ�Zν�����C���8��pƾ66�j��?+i�?v)R���������*������=�=�J}����¾ �k�.�Ӿ��վ��(��ͩ����w�d;�TK�>�s�P6������s���<�1�>;�}?2ⷾ�2 ��'s�	A�]��>yr�<|��<꓿KC���v�91)?��?0оg������"k;��>\$?�=�Dp����>�ֈ>���>�(?+��#������{�=�?#��?��C?�9%��:����\��}Q�>���>�I?�-��Z�������>P�?�Ff>ƿ(��ᙿh�6�tk5?�c�?.5{�^��>`?�0�>�=���1���I����^W��>v�>ww�-tξ�Y��v!=Q?�>W�q>�N �����yU ?Z0I���{��Lu�[z)��ѡ>��>�?�/������p�>�N?8��\얿�@��;ڽ2�o?.[�?��u?�?n�+�Lc���$�Ԏ�@L>P}�>2��=�	���i�>
?���zm��z�'��?��?���?�Ay?��[���ҿ�e��������g��=K��=�@>a��;=�=�CF=�b���1���	>j��>�q>��w>@�S>}�;>7->ft����#��(��J��EsB�"	��,��Lg��J	�Ou��@�����`���V���u��%>���H����
:�j�l�3;�=m�>��?��>��>9K>��2�Y�J�	���F6��o-�(�L��5�7����H�/;ޤ�"�����vC<?.����;�T�>��F=D�Լ�7->ڊA>��9>��>,��>�[>*X�>�>�U�= ��=Gy>�<���#Wt�R~��m���<�K�����,?SľZf�]$U�U��ʎ���!�>l�?��+>��8������@��G(?	\=Y��S�<�=t��>}��>��=�=e:��G�_���轋�v>,Ų=k�<V�,=��ž�<���=H�>;�վ�O�=��x>�1)?"*w?��6?�^�=��>�;_>{Î>"A�=݊M>�}S>fX�>�	?�\9?.�0?�%�>)�=�2a�V~=�a=�SE�`9X�������C�&�'Y�<T�3���K=���=��;�:S=D6S=�f���r;>�=~�?�}Y?q�>�?_i@������D�TR}���p>�+	<j
�>���>�?�G?�A�>�bX<z�J�����G���>|3>����hf�����x.>u
�>�;�?m4?Eþv�q���5:�?��?s�*?�x>�B=ք+�(^�s,ӿ�s��sA��ʟ�{^@�k��㤅����<��(=�(���½���=k�e>@֗>Qu�>F�7>�3�=��S>�4?&]>���<Y�ݼ���u����R�j�>���`1��㸉�er.=�^�<#�;���������l����c1?���>�J���=X���;�*��o-�>Ľ�>B�?�h?���!8%��iH��7���]���>R�@?+t?)����>�YK�a��p?6��>z�D��\���?6����J����>pG�>��?�e:��|��i���5�����>�>��D��{�?|*1?*��ZOW�>��xC�=��S>�.|��I�3�޾aX=��n;��.���4ݾ#.����>cg?�3�?jWZ��l���������d�!�_�2�>��l>�}'?�FT>)"_�p;����_+�l�0��&�q��>�ᾇB�>��q?��>�[�?'�"?W�G?�߾�|D?(}�=�qb>��%=y"?�N?	?䎚>��8>Y�^=��=����˾�h>�нV瀻ck=Oǿ=�.�<&��=��=��Ep
�{�н;~����X�S=dF
>ٷ�=�'>��>�_q?D֣��/�>`�>8��=��&��<��>-z�S(���+����>*X?k?
�>>��@��#���
�2�ƛ�-�?�?�>���>qW�=�� >�����s�)�=���>!�=��������B������͂>��>�>^w�>��?�9?�M?wt�� ��@���MK���(���>W�>��?�Gm=!3��������2�w��@����>鉔�'�c>��>��>���>�®=��)=�����
�9=^���8�=>�?)P>LX?�?�>P�1>}�t�V�#�ι_??���{��" �[�?�J�i�=��>wo�>��s��'?�hv>�i���ᵿ����7��5��?���? �?�o�Y+��]��>�=��'?�id�ʾ�ˋ���<��>˅>��E�SqѾ�Y�=�=�>�5��ܐ+�����������_ɿ�u[���n�p�;���G�1��\&��W>ꕵ��!��惾w�=�B���r���y=������	̾�@��{�?%m�?vo(���=hJ���/�-�S�g>>��c""�𸹾B��stؾ ���=l��'����x.4�E�5�p��>��Y�GO���,~�D��|��e��Hr?�fݾ8�ƾXU!�m:C>x �>����v侾p��������w)+?�	_?ʔ	��z��r�M#��3U?צ?5V�=�@���c� ��>SrH?��#?���z����������=d��?4��?'xC?|h6�v~>���3�P���>���>��><O]��������	�?�}!?���>d��?D���*�M��>��l?$GU���>z��>�R�>d2��rd��{���y���?����>�'��݁��{s��i�Id>�0�>_�F>�d��e���6n�>4��2�8�|C(� {��?���8=���>����	�=�BN>7	�=�#�%]���Ɖ�Φ"��{G?�-�?�hF?��h?Mp�s��<�x�z��;���>*�>�)�;�~̽�V�>���>�Ҿ@�K�P�Ͼ��?�?�?´�?��@?�cd�#Gӿ��/������A��=%�=��>>>�޽�ɭ=��K=�٘��W=���>l��>�o>#;x>�T>�<>H�.>h�����#��ʤ�,ْ��[B�� �դ�wg��{	��y�����ȴ���ȗ��ʢ���Г�|�G�r��\U>���=����>\<�=F�1>Eo�>��	>��j>��:u�꾙̳=$����2#�H(���%�7L�����I�m���ž��{<G��꿾�+�>��F�/�=�$�>�����>�,�>���<>)|3>��->mG�>���>|�e>ZY�=��c=`p=��>�\�=5��� o���o(�B���=��-?����<�����d�
�M�˾1AK>Ԝ=?%?6}��x���f�亱>�ˁ��o�]�N��">4<g>�C�>��N>j4�� g��D.���">=�!<��R=�۔=,�>����|��U���?��>�2�t�Ƚ�3�>1k?#h?��>;�'�$o
?��>�I�.�oi�>�>f!>Qx��Hjk>��u?��0?u!��^�]��'�<\�<=�q{<fs��L��c�3:�Ku��dݼ�>�r<��#�G���[A>���=x�'<h�E���=�:�>��>��;?��/?	C���J&�=4���ɾ[��9'���?l?'j&?��?���>���=W���{��I�@ؔ>��=�D���O�@�;7��>��?�n?Z�r>J"¾��Y�c�J��-�e��>N,�>>�x>-]>���=r3�>��Kӿ��#�K�!��n��{\��ˁ;�=��L��9��,��	�����<H\>u�>�p>��D>��>O	3>z��>��G>��=��=�?�;g�:VEF��
O=����H<�LQ��p����¼�r��S��y�J���<���/ؼ�[?31?>M�a/�]�m�? վt����><��>�#.?��?|����#���d���%�q�'�2�>��?l?c���?S>�0P�&i�<���>��>��
=
r����\Vɾ�,�i��><?U��>�D�D�t��Uo�Q�O�>N�1==(7���?Urv?�ؾ�Ⱦ�Y��=t��P���NV�\��� -&=���������e��ڒ��h�:�s���g]>m��?�
�=3wG>!�־����@���L���O >э!>5�>�%�>�P>�Gw���վo$��1��,�|���T��;�{	?�X�>)x�>1a?���>��?�bg=���>�ӌ>0�>9O>Q�>�Ԝ>;��>��>eaB>W;ͽV)>QU��=���=w��=á>��=Ft>�ʁ=R�(=I�=�!�������9�~�=M�<��=c=���=��>�&
?�?U=�t��^�/=��<�ϡ�=�_J>#d+>V��<p�����-(�=���>�1?ˣ?& 7=��񾺤������M>��?�u*?;�> �X�	8K<<����\�1>�o>(/}��ۄ�Z��X¾������>/fl>*x�<B�0>g�b?�-L?X�#?/'�p�?��U��M~D����=br�=O�>���>��>g徢9���K��Uk�$j��_��_�ͺ�l�>9 �=��
>���=3@>yd�=�	���Z��\�E=�X>= �>ꖟ>��>o>&�ͼ痾G����F?����"���ھ�/���x��]N�>!4�>��˽��1?��>����ᨿ�RN�$��>���?Q��?�}�>Jr��9��U�>�:�>��4>1������p�<`�<�,�>nT�>�(���J���8=�N�=�
�
a��Kދ�&�o�em伥��� /P>۾v�>0��ɟ��R���}�%�p���;k��eF���_��t����Ծ�I�:���wZ�k��?��3?^t�=�!h>��(�o?%�5Ux�O�=��NPw��wľ5}�r>���ؾ�;i�Ѿ�fľ��y��頾���>>���R��ݚp������=e�>>GJ+?_��F� �v�)�-�{=�f>��E>xF��$�bJ����I?�X?���Ͼy�����>C_'?��>4؇>�ӊ�kz��T>�q1?_LJ?g��=�`��L}��!���ɽ?��?�h?���q� ���t�<�??�L�>�?`�V>��%��߾�v�>��)?�?8?�Œ��v��wؾb�)?d�?Ix��*>i�>�� >˿��L������tþ��>~K�>��}��e��������<� Ţ=�D�>QU�>�Ѿ�򍾄��>P{꾍O�W�H��������[�<(y?u��^�>�i>X�>�~(������ى�� ���L?���?$6S?�\8?�����d�,ͦ�|�=:,�>]�>�X�=�b�
�>�B�>*2�qvr�+?�+`?�L�?���?gZ?R�m�@Bӿ&��h���F�����=q/�=��>>g�޽��=M�K=�$����>�Zv>���>o>�$x>±T> �<>Y/>�����#��ɤ��ْ�dYB�` �*���`g�=v	�%y��������N佾�\�������ғ�A{G�є�tZ>�z�7��կ>���>M]�>�$�>��`>&�>��!��K��`���醾����_�|c���9��F�e���4�@���t����{�B�^��>`�1�=�Ƀ>iG�M��=��v>7��=��=� >�,J>���>��>��%>-�>�@d=�M<��*>�n�;����^�����t��d�������e?bQѾ����=�{d辇o���=�>�F�>��>����|�1�J����>6U��T��X���2�=t[?�np>�f=32���"���о޺���O$>�f�>ʇ�>�p�60��Yw����>�-�>vl�wK<�>��?Axv?=�-?&����9>��>��>�n9>�~>)��<؜1=N�?<�A?e�>@��>:O<�꽣L>u��������н�]�����3�<T�>Ɯ����;����G�>�@=x�*��ѻ�$(�=U��>�R�>�]?���>J���5d��&��踾[�>ƞO�� >?�C?Đ�>�Ձ>���=�Y�>�i��Ou���޾>�>�c=����k��[��=�J?A�?�&M?e>H쿾4�ྫྷ� �U">��V>=�>�ӯ>�1�>�yy>�n;�����jӿ�$���!�w0�����ш;'�<��M��ދ7��-�����p�<�\>��>��p>FE>4�>G<3>9Z�>AGG>���=�֥=��;�2;�"F���M=�-G<��P��读��ż"�����cI�H�>�m��Qټ?��6?j��=��u%`��������T�>|5?|}?�P�>m��"%�_�P��4��y]�k�>�qq?Sw�>�*l��9>Y뽑%�=\C?��z>���=���N׻��䴾{mG;��>� ??��>�j-��te�e�x��iƾ�8�>��>%z���t�?�o?�N�ʾ��>�B�j��CɾL̳>�>��[>I�>��3���*����J<Ҿk���		����=��|?~H> >�%��Ú�hR��h����Ú>���!�?放>��a�x�N��`�۾˧X��Ӻ<j�>�:A��/?)Yn>�C�>z�Y?4��>�l#?->�8?�À>�;�=b�żʷ�<��	>���>Tu��9J9>�L>�W]>_ƾ\�j���ս��)�{bi=�Q>4�>�<>�G�=l8�HrU���=�,=�+3<�Wy�n�2�D[d=`r�<�B���?�p�>��=0RY=�"����=�7>���=�w�>�j>{u�������k�n�>�?rG?
py�*���k���0O >�-?f�?u��=讵����=���Y<��> �`=k��\���� ����>�7�>�0�>ް����h>~k?u�I?A�'?5�.��49���&d-���1=\8=���>��>](=[�і)�WX�x�`���4���O�L'E���<�o�=XC�=�F>x$�=wK>�:c狽$l��)/=#c<7+�>��>��>��p>�O<=E+������4G?�cn�W��֙����A
=��h>��U>O�u<�?k�#���~��⥿K�B��E�>���?��?�[?�nP���,�X,�>��>�y >(O��e^���w��^�ΣY>��=�}G�;*l�/a��N��=K�>�'��ҭ��瓾M�1���`�A����ʡо���� �m�����C�	��E����ξ�v��O�Ǿ҅o�0�O���y�=�/�G����?�]?/e�h|�=F�A�)t)�!Τ��o����E��Q����X���5�$q\�3{��� C�lþ�P�a��'܍>7������+=��6����*=��ڼb|?�"�A8��E�r�+��s�>-��>��v0������l%>�C?�J?۩����ZB,<���>�~�>�@�>��z>��=�i~��r]b>��.?��l?�q~>��\�IQ��"�9�4U�?�(�?
� ?��ʾ�+���Gn�>m�&?��>'i?*)Z��qr����J�>	W?�N?[�d�!4���Ⱦt�?��=�F��2��>��?�z�>}O�:ot=C*�=[�Z�6�>�?��o>7�L��k���Ծ���=�&?�φ>���ej��{�>x�zɌ��7�TV�3Ճ��f�="��>/(�{�>�X�>�e;u���p��䒁�cb�G�?���?��?�dG?�8�˴𾷚�<��>~��>�zc>�SV>���=?�>������ �Gܵ>24�?(��?��j?�%^��Eӿ~������W��l��='�=�>>��޽�Э=ۭK=z�����<�1�>���>4o>{5x>]�T>�<>��.>������#�zɤ�>ؒ�[B� �ã�x{g�|	��	y���
Ǵ�B�斨�<���gܓ�f�G�ь�s>��X4����=D��>U��>l��>��k>a+}>jI��M�о-����k޾�ݾ
#��N޾[o���G����8�h���:�S�����W�;���>�����Y>��>�k�$F�=2��>|�+=�3>�\>3h>��M>(��=��q=nI�=�m:>E{�=�|�>���{�{�ֶt�:m�c�i�a��=To+?�%�U6�O�A�w|���9�>��4?{�>�:(������k� 1�>�>P�<����&]���*>�;�>7�S=]�{>[M�6(��v�;�:>�K>�x,>D�ؽ� ��z��;&p�>I��>GQ��;W�= N>+�?q�?�(?��g=��>��P>�@�>���<m��=Ra>R�>6'?98&??(��>�P8=�RT�V�o=+v��,�b�]�`߽�ډ�!�6�yrE;6�k��>�E>[����u=�UZK�M]���G�=pl�<T?�>�%?[�f?Tc����0 �"r�u��+羙H�<&e���?5#S?y$?�w�>�aʾǨ��)��%6I>�=><�`�%r�{j�6�7>���>T�?_?��\<Ҁo���t��l���89����>�?޴�>�)�3���*�r�����޾�`�𝊽
<ѽrl���,�@C��U�j��C0�R��a�O=�>�΁=���65����=<��0��>��>>RJz=��*>��{�B���<����=�*'����=q�����!z�=�Nx=m*��R7~;��
�'�J�c,=��?��?� C��	о�C}�j$3��c�=BS?(A$?\T?$?�	�>%A��Dm��=t�zj۾٘.?jU�?Ϗ�>d�x��P�>LL�=c\>[R���ཊÍ>�],���|�n =�j=B?�j3?6;g>X+��o�{��Qx���·�>p��=Q.%��@�?�O?���d䀾#Y=�K�a�le�{a���Ǿ�`u��d���忾h�پ�7ž��
�ymM�!\k>ב�>[�?�ŉ��T>���xI���7������(aƽ��q�m��>���>;~>/>
����������W���(V�>'U2�`�Z?�Na>��>��r?ҟ>aN?�+@>� ?�'�>.?BG?��?��=
`���g����>�P��hc=�k������˼=�<�N����<�	p=l��;�ѭ<Ѵ���~|<����-�^_o=YW�=��2=��y=���<p%c>&H?P��>�8�<��q��a=��m�{q;=�U�>��b���ܾ'���3��Ӌ�>�q<?��0?��_����劾_��+�=��>��?c�>�>U�<��,Ӡ��,=3��>)筼����E%��*�վ�����>Q�>(���ޙ>��h?2>?Pd?����o��Rf�3�4�.�����<rfx>� ?�]�>-�5�o����l�̖U����]�>����y>�1�=~�g>S۾>�pt>���=�>�;�ە��*����<�m����>n��>���>Es�>ă=c;���徏�A?�]��}],��d��7�=c\�>)��=ϖD>�0G��>��->�o������#����>�?#�?U�2?W\���Gn�佔>��;�;=�Y���c����G�e0>L�/>k��K���������> y�>�ڄ�;������x�GEÿ����*=��]�
��b�UQ��m7*�Kc��vi�M'�Y��d���ս"9R�娝�U&��gy9�(S,�Z�?�d
?�%l�A~1���'���Z�y)��Ǿd8>�XJ�� n�*9X������۽�R2�a�w�@�ž}����+�>�t��뒿�]y��r2�@DN�
F@>�[#?i�վ.k�������<�>�D�<-ӾԽ���������0�O?h�>?�t����Q=�n��=ym?d��>ف:>�╾H���3�>�0?+�%?}1��򽏿7����=	ɽ?;�?��4?����5<��
����?Ź?d��>R�j��s�����?�8?}��>���`���a���>��R?��^��x>ؗ�>`6�>���? ��ռ����T���&?>�n�;�P
�8PU��m0��$�=y�>�l;>��p���{����>B��ܻN��H���� ��\!�<�}?ߌ�MV>�ai>�L>��(�3 ��k���Ӎ���L?r��?�=S?¨8?Z\��?V�3���l�=輦>��>#ǯ=���KО>C��>����Hr�C����?��?��?�EZ?�6m�I�57����־��žHV���G��J>WG��� >[���	=�Ɔ=��
>U��>���=��>1br>�m=�>��t����+�;��cz��3��5
����nD��(ʾ�^�����7���O��*���jD��]�<���I�8� 8+����?V��>���>g"�>
�̼F��=A��t������N1}����"�� � ������/9`��3$��v˾���ؒ���O�>V�ν� >��>s��<0~�=xUi>���>>�{=�>�ƺ>
�>�>��=��>"��=S#�>�1���n�����%�N@��5��=Du?%�¾����aQ2�GN�u5��S��>��5?�B?B�����������(�>����:i��ً�<؉=��U>��M>�L>N<ɼ-S>_0;h���|*4=��i>~�>�)k:|h��⊾�]�>�8�>��6?�=oq�> t?w�?��?��; y�>zax���=��=��>�j�>��>E�>��$?��F?/�*?�=lZ��&>;H	�=�mȽbi5���Q�#��=܉�wz�=��]=��:Z���^���;j���=tG �n{=F��=���>q��>�:? �>�����I�=�f����l?>W�=�a�a>w�>��>�>o�>� �>�4�.���{��g��>(�Y>Z�b��ڍ�{ͫ��f�>�nC?�?Y�r?Mr�>_=l��O�g�p��<k֓>Fg?�>(�����������ο�W+�I&�A_��
i��#}:L�?�4x<&�hj3��<��l�<VKL>��K>�O>��S>���=��=��>(k>���=y4=l\(=���=������=p�<�xϼ՛������r
J�0���9�q�x���M��%�a��2�<<,?f�?�H=���kw���
� C�=���>�>�>�v\?�_?|p�>��$�&��:�{�Y�W��>U?��s?�EE�O|2��#h>.�<�tu<�s`="�>��)���M�`�����:=��->��?~%2?���= M��c��$��W�2D�>"
�=�d)����?��q?o�������XH��\��L�G.B�*���?0�6gu������}�侣/����=G>�j�>�S�?�&��x��=�U���씿�z����Ӿi�Ϻ�W;����>��>�Xi�;�}����G⓾�{�M૽��>��F=���>��	?��!?W=a?�?��?�E뽹H�>�v<���>R�>���><��>gZ�>�s>�%D>��[�.Zս\��r��~�<�k�:��=t9>]`=�t� ��V����1$=aG��?�v=��<�
�=��=�= >\9>�4?ؤ�>��>Jb�;�g��W��e�m>+�>���>����gQ�w\���&�9�Y�>��*?�8?���Є�@���P��z�U>7�?�`+?��>n��<'��i$��N��1���u>�Dq=���������ɾ���<�>d>u�>���1+�=p[�?m�+?�6?�𽞠��^�Ia᾿O����@>l�?�?ˁ�LK0���k�߀g���p?����1�o�N�]>�8
=��>#�>�X>�>ୣ��Q���	��f�S��;�<�e�=���>S�?1tx>{��t��5���3F?Ԛ��Ž�$W����ľ�AU��s=>u�_>�Y?���r�:ѥ�q 9���>r��?��?�0]? J���xJ/>�">~ >�2=�O�]�-������&>�"�=3�m�Az��3&<}F>�h>Cr�G���]{޾�]���ȿ[�aH�=	㸾�B����QؾUe��௾��"Z���(�ۈ�m��9���m�3���s=�Mi�'��
�?b�H?��J�ñf��"�9~(��*�I�=s"����*��~��������eWp���O<�򬾟����ܶ��������>`���F��K���>���>����I?ȣ�w�6��[.��!���"�>[B�>6i��̀�p���XC�uށ?g?��׾<����%q�j��>K3? hq>�\>�B�=�+�����>��
?��m?��/>&�s������u�?9.�?Zd1?F3�E�(�?���ی>qJf?�?�>�S>�]�=!��c���t��>���?��0?�Խ¢��fD���:?]�|?g�񽔑�>�M?�'�>�^���w�I��wҾ�������t����j>S�,��υ�
��=}��>�f�>��?�m#J�A��>�@� O���H������9*�<C?j��$6>/i>8>��(�Z��Dˉ�$��L?䕱?}�S?`l8?�V��l����C��=I��>b٬>"֯=J���ޞ>)��>�j辝ur�����?_G�?7��?WZ?��m��6���7z�"�׾�r�=���(=\v9��`�=���=��;�@.=���=�\>�	>�[>�qJ>L�%=��>ׄ�S�1��פ�����(�^���F�-�Hj��N2�q񽋡꾉T��{J|�"�!��H���'��i�g@��GA��tǾ ��>�� ?-�!?�J?��z>�&|>W��̢�������k�Ek�B^ �f�	����-=�}p���:�L���⍽�K�jXB?=�m=H9�=t��>u�T=s���W>^�|;K| <\�&>^H>7�+>�q=Ǯ>�n>!-�=A3<5��>�xm�W+���z��6E�\5P9����>�����}�47�h�ھ����hM>��?攜>U>���9��N�1�F��>���ׄe�I��m7>�d�>���>�N�>&�Z�����%�������9�=���>��">&�V���V�޲s���)>�i�>������.<��K>`?gqk?0o?ڹ>���>��{>��>{�<A�=��>_~u>�i?*�?�4?p�>���<�{.�Na={.�=��,�B"��V���d��}R<�Kk=�1��b�=�3R=�&���l"=r�=�wϻ�]���?</}? 5�>��?��>*.�(A��0U��"��˭��I̬�KS?ǔ@?�?��>_��=�]��g*=����&P��~�>��)��c�������>�?T�>�Zr?��]>���ٌ�1T�@)K���=q��>v"�>�v�=Aj�>'�����lӿ�$�~�!����_��Nt�;��<�p�M�M�8y�-�Կ����<z�\>E�>�p>YE>�>y;3>�W�>�GG>�Ą=/�=�)�;CD;��E�	�M=K��!G<R�P�N����&Ƽl�������I���>�v:��:ټ��?ô?L+�cGʽ�S��������K�?�?ƻ8?$Č>C�b���E�٬i�<�ξ٥�=\�=Cp?7S?�g~��C=�R�����f�>G��>cL�7���#���Y�ξ�k����>�0?�?D-�r�V��)]�[o���y�>��=b�<���?/,Y?L�Ҿ�>˾�8X��HX�Q߾}Ɖ<޳�;�:�=��'=�)�.��پ��g�����ٽkm�>��?\�=��=}�����SΥ���Ӿ+�'>�x]>�a?��?6:�3�����޾�l��\����)��>�!���L?/��>Ɖ=?#*$?��2?�?|�>��-?���>�:>Qc���N=Jٽ�`>)�^>�nܽ���>�ޑ>q�P��~ƽ+��=�+�=3�>Pn�=�H�=!b��C?.=ؒ
�g�j=v	u=,�=X3�<�]!<ʞ���0;]��<�bk�M?���>ݮн.wϽh�̽���?�>L3�>��>ڄ�=i⃾�]�a�|�E��>�6?�P"?]�
�*��W�B���Ѿ,�>�>�6?jc/>'��{��<�t��8P���>4*>�����౾��\�žz�>�?i#>��=C߈>�\V?�<Q?�1?�����H��r�ơ@����� ���?���>rtf>Sh�#�L��mY�	�%��=R���F���4�o�S<>�oL>�x�=Q��=���<�갼A���f���=���=.��>�w�>C%?�V;>@G�;���W����G??R����Ǿ�޾ ��4Uܽ���>�.Y>�ͅ�vw?��v�9���v\���P����>W��?]+�?��?G�L�A�%�V>���>���=�꼪���{;3v�=?�>���>��[���ڽ@e��6��=K�$>�C��������'�b�;�ο�9���
���°���:�Z\p���ܾ�x�����o�<�V��U<��[�.
�;�����<�?<�@��v��f�?�?c?[l������L	��T���#��a�<�n��L��?��ڰM�����_���/R�К�����<Ҿ ����N�>��ھ����F��oY��A�>��=�@?F���3��33����#�1>՚�>QIB�;r���Ӂ�u4껴�F?]�?�1��{ݾHF���]�>(��>E��>���>�>�uܾ\t>�L?�b?t�=���&����^<<Xγ?9x?�J5?�侖�뾺���xP>�]?�m�>�>��־Q�E�=�;�v��>v�D?Y0?���������Z9����>d�#=/a���!�>"�>1��>�{�7�R���=Ĥ��;�=�t�>�I���WM�8ˑ�{.ڽ;�R=6�?Ĥ=V�������>��.�,뒿Q}��z߾�7=���G�>_��h�v���>���=�.��t������!E<�J?(�? �J?=?����>�tB>�Xw>��>�pd>oU��괜>��R?�����|�bB�:YE?P��?!�@�}�?�G��WBֿ��������\̥��6>���=L�=3��$�=�ⱼ�(h=u+�=KK'>zi�>��>�~>pBQ>wo�=���=�̆��#�����߮��E3>��P�И��xf�Q������^ƾ�ܨ��A����{��X�E�������V9�Bsl>I��>h�>g��>�1�=��>x��ڇ�~�l�������a�՛�xB����<�[�=�+�������I��X#��)?<��=ē�>J��>S�L����>P?mR,>��g>u�>b�>�>��y>�T�>��8>W�g>�L��yz>W�=j��y"���z:���S�7��;|D?��_�"�����3���߾�ꩾ�#�>��?l[Q>N�'��政�Ux����>�g6���d���ӽ�b&���>���>�= ���9��7z��#콽��=�9�>">���������5��=Ww�>7�޾Z>��>7�-?gp?8�)?[��=��>��}>��>$�=bJb>��s>��>n?��6?�*?���>�(�=�vi�J��<a)B=�Z�R���((� 21�\o�<c]�=L3=�NQ=ɪ�=]�:�;)�=j|�=���:�<]==��>F*@?�5?�m�>�{���#�<�F���.=aCm>]Ҋ��N�>if�>b��>h��>f��>��7=�2����،��`��>О�=F-��@W�����1�>6>�K3?H_?(�>9�4�uei��%�>:6?(m�>A�!?���>61�>c�b=���'6߿��'��U�:A#���\�����R��=�W!>*b�=����7� <	>�Ƽ>@�?�Q�>)M>j�>A'
��X�>�V4>z�
���=ۻ�<C熻*ӽ��=��ּ��Q>���Atc���~��٤����Me<��ҼX)x=�ō=�i?%~?�CJ���g����L������1�>]8�>��>	�>�l�;O��� X���B�[�%�b��>�-W?�g�>�ou����=�_��x���@��>'�>?�i>\ȅ�\����������Y�>�?>r�>�wW�;�`���y�n��1w�>o6�=^�9�?~Pv?5�%�l���&;ݾ `{�E�0�$��>~��
`S�.���+�>�<��?���J���5��Ad���>�8�?�X��=^e�l쉿�r6������=�+���}-?|"�>m�ξ�ڽY���Ⱦ)�1�˾���R?���=V��+?��/?L��?�>�M�$�}>��p?�0�>�?�g??=� ?X�?�j?H?!ߞ>P+c��;��ͽ�ؗ�m����������=c�&>{�5<XG��aQ�I�=��4>��~<y_>&'Z=��j=��=!�>R�=�(?o�"?l��D�o�H�=kZw�U�K���۽��b>�޼���ܾ:彘�><g?�`?��>&�{�����ƾј��uL=��*?{`4?d2�>-7ֽ)iZ�c���X�c�l�j=.�I>6�:����������(Q@�b�g>6N>����e�>(�d?�Q?F1@?���`�p�9��*��Bd�$������>���>�����c��=��3��&Y����.��Ù><.�%9�=��/>��<胄>h��=3iQ=�j>$��dm+�)���4^f��>S�X>W�>��>\��^ٺ��̥� L?i��'�U��Zb������սR��>e�>����?,=>� ���ѓ�W����C>�,�?J�?�[�?I�ɾǼ��қ>��?�
�>�z��&̾��y�HL���x=�V�>�|���Ǿ�}��v�>"5�<�Q�%���P�h[�䦮���V��G� ���ud�����u����>�]���=���\�ӾpB�������8�����
k�H���v���3�?4h�?]V>��<�oqL��/��U�co>�c��˿�i�¾J�L�GY��̐쾃f�U�J��M�M�P���ľf�{>1�m=*x������m4�ֵ����>*�*?��྄�Ⱦ�4)��m���'�>�$S;/ (�E%��z���]�>x?�O?���U�O�־��->Hf?���>,�h�fz��Ž����-+?��[?�,=] ����U���]R�?�r�?�Y?Pס>��!�GZ�1�< 0�?�dR?�$���ּ7��O ����>/f�?ں9?4�
�oh{�Y}��B
?w��?A`o��"\=�c�>�J�>��>9/^������-׾��	�B�H�C�b�ý�H��^o��=�>C�(>ĩ\>�U��"松G��>�ʢ������oO�jۭ���=\T�<�.?ԫ���8=A�Q>�S�>*j˾c���&+;���4<�.Q?��?2f?({=? ���侂��<7Ɵ=��N>���>�y>{�s��

>���>���ڏ��r&���??n��?��?=~?/��KϿ�]������HB��#�3>+t�=q�Z>^�w�u5�=`�>���>���>���>h��>vE�>�_>�>Yrp=�^��8!��ߤ����g�D����40�I}���V������5���о���9������AϽ�V�<�`��q	�����-6=� ?e��>���>�=���>M^������	��p��5`׾��5�t(�����p߸��`ͽ�Cɾ��������c?��s���>M��>g�<(WF>6[�>�w�=&�>�{�>�
U>7��>��>��>��!>���=
%�=5*�=�c=Ӄ���τ��]4���i��]:��:?��|��㡾e`/�������?�h>�?�W5>/W6��9���Hz���>�,Y=�������¼�ۜ>c!�>g!>3l����A��������=��q>o��=���aQ���Q���k>s�?�P��O�=�?z��D+?~1�?9/?��hm�>�=@>/dy>_�`>v��>3��>;��>w�?�Y3?m*?�v?v��=�����=YU>�ļ���=S�7�7����(��>=���7�཈��=��>ӻ>7/ƽ�ѽ�jx�
��=XC?�z&?%-�>g�
?����h�����->&Ĕ>Z��>�'?!">*9�>�?Ҁ>cR>�[��q���{����w�>�s>�]m������[�?�>HFj���n?&�f?��ý�p�=�$z> �=`>�>j�@?�e?�wN>��@=V���iӿ�$�i�!�\�����z��;��<��[N�5���I�-�d&���
�<�|\>�*�>�p>��D>�a>�2>e_�>ӃG>®�=1��=RE�;��;��E���M=bO���F<�bP��5��)�Ǽ����_?��hlJ���?���G�ؼ�%?d�?Y���"��Fξ��Ⱦ���>,?I, ?ѓ�>�?=u0>g�ʾ�@=���9�,;�S��>�`B?�1 ?�V��Z�=Sf1��l��(?=h?�+p>�����P�����Uz��E�>Z%?�ȷ>0��+�D��M������>� �<�jo�W�?m�`?<���9)�8�8��j�ⷯ��"���>E�$`۾lb�
�8�F������h���vE�y��>�Ϲ?r���v^_>�Ͼ%6���ꂿc���"�8>�����?���>O#��Z���v/���	������כ�>�>��>�(?8�?��?�
?�6�>�?e�Zw?w>�1>�u\>�?�#?�\�>�O>+�>�>Ӻ�>��ƹE�����}=�����>�V>Ol�<#��=g>.�=@�>U8C�܎��\4�=3�=k�<=/X�=�(J>���=�7??�a�K�e�߇ =�z��%�=��=���>\���S�� 5���>�7?�� ?U�>�f�<�ᾴs����HȬ=�/?k&'?��>�ܽ�߬<Ȕ���$��0��<W��>追������
�q������șj>�qz>'|н�{,>U>\?%�\?�pk?`�	��Z��+�p�m�*�=�½�?d�?�r��LI���y�v{��ӭY�AI������n��|�PN���B�>�un=+��<.�>�T =�	V�)3)>_$��!��?�o�>���>��>!y'����_	���g-?����2/�N^���"�&���?>�x�>-(ݾ�>��uN��?����v�*�7?���?b�?���?����r��0>��?��o>���l��n���ֽ�=�k�=�����
�����A>�Y�;��Sm �0h3�'����ƿ�f���Y��ͮ���.c������־]��7��#�����oܴ�	�ʽ���8�	>;�\:�n�������c �~�{?b̈?]�U;�6ý�7�_�����#7������ �j����䉾~�Ǿ0���I5���)��C���2��9���=Eo�PK��pW��['�*y=���>�J"?�#ݾʜ��m���0����>?�R<Ǿ�Q��lӟ���ý��]?0YH?�����p񬼇&#>�(.?C
�>���=޷��~�0Jv>�fA?dRL?LԽ]���I+h���
>,��?I�?��T?L�L��d2��1��@oK=�n4?�?�/>qE�;��b�B��؂�>�X?��?��þ@?q�f��L��>Ƀ�?.Aw�)ߨ=@?��>�|ӽԾ�M��+�D�	�׽��>;#���Y���.�⩢����=�t>M�=sL������>��.�,뒿Q}��z߾�7=���G�>_��h�v���>���=�.��t������!E<�J?(�? �J?=?����>�tB>�Xw>��>�pd>oU��괜>��R?�����|�bB�:YE?P��?!�@�}�?�G��WBֿ��������\̥��6>���=L�=3��$�=�ⱼ�(h=u+�=KK'>zi�>��>�~>pBQ>wo�=���=�̆��#�����߮��E3>��P�И��xf�Q������^ƾ�ܨ��A����{��X�E�������V9�Bsl>I��>h�>g��>�1�=��>x��ڇ�~�l�������a�՛�xB����<�[�=�+�������I��X#��)?<��=ē�>J��>S�L����>P?mR,>��g>u�>b�>�>��y>�T�>��8>W�g>�L��yz>W�=j��y"���z:���S�7��;|D?��_�"�����3���߾�ꩾ�#�>��?l[Q>N�'��政�Ux����>�g6���d���ӽ�b&���>���>�= ���9��7z��#콽��=�9�>">���������5��=Ww�>7�޾Z>��>7�-?gp?8�)?[��=��>��}>��>$�=bJb>��s>��>n?��6?�*?���>�(�=�vi�J��<a)B=�Z�R���((� 21�\o�<c]�=L3=�NQ=ɪ�=]�:�;)�=j|�=���:�<]==��>F*@?�5?�m�>�{���#�<�F���.=aCm>]Ҋ��N�>if�>b��>h��>f��>��7=�2����،��`��>О�=F-��@W�����1�>6>�K3?H_?(�>9�4�uei��%�>:6?(m�>A�!?���>61�>c�b=���'6߿��'��U�:A#���\�����R��=�W!>*b�=����7� <	>�Ƽ>@�?�Q�>)M>j�>A'
��X�>�V4>z�
���=ۻ�<C熻*ӽ��=��ּ��Q>���Atc���~��٤����Me<��ҼX)x=�ō=�i?%~?�CJ���g����L������1�>]8�>��>	�>�l�;O��� X���B�[�%�b��>�-W?�g�>�ou����=�_��x���@��>'�>?�i>\ȅ�\����������Y�>�?>r�>�wW�;�`���y�n��1w�>o6�=^�9�?~Pv?5�%�l���&;ݾ `{�E�0�$��>~��
`S�.���+�>�<��?���J���5��Ad���>�8�?�X��=^e�l쉿�r6������=�+���}-?|"�>m�ξ�ڽY���Ⱦ)�1�˾���R?���=V��+?��/?L��?�>�M�$�}>��p?�0�>�?�g??=� ?X�?�j?H?!ߞ>P+c��;��ͽ�ؗ�m����������=c�&>{�5<XG��aQ�I�=��4>��~<y_>&'Z=��j=��=!�>R�=�(?o�"?l��D�o�H�=kZw�U�K���۽��b>�޼���ܾ:彘�><g?�`?��>&�{�����ƾј��uL=��*?{`4?d2�>-7ֽ)iZ�c���X�c�l�j=.�I>6�:����������(Q@�b�g>6N>����e�>(�d?�Q?F1@?���`�p�9��*��Bd�$������>���>�����c��=��3��&Y����.��Ù><.�%9�=��/>��<胄>h��=3iQ=�j>$��dm+�)���4^f��>S�X>W�>��>\��^ٺ��̥� L?i��'�U��Zb������սR��>e�>����?,=>� ���ѓ�W����C>�,�?J�?�[�?I�ɾǼ��қ>��?�
�>�z��&̾��y�HL���x=�V�>�|���Ǿ�}��v�>"5�<�Q�%���P�h[�䦮���V��G� ���ud�����u����>�]���=���\�ӾpB�������8�����
k�H���v���3�?4h�?]V>��<�oqL��/��U�co>�c��˿�i�¾J�L�GY��̐쾃f�U�J��M�M�P���ľf�{>1�m=*x������m4�ֵ����>*�*?��྄�Ⱦ�4)��m���'�>�$S;/ (�E%��z���]�>x?�O?���U�O�־��->Hf?���>,�h�fz��Ž����-+?��[?�,=] ����U���]R�?�r�?�Y?Pס>��!�GZ�1�< 0�?�dR?�$���ּ7��O ����>/f�?ں9?4�
�oh{�Y}��B
?w��?A`o��"\=�c�>�J�>��>9/^������-׾��	�B�H�C�b�ý�H��^o��=�>C�(>ĩ\>�U��"松��?�/.�����aSS�����>��<>K��>,w��[Ii���>ZU?���Q���PG��Đ[��9Q?��?��w?SF'?������y=�S>��=m|>Jt�>��þ~cG>d�>��m�/n��n���,?�`�?�U�?2'{?�T����w���R��y������=U큺��d=v���B�=O�<=�Ѯ<�s<d�&>�|�> ��>h�>���>I%�>��=�\��9�#�j��1���Ǔ>����z��ќ�����#�O��_����䭾WJ�����<I\��潩R��EZ���Z�5>���>�q�>�[�>�1 >f�8>���=^a�3�G���T���B���b�  ���5�����_!Z��Z��;O�F��qe�>f�l=�\�=��>H��=v���ۖ>��V>!��>��>��7=e#�>,�>��y>Unv>9>�};>F*�<-�<>��d�d���S��|��)!>��8?T(��}N̾�ob�-�dpG�>E9>
�
?buA>R<=����Ɇ��?�,�=K�����ľ�Z�z>���>:��>�1�=EQ0��愾�<Q��:���=��<Z�����>2��:t�>*��>xg���=1B�>��3?!�r?Q�,?�f>���>�nE>"؄>5�'>�qH>�UT>Ϣ>+?�\A?��,?���>E��=S	��.�=�l=��I�&��T��KnG�^qI�/s�<�M��X�.=;4�=՗J=d��=�yn=g�;<C咼G>�<5?3�7?���>*q�>������B�}%(��DO�Y�S>�|>��> {>c��>8��>A<�>�=]V �!����㔾 ��>�p>�;Z��Y���|	����>���=��-?r�\?r>�==$��>ES�>�	�>��'>�?=�>�ۏ>a�<,Y�Rlܿ(��J/���w�Yߓ�\��<��(��½;�'9~�s�������=.g�>���>�s�>�>D*X>;��=�q?2c�>C�j��/�6�+�Ѻ��T�>=��=YP���<s�=U?��� =/A���ν�u�<W���6N��Φ;k?�?���׽׾�8оj���,?���=)�"?�>*��=L���n�^�T�;yG��+�>/�j?o�>qI�����=��=4)o���B?�u?���O佐e��p��w�{u^>�J�>�	?bﵾ��N��n�Vc�D>t��=����ߋ?Ħ�?K��"l����� L��R��֓�.ZL=��p��8�W��|�7����c��K����=y��>��?v�轓|]�0!1�zɑ���r��Y��À>=P�=Q�G?_��=�\۾������.������=q�?�ɐ<�ϼ�iE+?n�7?�f�?���>�~z>k*t>k�L?m�>X=?�
?�N ?��?]�Y?�1H?�?��y=��ؾ�ݽ�ƾ�UC�8I<��>D2,>��=�S�=/�c=}xC��d+��/Z<���=;">946>�O=?�=��[>���=U�	?|
?�p�=�["=oZ�=�S��s�ё�ǭY>?<a�ھ }�K�.>��?�?΄>0�;I\�$sҾ���� <l�?��3?��>������"N�5*u�����r�>��o;�bԾ�N �iMd�Jȍ=��a>T�>e�K�/�>^Ft?x�d?#x ?��h��"�������G���e��1��>�H˽۴ ��rq� z�����i�����N�r�>�<<�|`����<Tr�=l�>�<ͥx>�K{=�d�=���=�}?����p�>��=3?'��>�#>p����	�R?�fZ���C��s��Ƥ��%�j��>���>�ʚ���>WN<>��g�����z��@�>^��?;��?���?S�B��UH��C.>� ?)�>�c(��ߩ�M��<��W�@!T<ݾ�>�h�����|p$>{=�{1>aq�?7־8�
�����K���G���%���߾Q\��n��^\���d��>¾��(i��������.d�C{@='3��1cX����I��?b��?��>�=��Q����žV䂽�t��3󸽄cƾ��$%\��Dؾ9�t0�U�Q�$v��J1�di>���=
k��h"���R�Ǚ�<I��>H?�Ջ��?�^��`�k���>aC�;���8��㷒�
�@�\�t?�EK?#x��1�9�p;�g�
>�+R?���>4�@�����;W��(�>uk?�� ?���`���w�]�X>"��?2��?(�V?vOX>LQ1�ڪd����ތ?�Y�>~�󾣚�=�j��h�rd>S��?:�)?ɫ(�#������?��?�{�U��=?��>
g�=�WF����[%���),�kA�����VI���1�����n>0yE>�:>Ƃ���P��Ba�>���}���#u�ś.��7>����(�>X�C2�<��B>b�>��-��)@���6e���\?f	�?��k?�.?;�Ӿ������>���=���=�K?��>(�l���>��/?������7�:�j�5?�	�?,`@��?����Vڿ�̚��8�� !߾Y >k�=�0!>|�9�:t�=�8q=GÅ��RD�a;_>��>"f�>�!t>`r>�&'>��
8�/��4� ��?�����H9��� ��� � )��� ⧾�B���׾�x߾A�ż��:�ⴴ�[�I���K�^u��~���b>���>gS�>��>H�=���=���w-��>�a���Q�+�h��R�rO�We�z������~��������'5?R'ս���=~a�>'�^�[&>o�>��=�A�>B!�>���ȿ�>�Q�>��`>��T>�>�O>3~g>��=!n��NU��_A�����>�� u=?|��#���+4��M޾W��� �Z>u�?��7>�1�������u��#�>�S<�#l��d��-���>���>�{�=�s��t[!�[�o�v�?��=y�k>��0=�|9�.���:���=3-�>�o�P�>�ǖ>�-?�Ts?�E5?��=B�>6��>��>�z*>[�j>Q�v>w�>�Y?�,6?rA(?�n�>��=A�q�[+'�.��<j�R���9��Y<�A��<ͺ-��=��H���=��>9��=��=E��=�e<�}+<���<�Q ?�
6?��>�>������a��p���Q>�\w=A�	�VO?��L>��>b��>?o�>l:��[�ً�������l�>>:�>�m��q��u����=:p�>#\W?�*@?�?>K˽<�>��>Ga�>D8�>�f�>���>c��>���=J�	�^�ѿ���e���=[�H�k|��d��wD>�_2>&�5�ƻ��W��=��>N�>��>[P>��v=�>�P�>�<D>��<B�<ݾ�vbӽ��[�n���X����=r���Qa=tkW�=K�<T����°��M��@�;-�?6�?Bj��)�ӗ��Q������s�>�n�>a �>���>F�<�)�=a���J�Ւ=��e�>n�\?6��>1z�8C�=)�.=��J����>:��>�a>(ڽ����Ծ��>�
?�h�>5)h��b�(�w��/��@�>��=�� ��?��Q?�?���ƾ�.��TD���M�_4r�ǞŻ�_��e$��b3��3[��1��q���!����h=�>���?aܽ�O=E���i��3|e�R���c�=�_����>g^�=2�������Q(�),�9��TT��9�>\�>u6��Z�:?$=R?��?��
?3�?;�ݽ�ML?W�?��?��f?��?_??92P?�1:?�m�>�G	��Ե�t����Rz�4�95ػ'��=P�)>���=z͹<;��<�G�=�I�=��O��a5<�87=2G >�!�=�Y=��>;�<8>?�N+?�M�;��=�FF=�SE���4=get>�6=>�@��o��0w��9 g>��>�	?���>+�%��~�y媾{- ��Ő=�1H?,(?}S?����������=»��W>�	�<���d���d3��];P}�>@)F>�!0<�ہ>��?([?	�>�M��>"/�U�\mk��'L�ٵ ����=WZ���������xP�;�q�Y���T?m��髽����5�E��=�x�=��>>Zӏ=R�:�$*V>?s�= '#=΋Z=�d����>s}�>�B?Q�>�	�<�0*��:˾Q?3�PX�&3��O�:�^3j�d�>箽>��	�,6?ؠ)>�$b�]������Ci?>�\�?S�?�q�?as����F��=,B,?^��>w�N<b��g�~4�ֺ�<ژ1>�A �����N>��l>+���VX�����?US�"!K������/��I���ھQT#��⿾\ҽ��˾\�L������ a��
�>�s�>��\�O8�����뾾uj�?�f�?��=Y�ҽ�%=�%�K�Ӿ2ԡ=�ؾ��;Z�ɾTe��D��?�5>�r2.��k�0 2��mȾTN�>��F>t��������_p�_����>�?����ur��h��vl��Vt>����H-��{��@���+�?� ;?�k���n���+�k>� �?�X�>V��Ά>1>����?#?�'e?��a>�ʖ�4'�����>�?��?
�]?9��>��a���h��/W��)j?��??�o�>אP<��ӽ3��?�c�?�j?�P�-���Qk4�F�?7C�?Q#���<=P�>&?+@=�7�m={�<��ʾ�	���7�����;�k�[�����>9��>���=�i߾�־|��>�׾��J��p"�=�޾>�2�J2�=���>*e�*r��ft)>O�^>��+�tՉ�A"���2=�mW?�ҷ?�m?��?�T����o�:S���{���>/�>g�a�o�a?i�>������,���>"��?��@,I?�A���տ��:}��]����>���=Sgj>���c��=~��=p�i=��<{kB>��>��S>b�k>%[�>�UA>�2%>���;p'�86������0�;�����l�g�r��^�ھӬڽu�y������ >�F$ͽ��&@����>~W���=� 0?��?|�>~	>@�>�<����,R<�E%�h�ƾ3��W�0���jT���e�����!�����\�YX�>1����,>O)�>w˔��#?=��><�=�h�=9�=r��=t�>< �=z��=�5��Q�=b��;̧�=a�>������.���;>���d=?��F��V>o29�F5��9��$>'q?�6�=L&��=ƒ�㝏��l?��?���ǾU�޽�<d>	?�[�>������=�k��?ھԟ��~�s>��>�:�濿�¯~� ¾"h=�/�>�Ӿ�(�=�<u>��&?�v?+�7?r�=n�>�R>�֑>-��=
qR>�V>�>:h?�]7?51?���>�={p\�6�=X�A=~@���T�6��el�������<e�A���:=�6�=x.)<<�V=r%`=%���B>��<Q?&�4?I��>�Z�>�T�
U5���,>lL�>
�T�:�?:�>�M�>ܠ
?tF�>/q���������Kz��[�>vա��͇�����Q�g>	??��?��T?�j�>`o}�xU��׍���*ϼ|��>�YD?�g0?�0e>\^�<� ��A��0�ڿ����tn�H}�=ͩ�=#
>�-��Y�|��'s=�O����=s��>��D>nh�= o�>?�?.I>��}��>�v�>���;�}���-�=��;cQ��Z�=���=��=�K`�[q%�O�߽y_z�D�;�2=\Љ<���<B|2���?f�?�[%>%>�ɷ��1��_v�JZ\>G�>�/�>��>\�>.��9`�5�\���Ⱦ�@�>'O?d?���G�<AK޽{>(�B~?{+�>�I@<�0V>�n<x��c*>�2?}y?��>� Y���_�é�������>���=���H�??�?$��=��Z���2Wt��{���;=c�x�h!�ć"�>!A���b�[��-.���t��q2>d�>�g�?ǚ����1���:��sh�*�z����>*�L=iOS?��	=Զ���Xl�l�����^"��e��>�m�>��=��>7�$?��#?��J?4�?��?w�%�F�>	�<Ѻ�>p��>.�?L?�?m��>n`>B)H��Դ�9�!�܋��b�5=n���	��=�>>R,>M /�aь=��<1 �Q��4+��4T�;ppR;+�:c�A=� >���=u?��L?�5�=m:[> f���b��(>�>ߘ�>�ZA>Nɾ���>E����?޼j?��p?�L?N���4��Ӷ"������>=�?ډC?���=�	���!|���*���ƾ:9�>7��h�<w2�Q��ڭ��.�z��>�=��@��̆>�z?k�M?F�?�Rw���L���}�"�����>#��;Fq�>`?�V>�k��*.��9����b�K��Qy�<߬A��$x<��>v;�=��>�+�=)->|��=�	�_I����X�B흻U|�> W�>�*�>��M>���<>��LO;W�C?��x�������P� ��}]��ks>�hC�,�����?�6���zs�:6��$A`�,�#>��?��?�?ӂ���J�K5>�M�>�Ț>��;�R���6�YI����
>�C>9�̾�����I�Zg�����>*�7�ݡ׾}X	��[,�!T���-��m�)C	�SX>�#����^���+��u����=�Ҿ����W���SE�7;=1��W��r�}�x����	�?n�?ôʼ�=5�:B&����Y(���{>��C����=W�;�T�n2�9���}��������MQ(���
��L�>z秾�"��:w�Q��<��>�[N<C�?9���b_ ���'���=:+>A�ӽL��:y��䋿�D��۠S?r�/?
"�v���1>Vd�>q@d>L��>�Y�>
�M��S� ?�>?l	?���%���x2��SD��)��?���?o4F?��4�@�1���Ѡ=��>���>*:-?yW2�ͼ$�v�>g�>�)?���>-��w�t�}K���?�c?��$��J�>V��><R�>-���4.��l�>"D+�zig�KF����=Ud���当qۼ>I>7��>a�>C�¼xp��|��>�׾��J��p"�=�޾>�2�J2�=���>*e�*r��ft)>O�^>��+�tՉ�A"���2=�mW?�ҷ?�m?��?�T����o�:S���{���>/�>g�a�o�a?i�>������,���>"��?��@,I?�A���տ��:}��]����>���=Sgj>���c��=~��=p�i=��<{kB>��>��S>b�k>%[�>�UA>�2%>���;p'�86������0�;�����l�g�r��^�ھӬڽu�y������ >�F$ͽ��&@����>~W���=� 0?��?|�>~	>@�>�<����,R<�E%�h�ƾ3��W�0���jT���e�����!�����\�YX�>1����,>O)�>w˔��#?=��><�=�h�=9�=r��=t�>< �=z��=�5��Q�=b��;̧�=a�>������.���;>���d=?��F��V>o29�F5��9��$>'q?�6�=L&��=ƒ�㝏��l?��?���ǾU�޽�<d>	?�[�>������=�k��?ھԟ��~�s>��>�:�濿�¯~� ¾"h=�/�>�Ӿ�(�=�<u>��&?�v?+�7?r�=n�>�R>�֑>-��=
qR>�V>�>:h?�]7?51?���>�={p\�6�=X�A=~@���T�6��el�������<e�A���:=�6�=x.)<<�V=r%`=%���B>��<Q?&�4?I��>�Z�>�T�
U5���,>lL�>
�T�:�?:�>�M�>ܠ
?tF�>/q���������Kz��[�>vա��͇�����Q�g>	??��?��T?�j�>`o}�xU��׍���*ϼ|��>�YD?�g0?�0e>\^�<� ��A��0�ڿ����tn�H}�=ͩ�=#
>�-��Y�|��'s=�O����=s��>��D>nh�= o�>?�?.I>��}��>�v�>���;�}���-�=��;cQ��Z�=���=��=�K`�[q%�O�߽y_z�D�;�2=\Љ<���<B|2���?f�?�[%>%>�ɷ��1��_v�JZ\>G�>�/�>��>\�>.��9`�5�\���Ⱦ�@�>'O?d?���G�<AK޽{>(�B~?{+�>�I@<�0V>�n<x��c*>�2?}y?��>� Y���_�é�������>���=���H�??�?$��=��Z���2Wt��{���;=c�x�h!�ć"�>!A���b�[��-.���t��q2>d�>�g�?ǚ����1���:��sh�*�z����>*�L=iOS?��	=Զ���Xl�l�����^"��e��>�m�>��=��>7�$?��#?��J?4�?��?w�%�F�>	�<Ѻ�>p��>.�?L?�?m��>n`>B)H��Դ�9�!�܋��b�5=n���	��=�>>R,>M /�aь=��<1 �Q��4+��4T�;ppR;+�:c�A=� >���=u?��L?�5�=m:[> f���b��(>�>ߘ�>�ZA>Nɾ���>E����?޼j?��p?�L?N���4��Ӷ"������>=�?ډC?���=�	���!|���*���ƾ:9�>7��h�<w2�Q��ڭ��.�z��>�=��@��̆>�z?k�M?F�?�Rw���L���}�"�����>#��;Fq�>`?�V>�k��*.��9����b�K��Qy�<߬A��$x<��>v;�=��>�+�=)->|��=�	�_I����X�B흻U|�> W�>�*�>��M>���<>��LO;W�C?��x�������P� ��}]��ks>�hC�,�����?�6���zs�:6��$A`�,�#>��?��?�?ӂ���J�K5>�M�>�Ț>��;�R���6�YI����
>�C>9�̾�����I�Zg�����>*�7�ݡ׾}X	��[,�!T���-��m�)C	�SX>�#����^���+��u����=�Ҿ����W���SE�7;=1��W��r�}�x����	�?n�?ôʼ�=5�:B&����Y(���{>��C����=W�;�T�n2�9���}��������MQ(���
��L�>z秾�"��:w�Q��<��>�[N<C�?9���b_ ���'���=:+>A�ӽL��:y��䋿�D��۠S?r�/?
"�v���1>Vd�>q@d>L��>�Y�>
�M��S� ?�>?l	?���%���x2��SD��)��?���?o4F?��4�@�1���Ѡ=��>���>*:-?yW2�ͼ$�v�>g�>�)?���>-��w�t�}K���?�c?��$��J�>V��><R�>-���4.��l�>"D+�zig�KF����=Ud���当qۼ>I>7��>a�>C�¼xp�����>"��]�G�3x?���	���E�#�<1��>�� ��%>�>U>Ch>3�)���������7����H?k��?�X?V�+?��徤�Ծ@8Z��{r=Uh>G��>�у=��Z[�>&�>#뾻�z��^��~?&h�?��?O?��n�l%ҿ���͊��t���U>�=�]>�"���=���=��J����|{>��>Y��>BI�>E��>U�$>��>���XD(�n᯿a��tC��6�W��S�� ��-^�4�0~˾����"bȽ�D���&��x�{4�oS�r₾8^�=�?L��>p>�b=
`>�I���*ؾ�G��-�F�1������پ�<�IQ�LU��R���>���꾍�?�o"= �->��>�����<�
?�>�z�= �ʼt��=Ǚ>5�>X�>�'�=h[�=ܦ�<[�:��N>����b���9B����>L�r�&�>F0F��>�QF����òξ�>,�>�>������)*���?���q��'Ի���>�H�>�$�>�u���� >�x뽤�Ѿ��5=��>n
)>l���n{w�8���Xl¾�l<�>�>��Ҿ�7�=p�w>߬'?��u?B6?#��=}�>��[>�>�=�Q>�YW>���>��?��9?��0?�z�>~��=��b��	=4 7==��N�����sڼ�����<�3$��sN=��=Y<�;o=��G="ۧ�8]�;��=�h	?�j+?g��>&�>VA���GI�F�X���<P�>�]Y=�?P�>Ĝ<>M'�>W >�Խz���rk�"������>A��<	.��� ��#�>�@E>���=�7?q] ?���X�n����=�>�s?^�'?mz;?K]�>味��ar�h���տæ$���
�f9�;���g�<謾�ֱ=�v>�B������}�	Z>�Ҫ>i��>�S�>W׼=Z>�V�>o�Y>H�<㫰:�����=ݒ?��E��%��<v��=�s;��ݽ�/6�^�:�p�<7�l��(��=�������?��>+Z=#�=���5(� Z��<��>/j�>�c>x:?��n>w E��T��'4��ξ�'U>��i?���>R�O�Ȯ=Z�)h!��@�>[ܠ>6?ʆ�=�䐾D	���L��?̓�>�L�>(�,��7��]��3ž�P>�0~=�(��|�?Z�?/;A���㾼w�8Bj�����=�H=�Ki���ξ��;���N���D���!s�}�M>K�>��?�W���<(�4��$c�g�s?�<o�>h�#?L���N�aGV�%=�����,�eB/>W�>������
?R�B?A�?~�A?P�?�s@?�-ӽ�>�/�ܶ�>��S=I�$?�B4?.@7?�?U�?��%>0�O�0ꂾڢ���>��r���3*:>��9=ɖ=>^o��]�7>[,>(">k�M=���{�|:�ڋ����=k��=�R1>��
?�2?�v=G7>�m�H�P��8	��|�>;d>m=V=2�>�m��G6!?��L?�>b?U�%?o='>�1��,�B("�ˎ�>��?�Z?mG>���=.�9��������W��մ6>4���G��־�]@����l��=B��>�U��?r�>m[?��1?VN?GHv��C+���i� ��:�#>P�<M�>"�>B.��c;�]55��r��;O�����Q(��o#��M�����=Yͽ<n> {/>��D>}%{=�k=�D�<+�����;<�>V��>l�>?n�>�O>g�Ⱦ��پ��I?�ʡ����^��M.Ѿ�1���>H�<>��u?w4�}�+$���>�\a�>v��?jr�?�8d?"9A������\>#X>�h>�X-<�!@�/��ꈽ�4>�Z�=��z�� ��'6;s�V>bx>��Ž"�ʾ��侌�R��ȿw�2��}���#�B<v�A]��
۾�r��d<X�2�>}����ﾝ���!�ｘ�0>�]t�ܫ�;>7���ܾ���?��?�)Խ"¾.��[�]�ҝ��|>h�ɾ}7<��Hɾ��_�f+s�J �)�����徐�ľ�����
�+%�>����u]��:R����>�$=�T�>��ھ�'���c^�&(>2I6>�J6�|������=���.߾ޕU?VK?�[]�r�o���	>�/d>�R�>���>b��>�k�:�PR9>�"x?ͮ&?:�׽��|�#���}��)��?v��?~QT?n?�C�+����M�=�" ?;.?}�?�	>��';��{���})?��?�1(>J�Zk��7 �:)O?�]�?lC1��9�>��#?�>Z'�_x��=��H�>,���%�>E.�=rؾ���x����!=n��>�_�>QYb�~��A�>5����?D�	5�����oU���<���>��
rp=�1b>�
T=|*�kY���G��_Y���>?��?�xT?}�?�I��pT��(j9��M�	l>?B�>��]���x�>}��>�y��^l��8�n�?��?#��?�I?�mt�RGӿ ��0������Y��=%�=�>>��޽ʭ=ԗK=I̘��Z=���>m��>o>�;x>��T>��<>y�.>^���p�#��ʤ�5ْ��[B�� ���Fvg��{	��y�����ȴ����������Г���G�m���T>�K�o�-7� #?w>?�>�B��oj>5X��a��N�=s��F����7$�� L�dg��y,��h����żu�ד�h�?혞=�5�>�.�>yt��d>su?H��=��=�.�>�;�=.�P=r�>Tkz>�r�=gq������$��B��>�i��}��������j�>1ѾOo�>�0[���~>7?E�Ï>��L^�@9�=3
�>;GA>N�S���-׆��"?�H�����W L=�xp>���>���>�Y���C=`�=�勾�P>�@>.L�>��N=Q/���J�pz���@"�T��>�/Ծ�O�=��}>;(?�t?��4?u�=H�>�a>\(�>F�=�G>ѻK> �>'�?lL9?�O.?W��>�Ϸ=�b`�ZM=kD=��=���X�@�����������<����-X=X$i=�F;x>\=X�G=X7¼ �:'=۝?i�,?<�>���>�WX�\=���!�H�>W#�>�/Ⱥ��0?8K�>C~v>��?<�>wzP>��w�R�ˀ�:f�>�>��\�<Y��<f(=�ݢ>�-?	s?E�>�>�r���.���;=<0�>6@D?�?���=}Th>53�1����ٿ{9"��<�8��:�[м��={��#�J��9<��"�r`����%=�NH>�ڀ>�k�>m�d>�|�=��.>�K�>�\V>�=�\=�-���=7�f�a�A=��W�����F^v����<)���ò��:�_=0��r��}���w�?m��>`)�=��M�/���X,�AՓ�I>���>�n�>��?��>�!+�oG��!J�����N�>�W[?�<?���[���w���WW���>�s�>�2�<��>>Pۛ���C����>���>���>H� ?<>njC�k�����ؾ��'>?��=��P��}�?v-i?�o ��ʾK>־G�f������=߁��=Ou��4SK�qjO��r׾Q���� Z��p<>T�?L��?�;�P�������~�[�c�ƾ��=~il�f�I?b�={B���2
3�n�������>)�>5n(�/=�>cH?��%?��x??N��>: ���>Ģ�<���>�,>m{�>O��>�k?�X�>�L�>���п��M��i��3)@�D�T�{�(=� >��q>��=7�N>�s�<�W ��@��9�=���C�����O��<�TX>��>��>��E?��>z2b>#ja��lP��aT>��>\WŽU!� ��;�1�o83?=5Y?�xP?��?���>�%Ѿ��0��:H�sj>Y?x`P?�ޫ>A�$>n����{�r׼f=�&>t=�=pm��������� C�U2�>���=)�y=l�y>{?v?c_<?H�:?rJR���0���������`%>�4��\?Zv�>����Z���e�,��o�|�N����S�<
B���P={�=�;
>��1>���=��>>��=u�I�/�ʼ�<�=x�;�NX>��>M�>h��>�� >�*;s���>I?M��|��b�����־{DL�0�>M�->�=���?S�>�}�Mp��01@����>,�?���?B�f?R<� y��]>R�c>>��Q<[�;�I��p��ܺ9>�\�=�怾�����:+�G>	V�>/߰���Ⱦ!q�2�O���ӿ\-1����w�]�������ؾ���m�<�|��p�ؾ�<��Y������۽Y��0?Ͻܚƾ�ż�Q��?���?xH{���þMG�7K���j@��?�>�y���=/����JϾ�b��:5;�����{�گ���������Y�>��������l���;<��>��=��>����4�̋1�:��>�>��⽕)�Pk�@,��1���e�`?M�:?��1��]b�ZxT= ��=��>�ݿ>^�>����}��/&�>�pH?���>�>޽�q�����Ί���F�?�X�?�P?�̷���	�l���	�I��>|"?�)?�n���Q��^>��>���>p��>��a���w�u�e��(F?�[?�F��Y�\>���>7�d>�����&�`�=���&˽�?->Bb��H���'>���q{�Wb�>*��>�%������,�>���?�?��3����%�X�2Θ<���>���>u->j4W>�=��0��������9��BB?
�?\�\?z"?��ؾw���2׭�0�:;C��>���>�����?ͽ���>���>j�k��0�H�?���?z�?p:K?�M|�a�ֿ�ɡ���������T��=�ɤ=JcP>���,�>��=��P=G)�Xy=���>D^p>��>�z�>b>,�>�Q��f,������㕿H�u��	���C�(��5G������¾Rؾt����Iʡ��3���Խ�{f���ڽ-/:=�5C?
v?*���u=���>`�Z���J��H������kA�@9��b��I8�J�~������XR�<I~�W���:��>Vu=X�=�/�>�l�=Ӆ�= ��>=
G=qJ=�O�>{C1>��>��>)��=̆�=��F=����G>ܞ�=q��鯩�$���s�?j����7�>��۾��K>1�e��3$��Wy�P��>��?p�=�Ӿ-�������R�9?,8���׾�M<&���=�>�>�<T>B>2�оޚ����a��!>�Vd=�~��aҽ1�ž�������>Xm��{�!>���>l�?l5g?��4?8[�=��>H�>��V>�>(v�>s�}>��>�#?Oj;?1�1?��>"�g=J�|���F:V7����+�ss��s��<��6�<b{�T~e=Ԏ�=��j��I��q�N篽���<��=��?<�0?�ҥ>�2�>s�H�z-�7SL�.K��o�>����$�>w;�>��?�<�>k>��=|ɽѮ˾���HZ�>�H=O�i�o���+v>U�>�N>��9?�=?|&?=4!#�G`�=$�>ʋ�>e#?���>���>	=��L����4�>;��þ�P͉����q����>�>�`R���U���n�4�O>*�>�}�>��?\��>�3�<n��>ڍ>�~.��ԃ:b�>�h�=Li��u��@伕6=c���νSϽ=T�ȽΔ
=v���3�[��b3;'p
=Tr"?�?� �<��<�þ"�/�B������>|�?��3>�V�>�t�>u(��3s^�Ɛj�����)�7>x�%?c�?��_���������eo?��>U�6>��V=> �<�G��[]$>�X�>�f?�?��㽑W��q�h���>�7P>�yM��j�?���?��c�Ğ�t���Y�U��í��=��Q���C��Qվ�U��j��,����پ��j�rڸ>��>pߩ?�XY�1r3�G	�� ��r��9<H��=��#�J��>D��=�4 ��������>�wk�=���=�ܑ>�Ⱦ(��>��!?��?�,l?ƴ�>+<_?�Yb�C�>TiE�E�>���>��>�s ?j�;?�H>?+A?x}G>:���lJ=�����=(�`�὏�9>uf>'�z>�c��~�=7�+>q�l>yP�=jvk�����/�=�7>`"�=;)����=���>rgG?�/>�Dy>��-����0���@�>��;�oPQ�%�Խ�Z���~?��"?� ?��>%A"=x��~,��2�R��>�'?h{4?T4�=�����v��3T�up�"�<ǽ���Y���⿾���Wl>д�>�J��:�>2dt?�w2? x!?�_��;�*� s�79��P��=:)����>��>��$��K��y�|�`�V��D�<=�3��	���Լ��s�u'D>^�)>�0:>��)=��B���;P^ =""�P�>>yn�>I��>�R�>C��=�ڜ��۾�I?�X��NH�HQ����Ծ��9�Ξ>�.>\����?����'~�Ȧ���?�%a�>b5�?��?�c?��=��	�@�]>��^>�>�G<o-8�G�c���д4>`��=�Nz�V��|aq�y�T>�F}>Œ��jɾ_I��Hs�����.�5����7��)_=\+���	��XL����Z��>������Bà�_����H�=�rg=�{\=q�S�����3�?9�?���='j��R���{�v;"���+=U$��~���������f�jy����Ūƾ��+�=�:��Y���>������li�&�V��H�>��=�E?���AH���|4�j.=��>�Z��&���&���8��k۞��B?ؕ1?[������ye>��+>�P�> �)?խ�>��߾z�	��+?|�?$��>�e>x��A����愽.f�?
��?f_?�n�M�,����,��<�r�>��?��Q?�฾G�Ͼ��>�#?Ti?�j�>�-�UM�¿
?ʌ?_�i��4U>��?��>�����!����g]��Q؉��A�>ўZ=���L#�'jc�0ʥ>�S�>��>C�ｴ������>.ِ���y%��!龁���,��]/�>�̲��31>s��=]><��9��.���タ��u�`q?���?:,?y�:?�A�,7�����D=#�h��>Ν�>�j�>�5j��O�>���>e��	Y`��)���?�J�?��?�`V?K�R�T7ȿ����Q����9y>.ӗ>��y>��=dM]>���=�ԫ��=j�>M>�As>>��>�_>�$>pc�=
G}��u �����2����!�^̾����� ���x�*�uI����}�[:������U��.�U�
D?���ɽ����We>��>R�5=m?���>`��f���c����Q����/\�19���h�5�=�@�u��V���@���֚<2�ƾ�k?�!s>�d9=$���
��wQM>���>��l5�=7>ź�=�v=��0��*j>�I�>�� ?��)>��W>��{=�R���������<�=ט��N�>��r�LQƾ1�9���A���S>��
?�>��&�����eS�?��>[�8�-��Y=�\�=h��>}��>7�O=f;����A���Խ�>�L�>b$<0�q�F�c��� ��};���>�ݾ:�=ߕs>��?�q?h8<?Q��=W��>�>e�}>xؒ=2�R>��}>���>de?*�1?-�)?� �>RT�=I�a�g�y=:=�W��x���R���`�l�s����<�PL�|�=O?�=Y<��F=� y;���IL�<؟Q=V(�>�9?U�>���>K���uA��eQ����t$>��?��j�>c��>���>��>A��>t�+>�v�.����� ��>\%9>"]���r�Goc���i>b�e>�P?-F1?w>��e�5��;ٲ�=Ο>�G?�b1?r;�>[�#>��	����ڿ�Y���&�r,->3��>�FH���O�;��=nj>pzo�@@P��%�>&9�>-��>j�>g;v>Z�@;B��<���>Kߎ>$>�+�<m����[�=�N<a�m]���KQ�<�W ����y=�M�,�$�oRo<7���< ."?��?�<ɼ�==i#ҾGB ��5��L!?b�>6PD?��P?�Mm>���M1c��o��4���>U�?\�?.l��q<�����Z�>�T�>�<Og켚k���1Ⱦ��=�T?��?Uv�>Z�.�o�r��ݑ�))쾍ָ>�`�=jܷ��]�?��a?t��u�����߾>S���ݾox��y���H�+���X��� ���"�ѿ�T<�^��j*>S� ?��?tľ�k�=���ۭ��Pp��̣�VA>(��><' ?
�>w�ž�f���%��m۾^�F=��>���>C��=���>��(?�A"?2g^?:��>?��/�j��>䖭=���>�N�>.?�?d��>�cw>ԕB>�[��k$��(�P������=���<�ل=i�C>|�Q>L�Q;��=M�=E�ڼ��rk�!٪<4)�;;<c�c�=m�=�>\Z?��>UbD=<E�=���;-�)�)�>�bG>�-��I��Z@��
������>�+?�t/?�?HԎ;t��8h��,-���>��"?�;? 3?�*��J�C�޽�Έ��f>J�>���N�ľ�o0��!���,�%�<���3�\���e>��z?��B?0�\?O˝��e[�I�C���1� <�� > �I?H}Z?Zg>��Ⱦ��'��]�SU�z.��H��T`v��-�=*Q2>uHO>D�>��=eq=cp��l�>ٽ������=��>PL�>+�>'��>��<>x鞾>��7V\?��Ⱦ1-��Tp���:��������>.��>	��>xK>����E�����7�پ��.?ǀ�?���?��U?��=��=^*�� ��&1�=_U���>\>V�>9�=8��>]r��<��`��E��=U�'?��9?@�!>M|��ݾ���>Ȑ��.���E˽}=��$�U����皾�t��\,��{�=}����C�Fq�c?B�b�N����Ģ��ԾB���ˌ�?Y�?Vi�=���t� ��Ӡ��y��iP<j�
� �g��ʧ���$4
�Р��]�r���Y@�"m�a�>��`� ���\H|�I=+���V�A�I>��-?8y���̻�����R=5k#>BR=!澈F�������K��KX?��8?�+뾴'���$ὄ�>�
?���>��>*����޽���>��2?C0?�㣼�W��^���Zmq�Md�?��?��M?�Ƙ��h>�6���7�����>3G0?,g�>��q�
�ӾA��i�>��<?�?Y�T�=uI�fP��߽�>'�z?��Q��|�>�?�L�>?�=ˇ˾-��m��������>>J-<N�G��A%=���ߠ<^�>P�>�}���_M��+�>�<�=�A��A6�*����+�e����k�>���r�}>̎/=~P�=t-��l���Q������tyW?���?h�S?��N?A����$���=Z)��<6?A��>XU��{f>��?�<?��K�edp��*ƾ��?���?t3�?�%U?x"���;ѿ�!����������>Sq�=Y�Y>ru��� >�Ӏ=\���sP�kc1>���>�Lf>�l>B�d>��%>U7'>L���4%�0C������J�>������y�d�3{=�e���e��������M�&����� �.��1���u�+m��]��1��>G�>>&�>�ď>��3>�kA��V:�)�׾�
��p*��W� H��l�� 8�D�p�����۬�;�� ��>���=���=��>5M �0$�=G��>s=B1>|�>�Y�h|�����A�Zl�=��>��>aA�=b�{��^��f��������
>��>��w?�k��ch���LE��
򿾉��>�K?`35>[�������\\���>#�ق��$>��=�>��?\�\>����!��3˾ܗ��z�>�]�>��#=�޴��z�bZ̽Ա��{�>]�׾il�=,Ox>�(?�av?�i6?��=���>�_>�ڎ>�7�=M�J>��O>��>��?�8?6�0?wQ�>,f�=��`�.�=8�<=�B�ȝZ�2ﴽ���PY!��͚<��8�r3I=m�s=���;p�[=�x>=M��^��;��='�>�;?��>Z��>N�;�^E��[T���߅>�PY�.�>C��>�}?\��>W�>P�!>����_ľ,�Z�>��S>��[��#�D��<���>��$>��<?L} ?G�3L~��w=�U)>i�>��?�(?k�>�|�=� �����jӿ�$���!�ż������;��<���M�s����-������<�\>��>�up>�D>��>Q-3>�Q�>LFG>�ۄ=<�=8٧;x;&F��~M=���+G<T�P�����0Ƽ������o�I�7�>�u,���ؼH�3?v}?r=����>\� y7�wV�<�G?�ȥ>�1P?S�1?P��=��t����U��������>��?�ů>�H�	i�=}�=��>ܩ�>�zO>e%μ���<}�D��U���%_>'?[�?w��>��콮EU�XD}���L�>��=1+Z�?ޠ?�eX?.��4�����-�6�vo�>��<`@R��u�J�-������Ӿ�6���6���=�Z�>�٢?����9�=�$�����C�s�&c�{��=�e>@E�>u��;�	f��K����&�i���M�D=�Ձ>�=�>�~�#?�>�n7?��&?k��?�:?�:?~��n24?s�=��8?8?. -?: ?��>��>o0�>Ę������/�j�@����y?��@��<�۝>���>���=͞9>��L�#=�ƽK�+����m���g=��=S�0>8ی>?�B�>W��=AS�=�e�n����R=�p��Y���G��5���r|?X?��9?r��>�]=-ؾ�ғ��a*��aJ>.�8?�?8�?�$_='�>=~�;9A[��=@�)>dU�X���K&�����W#�IF.>�>�I���8�>��i?�!C?��X?���:�f��$Q�ʔJ�Va=,�=�%?�F#?���=9=���R&��T���A��2�PI������q�=| ��w"�ݒ�>��:><$G��2��'t�<0���B��E�:*K�>��>?���>�,�=�پʞ��d?2����I������r��2�=/>l�:>Q^�=;I�>35�g����=��%�2�b?o��?�N�?PY?׍�4�1=��u�&M��?��=Q�H=����������>>�7�RN��6����⾣W��|?#�,?��}=:�Y�+�E��=8�ο�T>��O���o2�A�)���`�}� �����UU��k=����Ê��}���n��/Ž⨘�����پA	�iz�?�7�?9Z>�䷾��������-'���=�������EܾV>�����x��#�ʾe��C�.���M�
��dE�>aI�����av���߾��=��U<��"?����ݚ���31�6h�=��0>�?=�ܾ@���r��������f?1�&?_M1�nS���l[����Z�=N�	?��b>a����M��y
F>KTc?�vM?�D��/�v��/|��G%�� �?��?)�A?�e��;��S�	rj��W�>J?r��> A��I� �&����>J�Q?�F�>:��L�b�Eh�Q��>B��?��=���>��?���>��?���U���,��8�O��>%�ƺ���)q����F�����>Jk�>3����Q�;�>�~R������$��f����1{�<�.?�ʾ�>��>��ڻ$L5��u����r�C��;cc?���?��@?��D?� ��C��k�������q>vA�>.��>z
�=�d�>%@�>qS*���i�Ⲿ�H9?�s�?l��?�rj?��M�)pĿ�E���j������a�=C?�>%�_>��ͽ���=�	��-�=B�>I�e>K�>�s>4�">0�O>�.>|����}�á%�ˌ���N��fB���۾����첾;Ѿ�N�� �����̞����uQ�ȳ�R�1��]��������k8>���>��=M�@?:�*>'I���I�����2��m
���ʾ����H�۾du��4���z�z�¾�H��1ȼ�:��a"?�/�>��=�%.>	�=V�}>���>]G��b:o>�+�>�6�=ό=o�=K�}>;?`>uN�>&3�=Ϋ�>sF�<�쇿�W������ܬ=�+ڹ�';?�:�k���)-�b�y����>�:?#r�>a�?���u� �솼>.d��"=���7�<��=�>���>��=ݠi��R,�Y$A���|�GC�>��?��=*-q��S�������=n;�>�<־�0�=�v>��(?�w?`16?�ݟ=�}�>?*^>i��>�|�=�XM>�_Q>���>��?d�8?v0?nC�>�K�=��^�lK=�T==�|A���]�;8��_����(��n�<Q3�J�K=Tu=��<�U\=��<=�ӵ�}<-�=&8�>�9?��>pm�>=t�oED��OI����M�>�zu�j��>~Z�>vt�>��>� �>`:>��|����,�վM��>w�D>��`�Gs�w�2���g>��P>��L?#�-?�"o�>��H�<�n�=!��>�0?l�+?:�>�@%>]}�� ���M�zO������[z�E��>�J<W'Ͼ�gw>[�E=���a,���<>>�>�Ƃ>�(I=c=9>��=�z\�k�>�1x>f,_��o~�N���K�����<�h�<9�<�>�v���m�����]�v���g�-�+��#<�k�<��<>ee�>�4?��U>ñ5>z���=K��6��$�?�8?��?��(?m�<��C���\�@�I�;r��Vp?��?gv�>*�����=G���,.B>i��>A�=���=��2�(��������=S��>q��>%ks>��6�ǯ@�%\��n&�T�W>�Z�=fŽd�?)�]?lL�ͼ5�9�վ��)�pI
�o+�=1���.�N̝�cf$�\�g˽�~���VJ�Y�>I��>��?sj�]�=��D���I+q�ঢ়���>-:�>��>
��=~Ȭ��۾��X���ʀ>Ɋ�>���>�oP=���>Q�<?N�?�Bm?hO?�>tƶ����>C�^>3�?�d	?;?��?a��>�.>%(>���΁�v��OO���BG>�!�=ӳ=�{�>G�>���=c@T=�)K<�Ӄ��N2��v�t(<� /=4�o=�{�<{�>ۭK>��?�i�>��e<�j#�	Cڽ�-1���>}�=��ef*�E~���-A�;(�>Z�
?��"?���>g*�JB����R��!>x��>�_?l?�_�A{T=����$���=� p=I䔾�Y���D��wþ�� ����=�5=�:����#>7?�.?���>"5�>pQ;���r���1�%�=R>D^? �6?��(=!���2�_�f��+����gnd�7U̽(ש<�a<H���@d>9e�>�=�������p<�=8=>+[?��>:��>ǽ[>���=�ߴ��_[?�7�6�\����3��W<_��>��?nuB>�$�>c	O����MӘ�X�"��i?�\�?�B�?k*I?Wn�&�=�ԉ�����(���e�=ц>Zx���6���r�>����A�MM��B�=� �>&�%?
,>��X�O�_=n���#=��!F�> �����Y�������?��4�߽$7�=�ӾLI��s\���޽b��Pu���Me�,L�Ծ��\#�?y�?�O&>�,�|�̾u�
�r�?�� >�����q>�8
�hG��L�Ͼ�r��g����)��>4�[M��������> �k��%����y��*"��>S��>R@7?�o��q	�8����_��H�>�7q>8SX�\�c�����@�@��}p?8�(?��վ}弾nS�����<l�>	�>���=j����-�"C>��8?O?��>�9��9˔����n̰?c�?�U?'�z���*����j9
?�<4?�N�>T��P����R�1��>:x�? �J?��H�UU>�?��>�u?�ׁ�b�B>�P?��>���� ��9,����
{���ۄ>�t��3��>����	��d�2��=T>A>黪���־���>��P>a�҉�矨��@%>�͠�)��>1�]��á>���Q>�m&����Dw��>I���!;?�s�?�P?%�O?ѯ���
�j�;�fNl<�S?�ޖ>�?$>p�� �^>c��>���ߣ<�g����/?,�?k��?�P2?���EVܿl秿d��m�����T>4�=��Y>$��6#>��<�x��x�=��>�a�>��E>�6>k>���=XX�=e���M!������o��E04�G�����ޗ�~L�.�/����������w���;����Q��[�۽02i�-� ��o���<��9?R5�>�x�>D�>�.>�m���'E�E澀���z0�T������vYL���6�n���ʾ��h�-�'�X�?�H�=�#�d��>y���Bu���m>�(]>p4�=#6F>[G�=G��=���="�'>� =>��>��=}�>ǋ�<�Ȃ�k;y���J��g�d�=�B?�K�@��7��������Lu�>�?���>�%!�@���%gf��J�>����l,�J�����A<�e>���>p*k={弽�z��L���C����M>>�3>���]̖�t�0��o>���>�վt��=�p|>��'?�u?q6?6��=���>َ[>*��>A��=:�I>�EN>#c�>�0?��9??�1?X��>+�=��^�_�=Q:=73;���V������u��S��~�<�.�n�V=��j=Q�	<��[=D�<=���i`T;1�=�U? �$?9�>,��>�����@�z.�w�:=ˌ{�w���y>B\>>�F�>C��>��>��>f�=K�k�l���>^��>����Rs�9��=K�>�3>�K�?�[?���>R�v��=%7?�>{ڻ>�??o?���>P�{�2�
�"�ܿ�qe��7C��tw>ۯ�>�D�=����?���#>�ݽm2��T�=���>t��>7�3>�,�=@�ۼE��<�j ?��:>)%��"<Q�.>�H�=�ý.��=�O�����=���b��ol���q=�{<���3��6�ݼ���=O�?��?b��=���>#�˾�)�(+����.?]�>^�=�� ?������Gb�W�5��ؽ��?x^d?B��>�>^��R�=}�><�>�?�>�m>�X�w4��S��x���*q<r/�>��E?XG2>g�@���U�X�i��4����>�=Ց��.��?�%j?�j�l8��9�8a3�HK�T`������*q���������6��]�p.A�C��=R� ?z�?E�m��_)=M��t*���䋿��<��l>uy�>�? <�>�C��㏾�&�d2_�Tv��"g<�b֗>�^��@�>&]�>�-?O?���>)-?�;�x?�a>\`I?��-?
X?U?*�/>��(���^�!U�<�,�����G߽�V*��'=YA>��>�й<��=쨽y0�����!�$���+=!�Q<�0�ў=���>xob>d[?�4�>,u�=���;�/�0|_����>�>g)���Л���]���/>"�>?]�m?�X(?O�=l�k֑������>�)?��>�a/?ɦ�=����۾L��;c����=��=�U�u&�i����틜==��=��i����>j҆?қ9?��'?�+�=�-9����.�#�Nʪ>��?��'?�G=?<�?[Ӽ� �A���sd�e\��'Ǽ�$������Yv=L8B=_��>'O�>8��>������������=��x=]6�>5��>���>�`:>+�=�h��y�'��Wd?�v����$��R��U�*����=�!�>�2
?�>t�B>�F%�}�k�����(���> ? Q�?���?��]?�e��/�B��l=�nQ>j��>A�^��[�-B�>R��<��>�v��ȗ
�#>��v=<j?���>�[7>)3��A�=>�ؽ��Ul��x��Z%���=[�7���޾Ԓ��r���0��K��P]��_�����=_�����;پgp����B���?��?�*�>Q���@2��pJ�L��#�U=`&X�o6���Z�#h��ܾ��v��ۦ�4f�
���x�b�HA>h0��=���J��Z�/fս;��=z�?����+{���"��Dg=r��=���ʵ��B��e�����|?�=?ԃ���оM�7��ޓ�b_�>��>���>+z��˽l9�>K�=?`�?���n����x����=�İ?*B�?��??�O���A������3*?�?5��> ���C�̾�q�?4�9?�>� �2h���;��>�[?�;N��yb>���>]4�>�$�,����7&��.���8��s�9>]u�!���Dh�V+>��ҧ=��>�x>J]�`����}�>ԧa�|���N*�L;ݾ�K����/��9�>8L辧�J=�������?��V��{�i�@��N?냭?�k6?�\?Kz��s�^�!�"�o����?��?���>���=�g�>���>� ���L�y���k'?3�?t��?J9x?6�d�>Gӿ����������=%�=��>>��޽�ɭ=��K=^ɘ��Y=�q�>���>o>A;x>x�T>͛<>��.>q�����#��ʤ�4ْ��[B�� ���wg��{	��y�����ȴ���M�������>Г�x�G�[���T>�<��>���F�+>���=��B?��5��0�l�;�f��ƾ�}#��9��u��	���i��*ξЁ��쾌`ξ�dQ=�񥾮P#?O��=���ݷ ��H�Z%>��>n#�����=O��>��_�lc]��L=?��=h5�>�1�>�7O>_�>��#�lF��}�y��6�NQ�=�+]�!Q?�3q�����B6�%m
�S����i�>@�:?`��>���ˋ�$�)��թ>���I�q�%)�Ya=��=6E�>ߕ<Ps��t����n��� Y��E�>(�?	�=��
��k��9���꓁=��>S�վ�+�=�<x>��'?��v?)%6?���=*1�>E}`>���>�@�=�zJ>��N>���>.?]A:?�2?c/�>�l�=P�^���=��1=%>��Z�$-��PoӼ� ��t�<�'��L=D�o=x�<��[=�XC=�ù��$�;S��<q�>%9:?d�>m�>�
<���E�O�~{�1>nI���>�>7�>�@�>Z$�>�g>��v��_�� 1۾]�>џL>�`�Vt|��j��>��F>�VO?a�-?���C�A���=���=�s�>3C�>~$?��>>L>(j��-_��߿��7��!1���;O|B=J�K<F��UG��,�<)w�	����=S��>^!^>�d>R�.>],�=|��=Vx?E�|>�s�<�0.��#�=W��=~�[�Ĩf�Zvj��YR>ٗ鼺�G�:����]�г	���<ITI<5�=R�?jI??�%>jE�>����9I���;4�?�!?��?q�>?�Z>��0��P��]>�b�'�r�0?���?�>�����p�=簡����:���>Pɇ;ݞv�ة꽡�<����M ���?7��>H�>q�D�R��a��H)�	�>�U=�Z*�D�?nc\? d��V���5�Q�:�3��}􇼊z(��ay����w�(�X�/������ �2VW�)��=�h�>Xo�?�4�KkV=����A�����~�����6s=���=���>�%+>p3\�yĳ�V>�1ّ�ޟ����<>
-�>��L��-�>3c?"��>SF)?��%?�_?�E��x�$?��5>��9?7=?2?��>�>Ú��LQ>e,�e"�=O��iiھQv
���
�R�>JW>c�>��>�~$��hb�C���X���l���<��Z=;���Q�=
��>ah?N"�>z��;ӧ�=?驽O������=0Vu��`z���<�H���-�>�?�?�C$?[�>�c�����}��}�Q���=Q!4?�; ?>�>�� =���=j�|��=}��=P�b>9�����,�w�*�>���N��n7>x�=e�V[�>x�?��*?���>݉�s���}��u���">0��>6"�>n�*?��>����$�4os���C���?���S�����01=[>8y�=]��>�*�>��>``��*�X�����w�ܻ�k�;���>��?D ?X�r>�P>���
�X�V?�sB�̴�����l�(�Z�{>�L�>R?`JK>Ͷ�>:����t������-�"-�>���?��?#�v?򌓾�E>;[�s:ݽ�2=�����0��a�=���>ᴽ>Zg���9>����|=7h�>x?��>�.־�D����<2�ÿ(�8�y����oN��~���X��ED�0兾���a[�=�R��;}A��Y[�?V&�� =�Vܷ�����¾R���D�?x�?�X=vq<�!��'$�I��wN�=�����)�����X��鷹����A��3��&.���-�n��zB�>#꙾H���(�v�a[.����<�)h>99=?�8Ӿ�|������"8��^>m�)>"��M	r�>���
�}�a?5�&?��ݾ��;����Έ=��>գ�>`�p=���`@����i>�>*?z�A?�*d=K�zb��l	�Ty�?�j�?bZ?Ѿ2uH�$�Ӿ�K��O��>fF6?�`�>D������g���\�>�F�?�9@?R��F]-�'��D�>���?�1���^�>�1??Y�>�-�&��=ᏽ��&��`�{:�>jƅ�NH���fF=�ɕ��� ���>��=��$��1�=L�>qR�b����Ɖ��qp>�܈��R�� N;?R���d�Ͼ�V�>��>�FT�9���Z&���MϽO�[?E��?
�_?�<?�	�vf�>�a����=�GҼ9Q�>��?>w�=�z�>�=3?�
��_��������;?�o�?O�@��?�<���!ڿ�G��w@��&t����=�̘=[�'>�񽷗�=$`�=��ڽ�Fƽ��>�9�>��>'f�>J�;>�A>�|�=an���(�9���B����1���G���c8{����m�U����쬾A����~,��{�Wk}��(�ہ��n�$煾���=��>�8>-LF>Y��>�s�=�ܭ�S���[�O�>㊾��#�o�y�i���l�2<јE=��n�Pw���ǽ �
����>m��=pw�����>�0<�R>>�T�>�ug<�d�=�MK>Ai�>7;�>/ >Zq�=/�>(�=I}3>���>+>ou�)�p��&�M�P��Š���I?�Z�D���rD�۫ƾՕ��I�>�?kH�=F~-�E&��sNs����>����eL�w&���μ��w>0G�>�S�=��6<W˴�x���B��U`�=��t>�W>75�<!���#�@�=K-�>��־��=�!V>�V�>��z?5�7?�oƼ
,V>��>͸�>�&�;.�H>"�L>�#�>��?��2?yB!?�R�>A��=�<s���B=9�=yt[�2�e�V��Xf�<�_�<�-<�D��y�91k=���=,d*<C**=P0��-T���ݼa�?l�C?��>'I�>ǅp�q?(�d~S�$>̻Nf>S@f�Cڟ>���>��>M8�>z�H>1��^���Syܾ�B��,�>�?�>���������6>QZ�=�M,>J��?:�?���H����u<�$>c��>Ӱ3?M��>���=��^>��ʽ4��ޜ��>���'��b��=H��>�1�����;�>�H���t>2�?�l�>��>%.f>_�]>'��>�S�>�xZ>�k���C�<]8��>6�;��=��F=��D���m�<�S�=;9;m��dG-��l��<>>�[<!N?�$&?{B/�k=f�&踾�4�x�㾽"�>��J>֧�>�c?7g0=	{�'�r��p�g�m��>�6?Iv�>�A��'V=&���ļ�Z�>��>�� >�4��n���*_���b>P�0?H�5?NH�>mig�c�{�꜉�"���j�>���=E������?R?Vg �<����� �8���cԾ���=������T�ds:�o=l���߾`O��&ͥ����tl�>�?z��y4�>��������� ��G��1��>��S�ܜ�>Q:�>n�߽��þ�`��X)�����}P�@��>�k>�?�!\D?U�9?6��>=_?*K?�%#��?��+?��?v��>�J?��:?���>OC�>���=����"�{>�$���^���YH���ɼr�I=I��=c�>��,:�=Em(>������Mԙ=gn<9��y�B=�!>)>A
�=tB?��:?�,���B�=��>0�&s�&�t>�޿>��R�� 
�Lv��U>5�>U�7?e`�>ǠK��I8�������!?�a�@?^�(?fk�>l=>L�U>�� ��5L�>q�??G��ے��t��h�g��) >zے>Ewq>�>�r�>��V?�Q8?��2?�Y�,X#��臿*����7=�܌��� >���>�V	>"(�P��<��4Sh�?m;��w�;�DM�0W*��j>�g>�#>ذ>���=��b�S��q�����
1���H\>y�k>�a�>���>I >�Q��پ^0?�˽Ib�7d;�I����þ�c>�
?eʾ�>����5���vɿ҉,����>9�?	f�?7̃?lj@�5�k���`>"?n�> �����3���C˕���5�n��>Zؾ���~��=8s�=
g>A�"�9�
�8iG����;����M�K����r[�5�8�}���)s����O�HN?���9���޾I�d� ���k�e6��4�+� �^�J�g������?i��?�A��y��	Ql�v�����F�>^�����5Cؾqb��T��bk&��(���-���C����h����q>"s⽜љ�QĊ������y�^��=��;?�����/���$�?7�=�.9>��_m�� ��\D��Q�?���u?7 c?ռ,����H��t�>5��>��y>-a>"���Lũ���>��P?k�>azX�'A��sՁ����s�?���?M�C?��s��J:�f��i���3�>���>�
?��d�B���!ʾH	?m-?�L�>.�Ⱦ�h����1��ܦ>O� ?�:@�`Rb>G�>C�>���v��!�c�_����2̼�T>����) ��t5���*;�=�,�>�`k>�Ҙ��������>��p�E!��6홿�8n>C������:?m������Bw>�j�>���kÜ��֝��ʦ�"�h?4�?Y� ?}.@?���M��hl=��<��>(�_>�Ѳ>�����9-?X�Z?��+ਿXa����:?�h�?�g@\ē?}���z:ݿo������'�Ǿ���=M��=q��>Yo#���D>t�=E;C=�N�=�ƀ>�3�>D)�>��g>ъ{>�j4>���=x����1�������B�C�3G�,w��]b�Y'���<=�ه��|پ?l��=���Xy<�6����!$��艾��^>%�>ьS>�5n=P�N=�>>}7��@C����*��(%�mS(�� R�w׽�=�1�=�4��֫D�M������E?�6"���>d�?N��<8�=q�>5�=�Z:>��Q>^�	>�4�>�n>΁�>��*>�̌>�5=(UW>z_=N��<\��Cx1��1R�#�{�i�G?i4�����>�%%�r]���g>�?[�J>L�$��D��r�w��`�>W�N��CS����@��-�>w��>��=ԃ޼�k�N}������=vP�>���=Ʒ�����h��6c�=Q�?��۾�E�>}U�>��2>�x?�?�@%>9��>e��>3ŗ>x�1>��~>��>Zz?�-?6�?q�?\ظ>s��=��&�=! =�-���my�����:S� ������j=7	�=HK=�L�=�jj=��j=i%�=��$;�sݽ[��>h�=?9��>N��>Ψ����>0Q��@��%�>�<��@H�>Z"�>Y��>q5�>�1n>����`� .�2ξ�?}_>���K����-h=�>�!>���?s?)KӾ�M]�$� >8SA;�x�>x�?���>��=�WS>��"=M���c� <��$����E�p=�R�>>_��Lll>�=|���Lʾ�xH=$m?>@��>X=�>�"�>�4>�+�>���>�٥>b�>��=�/�=�pS=J<����+>���;�˙�����M<Q�ɽe���y;���̽�.����=0o���>�%?�hݽ��½J����1V�����>�FY>u2�>v^�>|�罰�'��?q��2�^�	��?��X?+��>P;��6[N=z�=�:>�a�>+6�>��w>}7.�`w����5�U	��M�?�?��A>��<�טe��5~��� ��_�>r!�<mԏ���?y�R?�K8��}�� Z�L06������V=��!>ކ��)���5��<j�����s�.�6�_�z;�_?	��?y٥��o>.�	��d������[�O�3>�!�	�#?G��>g�'��G��E�u�q�q����������>���>H� ��b'?�!?���>�BY?g�1?蓼���>���>�R>Iq�>��?�W?��	?�G�><�1>�yҽ���=C	罆>���#�����Uۣ=��=��m>D��<n�R>��=�F����R<�o=�<��?<p2�<���=�Е=F*e=��?m) ?Z��=� >Sd���Ԧ�	�=v t��M+=���Jބ�-_H�ba�>�6 ?�?E��>e���B���ξ������7�8Y?vX?���>?��=�cL�������e�|>�T�=�':���i�0��h��-Y��M�>9o>�=�s)>9�?��E?}/;?�y��o^���a��L���+����=T�>��=��=.�+��a���t�,t��j�;��ԡ-�� 	��+>��>�I�>�>N�>}=y����֪�=��� Yp�$��>���>~	? ��>k�=���ԾY�?��4��V:�9���k��
X��2/����>w�'�Q�>tm�=q��vĿE$Z��r�>]~�?�x�?K�?c�X0G�ҨV>��?٣�>�>��v=�E�=&@��Q̐>�G*>6þR.�#'�>oR�=a�?>��b������I����=a���P�S�"���=/~��`0��z��>s��>�
�+>������g�dh���4�L)1�A-���9��Jf��#��?�ҕ?K��+7��fw׾t�����`(>u�D� ��T��ѽ^���8�������HV�.:Ҿ�s>��N><$��c.���2%�$&����g��ZY?��R��e�a]Z�m��>�9�=xy,�#�*����R���r��]F?a�<?��N�)�֚����?I9y=A�k>�_N>z��-���%�~>ԴC?���>�������p}�G\�<i�?��?�r@?Mf>��_�,���:�=U��=��>�#?�0о����$��J[?�L<?�{�>p+�q����#]��ԟ>~�?g�]�k��=N,�>xn�>�hk�/z�L�>)�վ��I=��z>oW�;����:#t�0/��E�>LO?�>����ۜ��=L�>qR�b����Ɖ��qp>�܈��R�� N;?R���d�Ͼ�V�>��>�FT�9���Z&���MϽO�[?E��?
�_?�<?�	�vf�>�a����=�GҼ9Q�>��?>w�=�z�>�=3?�
��_��������;?�o�?O�@��?�<���!ڿ�G��w@��&t����=�̘=[�'>�񽷗�=$`�=��ڽ�Fƽ��>�9�>��>'f�>J�;>�A>�|�=an���(�9���B����1���G���c8{����m�U����쬾A����~,��{�Wk}��(�ہ��n�$煾���=��>�8>-LF>Y��>�s�=�ܭ�S���[�O�>㊾��#�o�y�i���l�2<јE=��n�Pw���ǽ �
����>m��=pw�����>�0<�R>>�T�>�ug<�d�=�MK>Ai�>7;�>/ >Zq�=/�>(�=I}3>���>+>ou�)�p��&�M�P��Š���I?�Z�D���rD�۫ƾՕ��I�>�?kH�=F~-�E&��sNs����>����eL�w&���μ��w>0G�>�S�=��6<W˴�x���B��U`�=��t>�W>75�<!���#�@�=K-�>��־��=�!V>�V�>��z?5�7?�oƼ
,V>��>͸�>�&�;.�H>"�L>�#�>��?��2?yB!?�R�>A��=�<s���B=9�=yt[�2�e�V��Xf�<�_�<�-<�D��y�91k=���=,d*<C**=P0��-T���ݼa�?l�C?��>'I�>ǅp�q?(�d~S�$>̻Nf>S@f�Cڟ>���>��>M8�>z�H>1��^���Syܾ�B��,�>�?�>���������6>QZ�=�M,>J��?:�?���H����u<�$>c��>Ӱ3?M��>���=��^>��ʽ4��ޜ��>���'��b��=H��>�1�����;�>�H���t>2�?�l�>��>%.f>_�]>'��>�S�>�xZ>�k���C�<]8��>6�;��=��F=��D���m�<�S�=;9;m��dG-��l��<>>�[<!N?�$&?{B/�k=f�&踾�4�x�㾽"�>��J>֧�>�c?7g0=	{�'�r��p�g�m��>�6?Iv�>�A��'V=&���ļ�Z�>��>�� >�4��n���*_���b>P�0?H�5?NH�>mig�c�{�꜉�"���j�>���=E������?R?Vg �<����� �8���cԾ���=������T�ds:�o=l���߾`O��&ͥ����tl�>�?z��y4�>��������� ��G��1��>��S�ܜ�>Q:�>n�߽��þ�`��X)�����}P�@��>�k>�?�!\D?U�9?6��>=_?*K?�%#��?��+?��?v��>�J?��:?���>OC�>���=����"�{>�$���^���YH���ɼr�I=I��=c�>��,:�=Em(>������Mԙ=gn<9��y�B=�!>)>A
�=tB?��:?�,���B�=��>0�&s�&�t>�޿>��R�� 
�Lv��U>5�>U�7?e`�>ǠK��I8�������!?�a�@?^�(?fk�>l=>L�U>�� ��5L�>q�??G��ے��t��h�g��) >zے>Ewq>�>�r�>��V?�Q8?��2?�Y�,X#��臿*����7=�܌��� >���>�V	>"(�P��<��4Sh�?m;��w�;�DM�0W*��j>�g>�#>ذ>���=��b�S��q�����
1���H\>y�k>�a�>���>I >�Q��پ^0?�˽Ib�7d;�I����þ�c>�
?eʾ�>����5���vɿ҉,����>9�?	f�?7̃?lj@�5�k���`>"?n�> �����3���C˕���5�n��>Zؾ���~��=8s�=
g>A�"�9�
�8iG����;����M�K����r[�5�8�}���)s����O�HN?���9���޾I�d� ���k�e6��4�+� �^�J�g������?i��?�A��y��	Ql�v�����F�>^�����5Cؾqb��T��bk&��(���-���C����h����q>"s⽜љ�QĊ������y�^��=��;?�����/���$�?7�=�.9>��_m�� ��\D��Q�?���u?7 c?ռ,����H��t�>5��>��y>-a>"���Lũ���>��P?k�>azX�'A��sՁ����s�?���?M�C?��s��J:�f��i���3�>���>�
?��d�B���!ʾH	?m-?�L�>.�Ⱦ�h����1��ܦ>O� ?�:@�`Rb>G�>C�>���v��!�c�_����2̼�T>����) ��t5���*;�=�,�>�`k>�Ҙ��������>��p�E!��6홿�8n>C������:?m������Bw>�j�>���kÜ��֝��ʦ�"�h?4�?Y� ?}.@?���M��hl=��<��>(�_>�Ѳ>�����9-?X�Z?��+ਿXa����:?�h�?�g@\ē?}���z:ݿo������'�Ǿ���=M��=q��>Yo#���D>t�=E;C=�N�=�ƀ>�3�>D)�>��g>ъ{>�j4>���=x����1�������B�C�3G�,w��]b�Y'���<=�ه��|پ?l��=���Xy<�6����!$��艾��^>%�>ьS>�5n=P�N=�>>}7��@C����*��(%�mS(�� R�w׽�=�1�=�4��֫D�M������E?�6"���>d�?N��<8�=q�>5�=�Z:>��Q>^�	>�4�>�n>΁�>��*>�̌>�5=(UW>z_=N��<\��Cx1��1R�#�{�i�G?i4�����>�%%�r]���g>�?[�J>L�$��D��r�w��`�>W�N��CS����@��-�>w��>��=ԃ޼�k�N}������=vP�>���=Ʒ�����h��6c�=Q�?��۾�E�>}U�>��2>�x?�?�@%>9��>e��>3ŗ>x�1>��~>��>Zz?�-?6�?q�?\ظ>s��=��&�=! =�-���my�����:S� ������j=7	�=HK=�L�=�jj=��j=i%�=��$;�sݽ[��>h�=?9��>N��>Ψ����>0Q��@��%�>�<��@H�>Z"�>Y��>q5�>�1n>����`� .�2ξ�?}_>���K����-h=�>�!>���?s?)KӾ�M]�$� >8SA;�x�>x�?���>��=�WS>��"=M���c� <��$����E�p=�R�>>_��Lll>�=|���Lʾ�xH=$m?>@��>X=�>�"�>�4>�+�>���>�٥>b�>��=�/�=�pS=J<����+>���;�˙�����M<Q�ɽe���y;���̽�.����=0o���>�%?�hݽ��½J����1V�����>�FY>u2�>v^�>|�罰�'��?q��2�^�	��?��X?+��>P;��6[N=z�=�:>�a�>+6�>��w>}7.�`w����5�U	��M�?�?��A>��<�טe��5~��� ��_�>r!�<mԏ���?y�R?�K8��}�� Z�L06������V=��!>ކ��)���5��<j�����s�.�6�_�z;�_?	��?y٥��o>.�	��d������[�O�3>�!�	�#?G��>g�'��G��E�u�q�q����������>���>H� ��b'?�!?���>�BY?g�1?蓼���>���>�R>Iq�>��?�W?��	?�G�><�1>�yҽ���=C	罆>���#�����Uۣ=��=��m>D��<n�R>��=�F����R<�o=�<��?<p2�<���=�Е=F*e=��?m) ?Z��=� >Sd���Ԧ�	�=v t��M+=���Jބ�-_H�ba�>�6 ?�?E��>e���B���ξ������7�8Y?vX?���>?��=�cL�������e�|>�T�=�':���i�0��h��-Y��M�>9o>�=�s)>9�?��E?}/;?�y��o^���a��L���+����=T�>��=��=.�+��a���t�,t��j�;��ԡ-�� 	��+>��>�I�>�>N�>}=y����֪�=��� Yp�$��>���>~	? ��>k�=���ԾY�?��4��V:�9���k��
X��2/����>w�'�Q�>tm�=q��vĿE$Z��r�>]~�?�x�?K�?c�X0G�ҨV>��?٣�>�>��v=�E�=&@��Q̐>�G*>6þR.�#'�>oR�=a�?>��b������I����=a���P�S�"���=/~��`0��z��>s��>�
�+>������g�dh���4�L)1�A-���9��Jf��#��?�ҕ?K��+7��fw׾t�����`(>u�D� ��T��ѽ^���8�������HV�.:Ҿ�s>��N><$��c.���2%�$&����g��ZY?��R��e�a]Z�m��>�9�=xy,�#�*����R���r��]F?a�<?��N�)�֚����?I9y=A�k>�_N>z��-���%�~>ԴC?���>�������p}�G\�<i�?��?�r@?Mf>��_�,���:�=U��=��>�#?�0о����$��J[?�L<?�{�>p+�q����#]��ԟ>~�?g�]�k��=N,�>xn�>�hk�/z�L�>)�վ��I=��z>oW�;����:#t�0/��E�>LO?�>����ۜ��b0+>�x���}��Ss���=y?��">��?��w1�-!;�Y�?�L����Q��ì��"�S?�j�?dd3?��:?�D�����f��C�=@�
>f�>/zE>�w��)�?Q��>=Rо����E��rQ4?�?L1@�'\?�⊿��ٿ�ƫ��ƾ��Ѿ#�=rTr>4b�>�ý�_(> �I=���A8=+4�>�h�>�9>1�y>��:>�6>�mD>e*��e�#�	�ɿe*��`|&�Z�	���	�s��ܘ|���h��\�W��¾�|���)�5�ط4�U�/�G|ӽ�e�L�>N?�V�>�K>�c�>[�>'NӾ�$���q��5��
�Ǿ�)��f"�����f½�\��z��<�.���0!?�}�<��$>AE�>��K>8�<�]i>�3W>�m�>�ɜ>��x>��=㨈=Ll<>ED?>�Z>�P$>D�l>�G�=f����Á�8+7���R�篔;|eD?^V����?�7�S}��8���ۂ>Y�?k�O>�f'��ɓ�x��>��!�q�d��ͽrq�"̃>g޻>��=#���*�#�]n�f�罄ʵ=)�{>RN�=��Ҽ8"�����if�=�e>c���lv>}>{x�>p�o?uW?���p]:>���>UL>�@"�y>}>�T�>�8?DuJ?`.?�>�X�=h�j��.�="��=7����D��.�i�><~D񼧖����,���)>^��<8;*��x�����ѹ����A��y�<��?v+B?��>we ?[ap�fC���`���U�#�>M����$?C ?VQ?�|�>AQ>�5ɽҁ,��.�����z�>�kC>/�a��y���>=y�>�.�=�L[?��b?#�=����=>a�l>u�=f6�>5?��>a�P>���=У	�J㿧�7���/�j��`��=T��=o��>��!��NL�
����r=�ͦ>�ڤ>yn�>��d>`B>	��=���>U{>)^�:3�F<Dq�=$e�۴˽*��=�)<F��RT���b�����&��������\½��J��쌽c,?�7?�Z���'��$�, ޾[M��9?"'?ij?��?7��>m�����`+T�$K˾��>��M?&R?{ؽa�=�Q��HK�u��>��>��=�Т=l�8��g��0���	,�>�0?+U�=�� ��4�U0������>u��=\�#=�ш?O�P?Ȯ�q�̾+B
�7XU���۾f��=FF:>�"�2���+��(�B��j�񸠾 � =�m�>�Z�?��i��R>�ȶ��S�������N���>�<�&?Y�>��e��/ؾ��E�38��Ӿ
�.=��>4@�>bϗ;�S?�:?\
?��N?�4?7�� >���>���>~[�>�(?v��>֦>��`>��=&;0��忽���{K��bJ���>ּ�^�;�E�<�
>孢=v>�>D��=�e�=���=N�=�O�=!m<��r�s`
>�D>��9>�?m�?��D��3�=J�'�i$�?1�</���G"9�%q�	�a���[>�6?(�)?���>m�R<����J��ׁ�z�E=i<?�n'?��>�V�=��>��-�N��vRk=c#j>�#�=v����Ҿz�Ͼ��d���=8l�>��=�Q�>1[x?5M?T"?�P��;<O�iFf�s�������+Jý ��>��>� >��i�]8��Vt�M�x�4$2���������w���2q6=go>Ư�=Hܴ>(�X>���<�M2�W5B�mkN��A.�{��>��?��>���>q[=���x��~�?,���P���0��p���ܱ���F>	t$?�׬�v?����U��3�ǿK百רg?��?�b�??���E��Y*>�s�>LB�> �%��S�=׸�>q����Ur��+>]�E�Ҿ��/>� ?iV�>���<���Lj9����=%ÿ�Z�8��VG����pe�5t8���=��H=x��^� �d�u���E�C��νg˯�����5���(���镕?i��?=�="������-���3�<�6��C���^���ح�wl����
����O&�|�I�g���W��=���ZƘ��'��j��}����=�(?�a��
W'�OI�9��5R�=ľ���}�,3��9뗿g=����=?s&8?���ʉ���6̽���>�3�>_(>���<����L����>E`'?�
�>S!$�.z��;6{���=��?��?��V?Yƫ��+�PM־�V=�.?S�E>�	?νt��^ͱ���%?i�U?���=)��c���G�����>��a?գF�0�F>�<�>��>���%�Nz>Wɾ�B��-��Lb�� �̾;�.E<;:�>D�>s�=�o��� ��>84�n�N��H�������5�<��?k���m>B�h>�>��(�Z���Ή�6���L?���?�gS?�e8?�>��&��A����=�Ϧ>���>���=v��]ƞ>s�>�P�Enr������?%<�?��?^TZ?	rm�Ô࿍쟿�w�����%*>��d=��j>�5�����=y�%=\�1<LY��;D�>T�>��>zy�>���>�>>�>�ހ�1�!�,�����&K�� �F����x���89���� ��g��'jF����=O ����	��S��x����8��SZ=��?��?��=�=M��=W��;-���'>�O���� ��˒��<��x��dmY��������� �ܹ۽�<վ/��>�Y>2��>>f>�ü�
C>�x:>=v7>ԙB>�>��#��>�o	>��>Yyf>�A�=E��>-��>���?��p$����T�]�����>�G?�赾�0c��'<���оd T>�_>&�>.Yb�����i����!�>4�=��*����f��S�>FC?��7�M�=oe<��������u?>�0�=��;�,�=Mʁ����Г=���>��.�h=��">X8?C��?�*2?�k`?��=�*<>�}�>�G�=�{�>OI>Q|(?��?2�@?��>�i�<r�J��У=�����0�va�<��ܽ�Y���Ҽ ��<�Q��r@='�<�&>v���W�>�%�@�'��	�=P.?��?B��>���>�ZR�� �(�"�J��=�!p=kfU��Y�>�Z8>�A�>ģ
?���>�� >!�#��'ƾ�G����>��>X~�������� >~�z>��>��?�X�?��p��&����=��B=���>�E?�8?&�o�2\�>,������fؿ�f��*;���X���*F�<Ǽm0ὼ��;�Ä�G@ҽX��=Q��>���>��p>'��>oQu>�!�>�8�>M�A>}9|=��>�N���c��(��j�=<���x�6=���퍓�.<ӽ���ozv����� �B����[�)�?4�?�`]=��*���j!��v7��x]d>y��>Y��>�,"?�7�>�޾7�b�ɧC�XOz ?y�v?���>4�p�c�=�u�<�|w=��>��>n�>Q�G��`��eĐ��{1=%��>�{)?�l�>��Q�J9��f��
��~��>R�Y=������? �u?3���Q����1��-J����>�v�Ŝ��־_���]G���"����t�?�o�<���>^��?�&ܾ��;��@�z����������:>�]�La<?ZV�>(3������𨸾�\Ⱦ���=�%�>�]黁\
?W�0?���>:�E?h�W?�?�-��k?�?�=v��>4��>�o�>�((?�7?�Ŏ>��>I�>�EV>%KB�]D���P=�v,�p�>'�c>K9>��>��=ym>�4���C�q�j%-=�>6<<���~>,&�=�v�>��+?�T�>-v���o��.K> �f>�Y;���>*�P���]>�>
��>D�?ū?8?����_�ƾ
��=y^/?J�=?�s�>�TJ<���̾�澠EC=���>ܕ�>�!p��&�y(ľ>ﾾ}?��>*z�=�4�>q�?ǡ>ŗ?��
??4K�����wq��Lw>2B���!?���>K}�>~fE��K5�7d��0Yk�VV�0�>r��,��x>��`>F�6<P�>.�D>�\�>��}�a��iؽ.b��ŏ>&e�>�?��$>u >/ֽ�-����cJ?�8����������վ��H!7>C�G>�����>wr��A[��k��$$9��>:��?ȸ�?qjU?p?R�l���_>x�a>��>��	<�i0��N�`X��'�!>��>� �� ����Vc=��[>(�r>$���eϾ��޾R���Ӯ�^_�z�F�b��"o�����r���>N��~�_>V���jl���侐�����Y=���vRٽ��#�Mrоo?�?�O?�*�h�u<����8��0�� 	�=�QO�ar��4A���x�,z��оI�����5ѾJ������ʛ>cyY��?���|���(�;����?>#,/?�>ƾ����L���eg=	g%>c��<!�:���Ǭ���$�TW?�9?�>�8"��Y��6�>c�?b`�>ݐ%>���4�-�>�?4?��-?�7�N��2�������g�?���?��@?�/K�(B�Y�	��O�h^?)?���>'\���_ɾ]���?'7?�=�>*l�韀�Ȋ���>�jV?�9P���\>�p�>g��>�0 �����6l�G��������r1>���s��)I]�)GH����=,�>��r>>Z��r�� ��>84�n�N��H�������5�<��?k���m>B�h>�>��(�Z���Ή�6���L?���?�gS?�e8?�>��&��A����=�Ϧ>���>���=v��]ƞ>s�>�P�Enr������?%<�?��?^TZ?	rm�Ô࿍쟿�w�����%*>��d=��j>�5�����=y�%=\�1<LY��;D�>T�>��>zy�>���>�>>�>�ހ�1�!�,�����&K�� �F����x���89���� ��g��'jF����=O ����	��S��x����8��SZ=��?��?��=�=M��=W��;-���'>�O���� ��˒��<��x��dmY��������� �ܹ۽�<վ/��>�Y>2��>>f>�ü�
C>�x:>=v7>ԙB>�>��#��>�o	>��>Yyf>�A�=E��>-��>���?��p$����T�]�����>�G?�赾�0c��'<���оd T>�_>&�>.Yb�����i����!�>4�=��*����f��S�>FC?��7�M�=oe<��������u?>�0�=��;�,�=Mʁ����Г=���>��.�h=��">X8?C��?�*2?�k`?��=�*<>�}�>�G�=�{�>OI>Q|(?��?2�@?��>�i�<r�J��У=�����0�va�<��ܽ�Y���Ҽ ��<�Q��r@='�<�&>v���W�>�%�@�'��	�=P.?��?B��>���>�ZR�� �(�"�J��=�!p=kfU��Y�>�Z8>�A�>ģ
?���>�� >!�#��'ƾ�G����>��>X~�������� >~�z>��>��?�X�?��p��&����=��B=���>�E?�8?&�o�2\�>,������fؿ�f��*;���X���*F�<Ǽm0ὼ��;�Ä�G@ҽX��=Q��>���>��p>'��>oQu>�!�>�8�>M�A>}9|=��>�N���c��(��j�=<���x�6=���퍓�.<ӽ���ozv����� �B����[�)�?4�?�`]=��*���j!��v7��x]d>y��>Y��>�,"?�7�>�޾7�b�ɧC�XOz ?y�v?���>4�p�c�=�u�<�|w=��>��>n�>Q�G��`��eĐ��{1=%��>�{)?�l�>��Q�J9��f��
��~��>R�Y=������? �u?3���Q����1��-J����>�v�Ŝ��־_���]G���"����t�?�o�<���>^��?�&ܾ��;��@�z����������:>�]�La<?ZV�>(3������𨸾�\Ⱦ���=�%�>�]黁\
?W�0?���>:�E?h�W?�?�-��k?�?�=v��>4��>�o�>�((?�7?�Ŏ>��>I�>�EV>%KB�]D���P=�v,�p�>'�c>K9>��>��=ym>�4���C�q�j%-=�>6<<���~>,&�=�v�>��+?�T�>-v���o��.K> �f>�Y;���>*�P���]>�>
��>D�?ū?8?����_�ƾ
��=y^/?J�=?�s�>�TJ<���̾�澠EC=���>ܕ�>�!p��&�y(ľ>ﾾ}?��>*z�=�4�>q�?ǡ>ŗ?��
??4K�����wq��Lw>2B���!?���>K}�>~fE��K5�7d��0Yk�VV�0�>r��,��x>��`>F�6<P�>.�D>�\�>��}�a��iؽ.b��ŏ>&e�>�?��$>u >/ֽ�-����cJ?�8����������վ��H!7>C�G>�����>wr��A[��k��$$9��>:��?ȸ�?qjU?p?R�l���_>x�a>��>��	<�i0��N�`X��'�!>��>� �� ����Vc=��[>(�r>$���eϾ��޾R���Ӯ�^_�z�F�b��"o�����r���>N��~�_>V���jl���侐�����Y=���vRٽ��#�Mrоo?�?�O?�*�h�u<����8��0�� 	�=�QO�ar��4A���x�,z��оI�����5ѾJ������ʛ>cyY��?���|���(�;����?>#,/?�>ƾ����L���eg=	g%>c��<!�:���Ǭ���$�TW?�9?�>�8"��Y��6�>c�?b`�>ݐ%>���4�-�>�?4?��-?�7�N��2�������g�?���?��@?�/K�(B�Y�	��O�h^?)?���>'\���_ɾ]���?'7?�=�>*l�韀�Ȋ���>�jV?�9P���\>�p�>g��>�0 �����6l�G��������r1>���s��)I]�)GH����=,�>��r>>Z��r���>[޾FOE�]I�q�����J���ü%�?Xv��t`#>A_A>Z2>��)�L6������:��H?��?O�F?�<?�ݾq 꾾���W~=�J�>�L�>�=�={���r��>Q��>�㾹h����Sw? ��?���?�O]?ۨo��wݿ���(���g2Ҿ�>p�=�Q!>����l;=r��;/�L�a�z=e�4>��}>��:>TE�>(��>�nl>ֵ<>^���� ��M��DՎ���2�hW����5���,��l�����7�������BC��Cݺ�9�)���)�A)����Ծ��=�?���>k�>�za>�i>���u�;V�=��׾�������վ������{=x�g-��J����ӾU�>�o=��->
j�>���=2�F>|Q�>A����H�=���I�ڽ�^�=-u�=j.>��>���=n�;>Л?V=���p�����T�>����?�G?'
1����E/�,g�[n9��>Q�7?�e�>Y��ڸ��!�����>�M!�:q���|����~�?��?�j�+U>A3�>Eͽ�X/0����>���D��<�4>��<�h%=�3z=~��>��A�<�m��1i��KP?ՠ�?��J?5�=��>��=��	>2��=��=s��<{)�>��@?��/?�*I?"��>������s����<�[�1_�<��6�`I~�����	+�aAE<�g,�*>��<fG��BƼ��,���������]=�H ?�=$?��>C�	?�����F��i"��ξ��>��.�Lq?��>�?�s�>b{"=�JQ>��U�m�ھ�����>�D=�wF�����!�$��Eb>9E�>��N?��&?ܕ�� �����~&�П>(@%?E1?�z=��*>��@�
���Կ̍&�ym+��`=&�����d�,	c�|�(�2Q{��T��i�<:=ʜ5>�!G>l�>D!�>T��>/�G>֙�>���=�ʩ=��=�ތ�D$��U˩���=��<�=�$��'�����<�����ʽ�
���ӽ0 �<dt?�V.?�$>�$>��0�V�T��O�?P1>�U�<	<�>��'?�3s>5t���O�z+C��a��H?W�c?m�>21��V�p>h�=�)��ӵ�>b�>��=����㽤�Y�>�=���>��:?�!�>�,��<XM�cN>�F�˾�]O>��-=��Y�?wq?=l3��૽O#��-�&ٓ�a��	A�կ=�C���B��Tn��B��-��d
�%��>�n?/�?T���U=�ϭ�f����㙿��(�>�\���:(?t�?mM�yn�����G����&��a� >C�>��y*,?y`?�?{:�?t�8?2�
?I�����>��c>�A0?C��>�T�>t�K?�~@?��&>��>O�O>�*N>D����a����=�����X>;��=��>>�0U>R�>4(
>9~�p�Q�w(�:��μ�x�=��>"?)��*>�P�>�? ��>�J���ݞ=d����r��l������j�M>��I�j�?�9_�=���>�>o��>q�v>X؏=@eɾa,��zM��|H=��\?�E�?�w;�5�����b?^�������} ?Q�=T̾p�.�r��Z��M%?W��>?}=+��>ᧃ?���>΄	?�#`=	F��?��w�k��4�>�>���>�%
? �?�D��G9����З����-M�>ŝH��M=����=��>�sʻ��=�e뽕K����>�*�!��<3)?Ȍ�>��?��> 8�=�Z��i��>[R?�����-�
�b���C��=#��>�m�>d�s=���>s��h�t ���1O�Q@�>���?�h�?��g?B���1��_A?>3U>Z�>�c�=��:}��ｭf[=9��=�v.��mc������C>%<>^�K�ʝ��m���{��9B��K�p�샾*����#��!�U!���O>J
�����о�*�e
��>�=��@�c��B��S��s������?!>c?�=�=�R�9{�����Ã��D΢>�l����=��оm��l�|��y�<\x��*��3�.�4��/!�rU�>M�Z����G�|��\(���|�#,D>u�/?d¾󼵾a��Y=|%>�b�<i�ZE��-/���
�O0V?#c9?uq��]����߽�U>΂?F#�>�!>�V��ݑ�[�>�+4?�,?����N뎿����i��m�?Z��?K�A?�N���D��`��轈?�
?>�>�$���5׾��W?��1?<��>	�����/"�$z�>��S?��U���a>Nl�>ȟ�>���;��ȧ��+卾��7�6>>%�<BS�3	j����k҄=��>�؁>�r�0�����>DW�P�N��.H������>Z�<!�?n��*>Yeh>�>��(��2��hʉ�g��BL?�j�?�nS?��7?x9���W�X!����=�ɦ>@G�>�Э=>{�|�>I��>�n辸�r����l�?13�?.��?��Y?��m�ѿۿYu���2پɳ��7O>>� R=U=��˽���=Ĩm>�[�=�+���>R��>��/>b/Q=PR�>�^>f!�>f��ƿ)�����zم���[�xs־&* ��G�O8Ͼ
�e�������C����=�ݑ�A���y⚾T�!��C��<3�1wU>��!?�?<��;��>���>�_��AYԾ���M2��},��Q��������Ƚ�*�ⷯ�Ȓ��9'���O?��=d	?>7m�>f�=��>1��>!Ƚ:[==��3>�?�>T�>w�=�>�\�>���>ũM>/��>�}�|`�������9���۾)",�9(s?6�����������2��e2>0?G�h>��M��N��w��c�>��$�0�Ⱦ��F��"�=ǃ?I��>N��WQ�=�Nr=��=�C=�6��B4�=p����=�=��$���}��>�QS>dҽ�uy>�+>�+J?��k?��T?kU�=b��>	@ >��>">>o۞>3ί>c�>�?U;V?8;?ǀ	?�nϺ&3��}�==����$0��I��4��l=��>=�J.=���=0��=��=6�G�=ECp>e@�K+���1>Du?�F?�R�>U��>ֱ��щ���/�������=֚�e�>;f�>	`$?ی�>qSw>��.�I��<}��kn侘¤>�>Q�Y��߄���*��4>��?1H?��V?�/��6Ý��_�d��=|`R?�o`?T�L?��a=�>(� ���|�񿇧>���P�<�Z�=�w���t�G�;�>��P�Wa���|M}>���>�(��Y�a>��a>�x>�C�>��q>&�8�kݐ<4>W2�(�X=i�=䰁�:f�=םF�'I����<�H��~�=�Cl>37�<�F&��R ���?d^?�h�<�H>Z�B��f�¾���>H��=��>��%??�M>�H徯dJ�w�=����=:?�&o?��>Η��P?>� >*�>�->�u�>�J>��f��;��?�TCn>$>p@;?���>��5��+`���%�3ԯ���E>��J>���/Ė?�r�?��#鶽��-��Q�����E�>�Oe���3>T��u%<�U���~�Wط�tl����h>� �>��?'�վ��>┽%�k(���}��K=0D�=���>���>�K���*����L�����������.8���x?L)?Nb?�r}?�R	?�eO?r�M��>�:B>�;(?��>�m<?ޅ?�|?�Ԃ>!#?��>��>u�K�ԃ�@�2�H��@�P>LE���1>2�0=�=�=�a�<��R�2�>����&J�_��2g=�� ����=�Ȭ>��/?�I?v��He�� /�>��=��r�%~�=��>����m�����>pqO�h�!?r)?�
?�y�=�Qd��������&�=��=?�|N?�R�>���=w���J����)�� �=�d
?����������������O�$?҅�>:�=_�>�c?�?"j�>�^�4kV�5������>v������>���>���>I��Dvg��o�$�D��оu!ݽ�]߽9p!��WP=�߹�>�=���=Z��=���=��Ľ�Y�f���q�V��2�>��s>���>�>. �=����{^��8J?.[��D9�濫��+о����Y>|�;>���?s�	��~�C��;�<����>�e�?��?O�b?{B����|\>��V>B�>WO
<�Q>�.��i
��`�3>Ma�=�<z�?������;�\>gt>��˽'ʾ�1�'TE��|��c�F��=��� �8׾s@�6���>��*2=|���S⾑V��b`��wm=�Ǉ�Ǯ���]���U��p��?l-�?��>����%|�ˤ[�Y龴9�>ò������&�!1��吽9��:����;��@���U���<�Ý�>�������Z���zH�Ym�=3g�>G$!?�-ھ�(����� ��=�?>��轗����~o������J��Q?�0?VŴ��6q�pV�=>���g��>R��>��~=�J����$fY�1&8?�lb?��O�����ψ���=��?E�?��C?4*����2�!���a���
?�?n��>�Ғ��)_�C^%����>q�D?t�=��M����1�](�>��d?BE��3g�>f�?f� ?X�=��͇���w��>���2s;c�>��l�]�=�i�����QO�;O�>�xA>l۽�ب�Vp�>m	����N���T����zkV��I
���?�J���y=0�L>Q�>����������������J?qٲ?%K2?p@>?�1޾�S ���ѽ��=rf�>���>�� =`�����>�>�侲�a����6�?ϳ�?���?��+?*6h�y�ӿYg��*�J��6��A�>wV����>�ꄽ��=�=mD��#�^=���<;��>Z��=�G�>��M>t�{>�=>�.��B�&�?���)���D-�6K��B�>A��@�����6���5�SY�������H���B-��ȉ<R��B�*�Uo;�Bg��`=[W?�	?@�=?�>��o>�ؾp���Rr>Ae¾�w��!K��3 ��ኾ�5��Ď��F�;k���f��h�+�?��=��P>�>�ꀾ�M>��2>ϫh>�d�<`�>B�9B�.>�2�>�U�=h)�>l�>l(_;��	?��ȾR헿�!��(c��z�=Er�>�@:?�gF�TU���
�f��O���>�=O�?�>i}ʾ�X��Ԅ���>tQ��TL�1PG<���<?�z?��{�-+�=�>JZ��᪚��FI;�ύ>C,�=4��=hg����~5q>�9Y>=������l�+�`�w?�)q?Q�R?�!,�]`�>�si>�J�>�b�=���=��?�~?s?C]?9�1?g�?3=x_�jZ��!���A��)g;a��M�<9�ֽT������=��=��>C�!��Ͻ�M��V�p>��	>����_	?%�+?x��>���>��s�k6�;�+�����a�c>�e��~�>;ɬ>���>j��>V�>'KX�΁���۟���3��o�>��,>�K�MPn���
���=��>>�m?��]?n���ֶ���/�,>��-?��E?m*k?>=�=n��T��[ѿp;"��%%�X�ʥ��\����d����k��:����5���սȸ=R�J>y>cq>_&Q>4�R>��>��>5rK>Ӊ;=�a�=���HT<���,`�=������4���n���a�p)��*�����
���L���#��?㼄a	?��%?��k�y�=��C���¾�&��ㅛ>���>F0�>Ii?S�l>���SJ���N����"�
?��k?�t�>��s��\>km�<��û)-�>~,�>7HS>a ˽�ӽ�p����d=ȶ�>��?ֺ�>j+����M��]���H߱>��>�uw��?�?�5��~�Z@�s�#�J�Ͱ�>�2���9��a����7C7�ѩ$�h�%��w���>��>-�?���;��):����cv�e����k�>PS���x�>�Fp>'&��1D8�{������d羹X�>E�n>��4\8?�-?�?*�?f[;?7 (?1j�b�>P��T_0?��>8�z>��;?�	?��X>�t�>��>:�>ۢ{�yT���e<�2�~�>�y����2>x��< M�;f�>�H�%����-��?�<�8=\*z=V�<�#f=P�>Q�+?<?A;����.�n��=�=���>���>&y���C7� >���>�L?�("?9�>�=CC���f��p����>�.?k�t?�i_>m�n=��
�[Ǿx"1�ć>���>{��=R��D"����H�>� �>̃����Y>�h?��?%�?k�{��^�Jv���O���=WK�h��>��p>#�?��-���X��H�f�����6�v��>�{��3�=-D!>��
>n>�q�=u�]>�k��9ͽ�6A� g|�3r��]oI>�U�=�v�>,ni=�)>�2ܾ��M���I?�����/��Ԣ�mxϾ�i�B> �>>����?�"�Tb}�v���{�<��7�>���?�=�?�fc?UvH�Y4���Z>�T>�)>��<;�:�}��3{��Fl2>���=�w�#���H��;��\>O�w>�ɽwʾI��a�M�ɠȿ�_w�.ܩ�h���{��{PO�K�#����>�g�p����#���<Aw���ڽ�	d�F�^�����z��>�����?"?5�������9��K���ӝ�uq�>ah�����+o佢['�M(���Ͼ����>־w+���ws������-�>q�`�����<S|���*��w�J>�0.?_Ǿ;ܰ���1=��&>���<���dъ��ƚ�f��|V?�v8?"��O�hzǽ�t>�
?Ի�>�	">����m软��>�i5?�#-?B��y������D�����?�-�?L^A?[����Z?�fq��焾?�'?�Ƿ>!韾�������+�>�X(?2@�>ϋ�q�O����> j;?��b�b!{>EK?���>7g(�d{��kƲ��8�����<�`5>L��<1�2l������=��o>�wT>��M� hy���>�U��3S<�c�9��N��s�j�=�v�>����2�>x �>=<�m��0���C�������?���?ͩ`??�>F������\l��tD>�Y�>��r>c��=u|�;��>h�?�)�E�E���)���?��?կ�?a"?jZ���ۿ�*���]����>�U
>R1D>������;�g编��=-��=���>��P>~;�>��>��z>��E>\w���~(��|���"��܂A�>���ɏ��З3�l:��U|��֕g�s�����I��
��ݗ=4jG=�T1��*��M5����>���><w�>+ n>�s>y�R>����H���f(��S;D=���=�ʾ����� ��e�� in��qu�����@��ys��?&�7>B��<�m�>�l�<3=%y�>;��>F�=�u�>��+=⎧>�>[�>~�>B�=	�>��5>�����������<8�G�N� ���q?ݓo�G����a�(a�Fƭ��<>�a?5" >�d;�M��f�~��?�M�=L�q�M�ŽuĽ����>�B�>1�e>⺽_�`����#*��\f���>�܎=u�-�h�:��A�>0��>�H��#=��>&�?O��?j�-?��=M�!?��>>L�>ܺ�=�>f� ?R˷>Sz?� Z?b�S?E��>j
~=a�վs�����><�u�5=+��=>>`��:�ʽ�=j]=m��yj���=��!>y����%�c< �?��;?�O�>'��>�ѳ��Y^�E�k�3$�<�>V�K=$�	?X��>M?|-�>f�?�.v>��J=(󾦒M�
U�>P>�9�Ic��z�O��J�=�+T>��$?D�A?@��=������>�#�>�
?�-$?��O?좣>iTF>������ �(Q˿�Io���Y��G��x�vU0����=Ĉ�@A���Ľy��G�ս�vɼ��>c�>�^>PXӽ�ْ<-?M�Q>�8g>˰�=�����Y��
׽q=d>t��=p�}<0#ͽ�M;��{ѽ���SL������,����ƽ��q�)�?�K?$M �9皽�bq�pZ ��ы�@��>I�>�%?&D?���=�!����T�4&K���d����>��Y?c�
?�IA���g=_�=���<���>�ŧ>�Y>Yc��D-�}�Ⱦ7��<���>��
?�W�>�
�?�F�R�\��E���>=gn���ך?f�}?� �������뾏Q��Ҡ�#��|��<�ަ�/�!�&�0�*:G�G���_˾pm߾��=>���>�D�?�@��/�@>�O�������v��'.����=���>��=������M�����Wi`���>����>q(�>!��>�g?s�??%͋?�1�>m�?G{ľ�c?	ɉ>�-I�~�>�n_?��Z?�?��>�.?���>�yo�����23�=�g�\�y�&�Z>�M�>��$�O,ռX�'��=�����Ǆ�sZv=�f>�U��ʇ��1Te>�Q >�6t>�&?�!?z����ݼ<�˽��c��=G��=���>C�>�����/?���>z��>��n?�<?v��>��G�`(>�վ��=��?�*B?��?��3=9k�>&��xֳ�����/t>��a=��������^���⽴��>�ӫ>Tm�>)W>�|�?��|?P-;?��i�sr���`��c�k��8q��ž���>5��E$���o���c��~+���C��3c�I�>����ѷ���H<�A=��
>C�Ⱥ8o�<7)�>}�������®���O�o4�>�o�>]�8?Ϥ=k��=�����I?ے���g��ߠ��jо|[�4�>��<> �ם?0����}�����F=���>u��?���?�5d?��C���\>�EV>��>8V+<��>��O������3>wv�=TQy������y�;�,]>�cy>��ɽ��ʾ�$��H�_���	�b�����T	����i�־i;ub�=H�����0���쾆���9n{�A2��$��|���9_��*Hž��� �?�?P�>����*8��v��(�ྰ��>�▾�sֽˤž�>�xi���ľ�K��:��4;�a)�y���m�>wЦ��������)�?���?��8>��y?�9>�	ﭾ����O�V罿�/=��̾劣�����jE�=a�X?9$<?�_��o���"�����!?��C?_jE�w�Ӿ��=�X�>?��;?ǫ�>�!���_��왾=�s�?NB�?�@H?E��Gi���������>�p?"��>iK�kh��E�����o>�,?+x�>�bK����\D��Vc?�`�?�N�����>�h?��?�^Խ~�E�<OH�ILؾ���=��>3ő��a����'z˾<ƽ4�>R�>L��gǾ@'�>;�羋�G��J���
�0,��S=��>n���8�+>,�>�ٮ=�	"�K䈿~!��ԃ/�1<?~�?7�W?b�"?��㾬y��T�{�%!>���>C؈>�Ϗ=q��(�>]�>k���Hu������F?!��?���?aM?vq�naۿ@��#���vy���IP>Ai=��K>1@��=\=�߫ս"��}�=�{�>���>�w�>�>�"V>�tD>��wW'��岿�%���;�h=�I��j�"���Ew�ć$�.���M���n1��I@ʼ"�F�e?���h�4�Y�㾎��U��>b�0<��>`�>��>�Ė�-M�� s>�����uM�)��@
�B�ؾ�����������s>o�(����$�>��1=P�>+)?}	>�:��>�>��;��t>3�M>_g�=Ę>yK�>��>���>���=4_���'+>�k�:.���χ���?4�[`I��ºF�M?�}�p��� :���վ��̾[U>��	?].A>�(0�9��Nw��A�>e��<9T�y��=�ڥ>H6�>�}>c���b�<Vw3�z���l�<��b>�X�= �.��.ƾK�:�R%>R�>uˆ�i>aF�>3I?IL}?]J4?GM=��>T&L>}>�V>�&�>�|>��>��#?�eU?/<?Vd�>r}c=�8f�چż�F��~/�O��<�:��𲣼V0��]KV=��=��=��t9�ԗ�[A;Z$=��(�o?��}w�=�T?v*?>�>���>��Ҿ	�,�=�\��?P�B��>F">���>�߻�@?;�?���>88�>�R�=����Q7��/�>�Ǡ=�d��ɂ��׷="v�=�|�>#�?��>V��B��>2�����]?�O?ޔ7?�Bw>��>��ﾟ���;ݿ)�\��j0�yc��WƾII�3��<�ai�
;�䢾tKt��u�3�|>���>E�=��;��7>�
>/7�>�o>�k�;-k4�N��N�������>a�=&;��o��A����D��P���?GZ����dv<�>н�d?Z�?�輼�r��e�{`�����ѷ>��>��>���>HZ�=L	�E&Z�dC�%E���>�)g?�(�>W[3��d�=X�D����<m�>�8�>|`>��t��S �����~<�]�>9<?�ؠ>2j	��Y���h���
�W��>�n�;�Y����?[�^?|�-��#=M�
�j�i��1&���X��c��,��O6��L�< پ������"t>#��>'t�?
����>!x��h��g��s!о��&��7�=m�9?Ot>��!��63������彛_;3ߎ>5�>�?��.?P�"?��?��4?��?�{����0?Wi�6��>�G�>�2?�??K��>�?�G?���>��:�]����cD�A)�O%4<ҪZ>��k>xa�<�����N=�ެ=ӎǽ�����)=�Y�5��:0�+��=�S>(J@?�(?�������=��>�Y��` ���W�>k�?��=�{	����>,|�>tw�>vt?�!E?��>XOI>J�P�MѾ��d>)�?>b2?z*?e(==�1>���ۼ���=<g��=}�.>������Ǿ|-Ͼ(�U���?<
>j�>ч>�x?��;?�7<?l�U�����ϒ��$t�L���R�>j�_?�}�>	g�Y3��\r����Q�;��E>b���%(�J�D��?�=X�ܼDs`=;D�<�ڀ=T{�=�i6>�=k��fU���?���>���>t�~>I�S>�MN��|����I?�~���m��䠾dо�O ��>o=>���ҟ?����}������4=����>���?���?3Ed?69D�'��\>+RV>k>`2</�>�d�����E�3>l�=C�y������;��\>@+y>��ɽ�ʾ*�7�G�y����7��U��fU������,Y����C�=�A����M��n������	��&g��Y:g�e,þ��̾������?�v?Z�>l6>�6O��>��0�ѾxD�<Ν����Ծ�Yܾд��o���E��<d�w�z�B�C��Z���#�H�>y���?���������bS>�^�>/^?MG�f4����-���Y�K�v=�׷�y������}x(���V?*.T?��Ǿd�����.�Z�.<��>�) ?8�
>!���?�X=��>]�?�:?�P>�ޕ��$�� "ֽ�?w{�?^�4?�����D�]?�Ʃ�`(�>s6h?��>����T���5Ⱦ~M�=n�,?C�>S�-�bĠ���B�e��>5j�?l��Z	g>{v?6�>��H����6ﴼH�5�}�u>q��>����5ps�����Mc�A[�A��>�b>����S���>�U��3S<�c�9��N��s�j�=�v�>����2�>x �>=<�m��0���C�������?���?ͩ`??�>F������\l��tD>�Y�>��r>c��=u|�;��>h�?�)�E�E���)���?��?կ�?a"?jZ���ۿ�*���]����>�U
>R1D>������;�g编��=-��=���>��P>~;�>��>��z>��E>\w���~(��|���"��܂A�>���ɏ��З3�l:��U|��֕g�s�����I��
��ݗ=4jG=�T1��*��M5����>���><w�>+ n>�s>y�R>����H���f(��S;D=���=�ʾ����� ��e�� in��qu�����@��ys��?&�7>B��<�m�>�l�<3=%y�>;��>F�=�u�>��+=⎧>�>[�>~�>B�=	�>��5>�����������<8�G�N� ���q?ݓo�G����a�(a�Fƭ��<>�a?5" >�d;�M��f�~��?�M�=L�q�M�ŽuĽ����>�B�>1�e>⺽_�`����#*��\f���>�܎=u�-�h�:��A�>0��>�H��#=��>&�?O��?j�-?��=M�!?��>>L�>ܺ�=�>f� ?R˷>Sz?� Z?b�S?E��>j
~=a�վs�����><�u�5=+��=>>`��:�ʽ�=j]=m��yj���=��!>y����%�c< �?��;?�O�>'��>�ѳ��Y^�E�k�3$�<�>V�K=$�	?X��>M?|-�>f�?�.v>��J=(󾦒M�
U�>P>�9�Ic��z�O��J�=�+T>��$?D�A?@��=������>�#�>�
?�-$?��O?좣>iTF>������ �(Q˿�Io���Y��G��x�vU0����=Ĉ�@A���Ľy��G�ս�vɼ��>c�>�^>PXӽ�ْ<-?M�Q>�8g>˰�=�����Y��
׽q=d>t��=p�}<0#ͽ�M;��{ѽ���SL������,����ƽ��q�)�?�K?$M �9皽�bq�pZ ��ы�@��>I�>�%?&D?���=�!����T�4&K���d����>��Y?c�
?�IA���g=_�=���<���>�ŧ>�Y>Yc��D-�}�Ⱦ7��<���>��
?�W�>�
�?�F�R�\��E���>=gn���ך?f�}?� �������뾏Q��Ҡ�#��|��<�ަ�/�!�&�0�*:G�G���_˾pm߾��=>���>�D�?�@��/�@>�O�������v��'.����=���>��=������M�����Wi`���>����>q(�>!��>�g?s�??%͋?�1�>m�?G{ľ�c?	ɉ>�-I�~�>�n_?��Z?�?��>�.?���>�yo�����23�=�g�\�y�&�Z>�M�>��$�O,ռX�'��=�����Ǆ�sZv=�f>�U��ʇ��1Te>�Q >�6t>�&?�!?z����ݼ<�˽��c��=G��=���>C�>�����/?���>z��>��n?�<?v��>��G�`(>�վ��=��?�*B?��?��3=9k�>&��xֳ�����/t>��a=��������^���⽴��>�ӫ>Tm�>)W>�|�?��|?P-;?��i�sr���`��c�k��8q��ž���>5��E$���o���c��~+���C��3c�I�>����ѷ���H<�A=��
>C�Ⱥ8o�<7)�>}�������®���O�o4�>�o�>]�8?Ϥ=k��=�����I?ے���g��ߠ��jо|[�4�>��<> �ם?0����}�����F=���>u��?���?�5d?��C���\>�EV>��>8V+<��>��O������3>wv�=TQy������y�;�,]>�cy>��ɽ��ʾ�$��H�_���	�b�����T	����i�־i;ub�=H�����0���쾆���9n{�A2��$��|���9_��*Hž��� �?�?P�>����*8��v��(�ྰ��>�▾�sֽˤž�>�xi���ľ�K��:��4;�a)�y���m�>wЦ��������)�?���?��8>��y?�9>�	ﭾ����O�V罿�/=��̾劣�����jE�=a�X?9$<?�_��o���"�����!?��C?_jE�w�Ӿ��=�X�>?��;?ǫ�>�!���_��왾=�s�?NB�?�@H?E��Gi���������>�p?"��>iK�kh��E�����o>�,?+x�>�bK����\D��Vc?�`�?�N�����>�h?��?�^Խ~�E�<OH�ILؾ���=��>3ő��a����'z˾<ƽ4�>R�>L��gǾ|_�>�
����
6���;64�N��4�>��c��ǔ>Ř>1�>�U�O���D����i�� ?_'�?r!J?��!?<�$��lF�d��=�ʾ��"�>f�>��o�xr�=��>��>=\��\x�0۸�22?:�?�7�?Y�?�k�l ۿ�}������ǋþgg >M�2��g�=����Ӄ>Nޫ>�O�����t>~�>mW>�?�>��>��(>�[�=���OX'�O¿�e����D��;*�u�/�Π���{�ʻ����R�ܾt�ؾH}%���5�1>�=u���Q�w����C땾52>���>�Ł>m�;>���=k�>?/y�~j��(�=�[f��[�������)����Dv޾"�ξ^��=��D�2��+�s�>>� �69�=�L?� ���޼>۬>��^>��R>��c>uɚ>�	>�Κ>?<>l�>$��>T�4=G��=����A숿s*��p�Z�6��ýW�c?/�=��]㾫5u�]9q���Ѿ���>�9�>�>585�1��nu]��K?����lr��@�5�Οo��>��>D�X>N�ս�"�ǆξ)�����=�/>)�� �+��ٷ�Z����,>!}�>䚾�M8��s>�mw?ُ?�s+?���=�?�?>�x�>.+u>���>g>�;�>��%? �V?�5?���>�a�=��������>�^���� =�wW=.WD�`<����b�a�y����<B,�.�ܽ�����𽣽��F��D��yJ?�U<?W��>{�	?� ��Uc��)%�,P>w#<�_��!�?V�M>�>�y0?g�?��s>lm�=���d7�9��>#>��T�:������f>٧�=)Ry?��J?'_-���e�P!>�>;}?-�#?�N?5�?�ٿ=�?�Nm�nĿu�m�K0���������ܟ�餀��2 >�k�=�4��lEw�~=N>���>fp�>�xn>:;��֫�Z_�>��>��=l�t��*><z�=�};�*XX=�ݜ�Y9q��!B=���=]�j�)R<}i"���2�)�9��|�\.���?f�?���3��4�n�����E�zK�>=��>���>��>��=9��D|U�d�C�r/W�e��>�Th?|@�>&�G����=
�e��zM�3ո>b�>:]�=����������<�:�>z?'��>8�ATV�m�k�W���R�>��2=�p
���?�o?�09�F\=�����'e�;������kl`�;
��Ѐ ��D���9�o�������c��qc>��>�Ω?`�$����>�eO�=?���@n�HV��8�,�瘬=R>�>k�ھص�����D���"Ѿ�����>�>�kR>y{�>S�?�r$?���?�e?+�?��ǽ�R�>?Ra���?`��>��;?;��>�r?M��>��	?$��;����Q���B��9�>�c��~��<�v�=��>�5=}��=�';>��4�����8�L=5�<k��s�=@&=Vgf>�J>j�,?�C?�-���W�pϰ=�=Ͼ^�G��>Ŏ@=GI����=Uf�>@�>?��d?�J?��?l@��W�>���Ͼ���=��?�*?�?g�=��>yY��GQ��H�E�U>��L>[�����������Sc��AZ>�_>�+9>�LZ>9l�?�ك?SW?B̋��课�e�*�^�V�>4s>��>��.��&��CU�%1�"�*�i�N��4�DA�=v
�g	�=w���#ی��Ց>�j�g�>^�>��a��>m@8>@��j�?��l>�9*?�a�>U��=�W��ѳ
���I?�����e�젾�wо�?���>�<>s��S�?����}�_���B=���>��?���?;d?��C�e%���\>2QV>{�>�!/<�>�D��򮅽�3>B��=��y�����Ξ;��\>B7y>:�ɽ��ʾ�.侎dH������ _��ᖾ�s��.����˾-�Ǿ��0�=�9��D*��=��q����2w�ku½�L�
|���䶾6�����?1�d?c�=<��a�,�3�;��|x>�+m�ۥ�����r'D����*x���wu�*:������Н�>�ɾ�����Ι����ܾ�>��^>��7?9���'�N�r��Q�=�B�= �=_� �����(��ü��[?_�4?G����3��g���+�=@�? s%?�I���	�=Ԟ�>��?�]+?�?]=?녿�%��������?�#�?��;?���'����"��:��%�>��?�2>�y��Z����Z����>��?V?ɗR�����%�(�d?�J�?:vZ���>t��> �?���� C.�C��	��d�}>)�>><�7>%��g���	�����c�X��>s��>6���;�����>Z较,�lq9���
���i��BK����>MR����=0�>��>�N,��z��$[��7����?3��?�BT?η?����/8���r�;̧o>JB�>�\�>�( >�G��fu>�'�>ʶ�=�P������@!?=5�?,2�?l�'?� v������I��%'�����qf>�&=>��>N�g���1�:�=hCɽw9�&�d>=.g>��[>���>��/>�K=�1>3���v��_���{��^ Y�b�!��q.�5&n�8�:�8�(�����KľY🾬�5�<^ƽ��L<V3�����C���X�j�=�'�>,�>�nA>[׽>�N�>����������Q��/m%��2�����ھ!�˾��8�Vb��Z�>�I�ټ����ȗ>�:>j*=�s�>���=QGa>v:?[�=�>)��=�{>t�?�?y$�>�|�>��J������C�P�վ�#���%��g�
������վ)�?�L=���\�����������>��>�f�>gU6>L0�K"��Z}~��0?��J���˽��%��Ku�>��>S��>!˽��ƾ����j=��K���=���=�擽��,�H!��w��=��>;����5-=�v>l�O?��{?��W?�����?��>C(�>�{>\��>�"�>j#�>q$?.JQ?��5?�?��=��m�^E��C�R�i���=A���[���l��`=��>�2�f=m�>Y�����*�0��=���<}�l�>�?˾?�R�>Kq�>�'�:�9�62������>��=x-?�-�>)�?��:?4�?�>	>T��=)e��_-�$�>)>�	w������Bֽ9=�i�=�mG?d�?��j������>"�1>A �>I�?�~W?���>�Ď>t!z�m\�7ҿ'�3��}-�����v���M�P��+��2ڽ�w�=pF��P0��Q=��X>I�>�Vo>��B>�Ǐ=���=th�>eb2>�Q�=�Њ=ObN;������&��=���<#V=X۝�Mx��(5�4���C�D�I_�9���CT�X�k�}V?�.?́)��q��ܔe�49������c��>��>�>$��>T��=�����T���@�[QE�Q��>��h?�5�>��8�G̿=�O,���J;.r�>���>c>��d�Գ�%G���<(��>'�?)�>6A��:[��-o���
�J{�>��ؽ�~ǽJ�?w�v?���I�>KF�Ԩa�%%�$ܑ�f7�N�ܾ�;)��>��?7�b��������;5p�>��>Ԋ�?��!�]��<ۃ���*��=Ď���;s�-=�mY>�C�>�μ)s������0�S�ON	��>�4ޭ�^��>x�> ��>iH�>.�)?���?<��>$];?�P\�;?-de>Z	?@f?:?�c?��,?J
?��?hE�>�;[=���
L��\�v
�Xyo<)�u>
�e>�F�='�=�F&��������-�=��+=�׽��=���=UA+;A�>�Z??䍾��,�>��#�Bd5=��A>���>��>��_���)?g�>_(?՚M?��>?*B�>4Y>P�=��H�����=7?:A?��A?V��<f&+>9��W�G�.G�=�z>6��<�}w�b�о�C��.��TL>ɳ_>�nm>鯜=wk�?�ρ?C?���������r��mA>��7����>p0��TOV�쟑�[�q�P,�Ri;����>`�s�b���_%�;��	>W� >��B>���>�=��ž��-��Fм�λ3�>���=�>�M>�y�=h�བྷ���� J?�_�����w<��F�о;v"��c>]=>�����?��Bg}�RХ��<�D��>ׂ�?��?�Pd?s(E�?��6<\>[?V>�7>�9O<�?��	��v��� 3>��=�z��o��%l�;�r\>�Wx>�ǽ4}ʾfo��I�u�ſf4w��/ľS����xҼ���̾�:;a��݄�<\��������RZ��C�?�r�ŽQBi��F��	Ǿ}��?
F?M�>�G<�.��3������M>���a��� վ���iȾ�cw�=�y�̪�gC���'��Es�>e�ƾA���_���I0��"O=KL&>��g?�Z%�ܡ��L"��~�=Ɔ׽���<�˾~��i���-���@?5&%?d�_�(�A��e=�����>J�
?�Q��t#ܾG�D�NA
?��0?-y�>KE����W����/�����?�W�?�u/?��s"�^��ȓ�O5�>0 ?���>M���H¾����c>?�c?
΁>���	��=�I��?��r?���q��>�
?�u�>_,@�`������"���Y=Z<�>XԈ��K�+��� ����˻�l>-��>�U3�P9��o�?Q%�z�q��YK�������>��=�i?��.�0��>�ן�B�o>t}X��}]��+��M�����G?G��?pI�?|�?�gþU�B��:>Yb����=q��>D�/<0��=��>Լ,?{�¾�D9���uN?��?���?L'1?��f��9Կ��6���W���r�<V�>zS>
5a�%��=�Eܼ	H=��q=`*)>}��>R=h>��?>��\>�>�ڹ=1���(�*����������kV��,���J����������i�[�Ӿ9���|����I��-��阽�1�:�[�����C������=#�4?˧�=[\�=��F>�k�<���oƾ��0=��UP��L ���F��#�i������s��t@��ݱ�"���jK?CS=��p=U��>��K=��=�B>Z��^>�^�>y�#< kg>L�=G�>�!A>c=\��k�p>yK�=<킿uj~�-38��d��~��;>?�"Q��0����-�-H˾H.��I��>P	?�!`>2"�)ѓ��:y�?G�>��\�)tk���潈JD�^Y�>dϾ>���=&�E;5H�!������dx=���>��>�ػ�^��L��݊�=�h�> ���U-+>�*T>�*?�{?�8?i�<���>0�)>�2z>lg�=��T>�9>m��>�`?�~A?��-?���>w3�=������=��;��9��<��*�O��u��Q�~��T�y��=`k�=݆�<��=��P�M�;>�l=)�	?'8Z?B�<�V?���}o`����sF>KQ�ꊹ�^$�>^<?P�3?�� ?�?@x>=5S��-�5�%���>,<>8I�T����|> ��>n�E?;��>4r�Yo����>%�?�q?W�? C+?�}>�#>��ľ%	�ρֿ]鳾�-	�z��=J̽���F��3۾�S����`�N�/z�ƴ�<��q>�om>�>��v>�g�=��=A-�>��>�Ǖ�@,�=/>�v��^TD=A��=�=�N��I��y\P�;��qTL������s=��r<�"?=��=��?��>���=�4�=�Ͼ.y�)�S���>V��>F'?���>\ ����X�h�Y"-��Ԫ�SL�>K�k?��?�r��B�>2�Ҽ�#�w?n��>�?>�'[����+��'�ľ���>�F$?�5�>�W�	텿C����z��+�>�2�=��֠?��?�e� �'�<6@���"�����:>\S��ۨ�j6;y�>���F���v=!��B7���>[�?ѳ�?:��M�>�ɾ�&���{~�Ҏ�=��>N5��bh)?�)�>>C��#
�b���2`�/�ԾB������>�y@��rF>�V?�)?i)�?�q?��x?���j�+?�5�.��>D=Z>�="?6�?��?H�	?0�>A�7=��1���UƾE��ё�>N�'>bL>��?>�
	���<��=>��>�*B�D��<���>D��=O��k�h�f�v<�×>F(�>Y�~?�90��R=�L>s�о��=Η�=��>~g9����iq>�> ?l;9?��y?�"?'��=�;���.������=n�H?@�
?�s�>��]>䶇< �8�e��:v�\��N=�/f�=��`��V��d+O����>��>%��=��>�ys?k�,?�?,���5�YM��D�#�}�;�^@�'�>���>�M0<gG|7��wm��|_�]�-�/?^;��"���,�h6�=dg>�T�=7�l=N>��@=��`����b�=� 4<�ҭ>�s�>Dg?ŧ_>af�=�Ծ�����\Y?�Tվw��r�/�&�>��I!��ۋ>��e>�ʽ~�-?�6> ����Ǟ��@]�6�=ݩ?���?���?���͡H��~�>I?Fh`>�Z�X����2t��W���|>_>;���B�ܾlk>��%����>KS��i������ng=��(��(9���a���
����nK־��
�O��j��A|��/ʾ&�2�쮧�����dy�G�2��d&�u;b�+�����?"p�?Ĳ˻-�R��b/�����"�v>e��Ț�%ھ���q�ľ|V�4��(��!;��3��M�8ġ>�䡾���䵏��Ҿ�]>��I��79?} ���ὶ�_���=%�9�DB��0�,��&��t��k�6>��m?��h?�}ƾ���H��
y�>��&?>�>��>����]|����?C1�>�F>�^�����6��x�?q�?�.M?ƇԼ�sh��L �"�C�R��>�;�>.*T?��|�M�+���E>�)?vW?;�?�X�([��4�Ğ�>F�(?��?��!�>�i�>��>3젽:�����½Z��9�1�%�?j|�<��������� (��̈́>5J�>^�>�澾���o�?Q%�z�q��YK�������>��=�i?��.�0��>�ן�B�o>t}X��}]��+��M�����G?G��?pI�?|�?�gþU�B��:>Yb����=q��>D�/<0��=��>Լ,?{�¾�D9���uN?��?���?L'1?��f��9Կ��6���W���r�<V�>zS>
5a�%��=�Eܼ	H=��q=`*)>}��>R=h>��?>��\>�>�ڹ=1���(�*����������kV��,���J����������i�[�Ӿ9���|����I��-��阽�1�:�[�����C������=#�4?˧�=[\�=��F>�k�<���oƾ��0=��UP��L ���F��#�i������s��t@��ݱ�"���jK?CS=��p=U��>��K=��=�B>Z��^>�^�>y�#< kg>L�=G�>�!A>c=\��k�p>yK�=<킿uj~�-38��d��~��;>?�"Q��0����-�-H˾H.��I��>P	?�!`>2"�)ѓ��:y�?G�>��\�)tk���潈JD�^Y�>dϾ>���=&�E;5H�!������dx=���>��>�ػ�^��L��݊�=�h�> ���U-+>�*T>�*?�{?�8?i�<���>0�)>�2z>lg�=��T>�9>m��>�`?�~A?��-?���>w3�=������=��;��9��<��*�O��u��Q�~��T�y��=`k�=݆�<��=��P�M�;>�l=)�	?'8Z?B�<�V?���}o`����sF>KQ�ꊹ�^$�>^<?P�3?�� ?�?@x>=5S��-�5�%���>,<>8I�T����|> ��>n�E?;��>4r�Yo����>%�?�q?W�? C+?�}>�#>��ľ%	�ρֿ]鳾�-	�z��=J̽���F��3۾�S����`�N�/z�ƴ�<��q>�om>�>��v>�g�=��=A-�>��>�Ǖ�@,�=/>�v��^TD=A��=�=�N��I��y\P�;��qTL������s=��r<�"?=��=��?��>���=�4�=�Ͼ.y�)�S���>V��>F'?���>\ ����X�h�Y"-��Ԫ�SL�>K�k?��?�r��B�>2�Ҽ�#�w?n��>�?>�'[����+��'�ľ���>�F$?�5�>�W�	텿C����z��+�>�2�=��֠?��?�e� �'�<6@���"�����:>\S��ۨ�j6;y�>���F���v=!��B7���>[�?ѳ�?:��M�>�ɾ�&���{~�Ҏ�=��>N5��bh)?�)�>>C��#
�b���2`�/�ԾB������>�y@��rF>�V?�)?i)�?�q?��x?���j�+?�5�.��>D=Z>�="?6�?��?H�	?0�>A�7=��1���UƾE��ё�>N�'>bL>��?>�
	���<��=>��>�*B�D��<���>D��=O��k�h�f�v<�×>F(�>Y�~?�90��R=�L>s�о��=Η�=��>~g9����iq>�> ?l;9?��y?�"?'��=�;���.������=n�H?@�
?�s�>��]>䶇< �8�e��:v�\��N=�/f�=��`��V��d+O����>��>%��=��>�ys?k�,?�?,���5�YM��D�#�}�;�^@�'�>���>�M0<gG|7��wm��|_�]�-�/?^;��"���,�h6�=dg>�T�=7�l=N>��@=��`����b�=� 4<�ҭ>�s�>Dg?ŧ_>af�=�Ծ�����\Y?�Tվw��r�/�&�>��I!��ۋ>��e>�ʽ~�-?�6> ����Ǟ��@]�6�=ݩ?���?���?���͡H��~�>I?Fh`>�Z�X����2t��W���|>_>;���B�ܾlk>��%����>KS��i������ng=��(��(9���a���
����nK־��
�O��j��A|��/ʾ&�2�쮧�����dy�G�2��d&�u;b�+�����?"p�?Ĳ˻-�R��b/�����"�v>e��Ț�%ھ���q�ľ|V�4��(��!;��3��M�8ġ>�䡾���䵏��Ҿ�]>��I��79?} ���ὶ�_���=%�9�DB��0�,��&��t��k�6>��m?��h?�}ƾ���H��
y�>��&?>�>��>����]|����?C1�>�F>�^�����6��x�?q�?�.M?ƇԼ�sh��L �"�C�R��>�;�>.*T?��|�M�+���E>�)?vW?;�?�X�([��4�Ğ�>F�(?��?��!�>�i�>��>3젽:�����½Z��9�1�%�?j|�<��������� (��̈́>5J�>^�>�澾������>����|_�z�,�w�����K�t�AW�>�����Z=�Ў>7 #>Ua�b��Wy��@��Uj/?�]�?��3?D!?N�����62+>xk=d�=>)��> o���ü-��>x�?�0���Q��^Ⱦ[�?���?D��?z<M?�L�U�ҿUߜ�ξ�fþ�<>u�=>{>��i�5�>��;IU 9f����>���>7r>���>��U>i1>H� =����*��Ͳ�b ��|a������v�}����۶�����#���u:��R[��2u&��B�;I/���e���;b����g�<i�Z?N��>��>� >�n������޾�Đ��Ѿ���W��2;�n���B��,s��qP�]���w苾s���Ծ��?4N��Su>@U�>U�	����=���L���J>=�>�P�>f^>�Ǻ=�!=�B~=!q>�>�=p�<P>sρ��2b�lL��
	�%�7?�z<'���g�[�n�˾n����=��>�vu>	��@ݓ���B��W�>a�=�4 �{D��|�<�d>��>���=ȁ�<�=���t��=2>!Z�>5<�Q��nɼ��쟽,�O>�m?w�ؾ ��=�q{>���>�ʇ?��h?��)>��>���=1��>f��> d�>\�p>�9>��>nQG?.?��>�v�=�'���(8����<�Q�����=���<�^S��н1]��+�d��&�=o1>J�=�PL={�Y=\��.��<	�>�:? ?��>.�?A�d���;�^���ȼ�>_�P>��>A~>$��> �>�V�>��=�J>�q��������>뵑=4TC��@Z���K��n�>��?=�&?"8?e���� >5O�>�9�=��>w��>&v;?�B�>�>LS������;ֿ�nV�0�^�P�x�]n�=��=y潘,p=�6��X��`8�:��!�t>��>�< ?�ϖ>X/���}=�8�>SS�>�bT�{���p�b��b#�r�>�3=��P<�
4�t��:���&������=�9���m	=��:��<�-?|X�>�n�=��>Dh��	�����4��>��)?��!?.+,?v��=��|H�(�,��3>U;�>s?,?�O?7�N�l]>>҅	���Y�)g�=QJ�>$$�=]J��JMB�����ڽ�?���>���>�ϲ�Q�]����(L8��#�>H6=�m8����?��t?r����p���#��	@��!��B$>I��atξ8�������^���>о:��S��=t=?J5�?^���_��>��ľ�9��V�:������CC=�W>ao�> �^>�W�i?��9� ��x�r�<��=�	�>��f�-?l�>�,�>j��?I� ?*��>�����?D��<H?D>�ޟ>��C?	m?�
B?S~�=$s���� 1~�������F�@�ު!��^<�8s>9�>ַ�Ӟ>$�Ｖ1.��슾����,O=l�h�1>���=K� ��k�=�+ ?�&K?����gF��˂>����h���F�.V�u}>���񽎘u>:��><?�?|?+�>��	���
�(=�J "��M�>& ?�l?DK?)U�=�V>=u�'��l���a>3�=�|�4�-���i���~�½��>���>�o=}ի>���?ȏ?m�*?~F����9�ء=�>����A>?�>͛>2��>�=M>&�ƾ�	�Cnl�s.0��$7����>�m��К���>.JK=��+>��=+~=�T�==�
�S�1Zӽᑽ�,->�Է=�/�>���=r8+>]O_���B?U�ݾ95�k0�:��ܾ�r�`6>Gq��6=�<[�4?�n>��~�����M8��j>�?f�?�N�?���Sh�f?�>���>��>�#�=�詾㠽�1ؽKt�>�UW>�7���.پ�r�>�r>��H>�+���վ�7޾47��h¿��(���ƾf����P�w�澡ӕ����P������H�8EҾs���ڽ_%u���=K�Z<"ξ*��f8�?1�?��r>���=�߼��;�Z1���=�5P�1:��оU���|ؾ���z��g���-�)�쾮Ⱦq�M>�p7��r���������%yp��|Z?fa����y�7��ϕ>ܾ켥ⅾ޼B���R�����_���dR?duY?B�~���֗=��Z�H�)?$��>�c�=@����wD����>��*?��A?�.Z�z�r�KE`��۸�t�?D�{?3�V?Ɣ����%�ʾm�A�L�^?�`W?�' ?�2�X4.��P�=�V;?��U?���>��z� �N�uT�>��1?}�c����>�F]>-�>m�G>���������·=4�>a�K=�i��U��E��=�2#? /~>VG�=�����qp�o�?Q%�z�q��YK�������>��=�i?��.�0��>�ן�B�o>t}X��}]��+��M�����G?G��?pI�?|�?�gþU�B��:>Yb����=q��>D�/<0��=��>Լ,?{�¾�D9���uN?��?���?L'1?��f��9Կ��6���W���r�<V�>zS>
5a�%��=�Eܼ	H=��q=`*)>}��>R=h>��?>��\>�>�ڹ=1���(�*����������kV��,���J����������i�[�Ӿ9���|����I��-��阽�1�:�[�����C������=#�4?˧�=[\�=��F>�k�<���oƾ��0=��UP��L ���F��#�i������s��t@��ݱ�"���jK?CS=��p=U��>��K=��=�B>Z��^>�^�>y�#< kg>L�=G�>�!A>c=\��k�p>yK�=<킿uj~�-38��d��~��;>?�"Q��0����-�-H˾H.��I��>P	?�!`>2"�)ѓ��:y�?G�>��\�)tk���潈JD�^Y�>dϾ>���=&�E;5H�!������dx=���>��>�ػ�^��L��݊�=�h�> ���U-+>�*T>�*?�{?�8?i�<���>0�)>�2z>lg�=��T>�9>m��>�`?�~A?��-?���>w3�=������=��;��9��<��*�O��u��Q�~��T�y��=`k�=݆�<��=��P�M�;>�l=)�	?'8Z?B�<�V?���}o`����sF>KQ�ꊹ�^$�>^<?P�3?�� ?�?@x>=5S��-�5�%���>,<>8I�T����|> ��>n�E?;��>4r�Yo����>%�?�q?W�? C+?�}>�#>��ľ%	�ρֿ]鳾�-	�z��=J̽���F��3۾�S����`�N�/z�ƴ�<��q>�om>�>��v>�g�=��=A-�>��>�Ǖ�@,�=/>�v��^TD=A��=�=�N��I��y\P�;��qTL������s=��r<�"?=��=��?��>���=�4�=�Ͼ.y�)�S���>V��>F'?���>\ ����X�h�Y"-��Ԫ�SL�>K�k?��?�r��B�>2�Ҽ�#�w?n��>�?>�'[����+��'�ľ���>�F$?�5�>�W�	텿C����z��+�>�2�=��֠?��?�e� �'�<6@���"�����:>\S��ۨ�j6;y�>���F���v=!��B7���>[�?ѳ�?:��M�>�ɾ�&���{~�Ҏ�=��>N5��bh)?�)�>>C��#
�b���2`�/�ԾB������>�y@��rF>�V?�)?i)�?�q?��x?���j�+?�5�.��>D=Z>�="?6�?��?H�	?0�>A�7=��1���UƾE��ё�>N�'>bL>��?>�
	���<��=>��>�*B�D��<���>D��=O��k�h�f�v<�×>F(�>Y�~?�90��R=�L>s�о��=Η�=��>~g9����iq>�> ?l;9?��y?�"?'��=�;���.������=n�H?@�
?�s�>��]>䶇< �8�e��:v�\��N=�/f�=��`��V��d+O����>��>%��=��>�ys?k�,?�?,���5�YM��D�#�}�;�^@�'�>���>�M0<gG|7��wm��|_�]�-�/?^;��"���,�h6�=dg>�T�=7�l=N>��@=��`����b�=� 4<�ҭ>�s�>Dg?ŧ_>af�=�Ծ�����\Y?�Tվw��r�/�&�>��I!��ۋ>��e>�ʽ~�-?�6> ����Ǟ��@]�6�=ݩ?���?���?���͡H��~�>I?Fh`>�Z�X����2t��W���|>_>;���B�ܾlk>��%����>KS��i������ng=��(��(9���a���
����nK־��
�O��j��A|��/ʾ&�2�쮧�����dy�G�2��d&�u;b�+�����?"p�?Ĳ˻-�R��b/�����"�v>e��Ț�%ھ���q�ľ|V�4��(��!;��3��M�8ġ>�䡾���䵏��Ҿ�]>��I��79?} ���ὶ�_���=%�9�DB��0�,��&��t��k�6>��m?��h?�}ƾ���H��
y�>��&?>�>��>����]|����?C1�>�F>�^�����6��x�?q�?�.M?ƇԼ�sh��L �"�C�R��>�;�>.*T?��|�M�+���E>�)?vW?;�?�X�([��4�Ğ�>F�(?��?��!�>�i�>��>3젽:�����½Z��9�1�%�?j|�<��������� (��̈́>5J�>^�>�澾���Cjf>���J�&��o-�$����4���=�>D���=���>i>�V"����y�8%��jW?��?@�?[�>3sG�!G���1E�/C�����>�c�>�ތ��u�>j��>%3��D����"�(?��?�p�?�c?*�X��㌿2ؔ��9����=T�>��N>�m��%��=
�)=?�f=�=0/>�>$�G>��V>i�;>J>��>}2��|�!�tx���]��z�L�����M�ǖ+��m��|n��>��ě¾<߾��0�8�۽#eݻd���+_�ƕ/��<�x�Y�??T�>��=��E;���F�3� �[�C�&�����(��d ��� �m����f�~�P>痆>>˾��<��Ѿy�?fQ>]�$>��>�>����<�+�=��ýK��=;=	=�>#|�>,��>I'�>�c2=��>g�<���>ƽ�=��b��qc��ɾ�7��֩�"�_?�����&�+�*�,|�6���d��>N7?2��>�N�;���S4�/��>!E^=<�ܾ�a��*�<M�>�>f>8<}>\I>9���|ӾaX>�-q>��j>(�<hί��*���*i� ��>1��>��о8��=B�`>�:"?1r?%6?��=�4�>��j>�#�>"��=��G>.he>�d�>��?��/?y!*?@��>J�=PaK��ٚ<�2�<L0��T#��>˽ՠ�<uvǼ�-Y=�&o�PW�=<�c=��i��04=P�j=r�.�K��<LH�<ʷ�>��
?���>XP�>�>:�s/�q�,��D����<f�
=?r�>�}:>q��>��?c?���>L&��NþZA����>�qu>Pr�8o��$�<�E6>c)�>3�U?�dH?�S���L��X�>8Y=H�>���>�?X��>��=�hc�&��ղҿJ�"��;"��Y����(�S��&�9��[���:2�/�f��+\�<�_P>��>|+k>3�K>pH)>�->�D�>yKE>p��=��=h<p��;C�<�׾0=�W��t�;��R�����R���<���j����S�P�Z�n��(U���u?cN'?�L���st=�/h�����ձV��b�>G]�>���>X��>q3�=�	�Q�R�K�=��K��c�>MU?��?~���̰=>�Q4>K��=���>�@^=�1P>}:�����Ͼ,N=��>K~!?�3�>�����l�r���߾�8>S4=
ݽv��?�^?D�������E��J��B�<'�ɽ��\���������}5�ޅ���� ��]��3�=�.�>��?{=t�H��=����-��Ɨt�mT���Ơ=�=�	�>��3>�z,���B�k�ؾ�ʆ��z^��p>z%�����>��2?d	?PWe?�U-?<k? N�ǝ#?^��=�??r	?;�8?�?��>~m >k�&>�ė=$|�.�<�[���\�=<�Ľ��=��e>�̇=�>�=�_$>,t;<���=iJ�;�^��0�<R-=]��=��>� �=��?�B?m���Ľ�V�;�i>'�'�`��>�-D>O&�>����C䮽U��C�>�F"?9t?~�>>�N��}[������[�>K��>_I9?�$$?� ?��l*�R琽��ru!=��>��=������R⾇�I��	Y>A��>;	>��<��?��L?F��?_l�>�*[����s〿de[<�k�{'?y�?�e�>,佾��r�����L��n*,�9ܱ��搾��="PI>Qn�=?���I�>�����2�I_�={��I�\>��I>���>���>���>Kc�=�xƽ�	�"��*?��w��8�������$�;>�
=>�q��Q?W2b�W�~��3����&�&��>{��?��?��f?3NU�sɻ_>�'>�z=��/<>A� 5���<���f�=�}>����|��6׼�	�>�L�>(P��c�Ѿ7���� �,~��o[�l����̾�XǾ従`��5f��ɼ���6��+������,�y��`��｠5��l ��ֲ���~?�,i?@�=T�޽����ܾ�w��T�<.����7�l����[��.z��03\��a����!^4�M�$�l��j�>��D�Ҡ��ZW����؍>��&>yKS?�!�w�&��oD���Z>T�>c�>h*��<U��ᒿ T��Q�?O�5?z;4�3�����\���`2?��@?���g6>�c|��X=l�?�-?���=�o�]Us����M��?�g�?<�d?@Qž2 m�>�B��d⾤I?�w	?a�.>O�>U�8���̾L�?�43?�t?�I�E�O�9.���Z>]�?�^d��V�>� ?��>P�|��~p����rB��{*_�=��>9�>xٞ��i�Iϲ�[M�=BW�>Q?6V��f�Ѿ�M�>�1پ�,���9��7���ݬ��}(<�^�>UN��=x�I>��=3*�~�� Z����ɳ@?�X�?QnJ?�E+?99��wG�F?����=�V�>\��>�V�<����>+��>�%�u�(����B)?���?sW�? G?(p�FϿ>���wɾ�Ư�Tm>'�ݼ4��=NQ�o�7>œ>�	>@E=<�>i>�>��=�&�=���=3؉>�f =XQz�	-0��i�����kD�$�8�cd.�������q�z ⾆�ɾ��骿���ར~Ƚ��!�>��<9�ǽ� ��=J G?���>���>��>�X>Mv۾�0E���ٓ+��֯��? ����=`���M3�ː�Y�����~�Ⱦ��>��==�D>��>��/��ߝ=�u>DJ~=u�>;�=d�ν/L����p<��=�:>|�]> 7=���>%���\W��؈��뇿d@Ծ�>V�1?1��<�]Ƚ&�ؾ��;�=ľ\�?�P?b�>~�ܾ3���#"�\=u>��{��Ⱦ���gU=J�>D�.>��<}?�<E���|m��Ƃ���>p��>��>e�ȼ_����A��>9��> �����=�ɞ>�7?:�|?H'<?Tۦ����>�>ꚯ>�/>b�4>A�9>{��>?��"?7�6?u4�>���=�/��v=�6�<H��g�;-�U��!=��&;{`�<����g�}=�N�=��<���ܒݼ��<C{�<"�|=Ap�>1N?,��>�G�>=^M�4
<�ǜ.��y���>�y���$�=���=(A�=@�.>pL�>n�>��H>�u��_�����>G*G>�@��oM�0[��&�<�A�>��G?K�A?=k�>�Ц��>���=<?�D7?`3?���>hS5=�)j������ܿ�bO�2;	��0����� F�+�>�� >�>{�=sx�G�->	W>a�!>"�M=�{6=�i>��T>F��>�1X>m;����>
��=�&c>Q0��ُ>]ݼ��a�g��=�9=��Bwy��I=�kI=��+�����"P�=A��>��)?���=
�>=����h���c��q=^s>���>���>��>~)�����3�e��S$��_M?"#�?�ht=f�4����=�$����?�"?S>L��>�N�=1�V�?L��d	��q�=��>X��>�s�>�����nU�ɗw�Wx!����>��6=D�B=�И?��W?^Ǹ�`K��&�о<�D�+�"��n�����x���9ѡ�M/*��L�I@�]��ݷ&�N�0>2��>=��?3I�����a�߾��-�o��n���f>*>>��c>�^��o����X�H ��x�{��fE�N`4���^>��= #�>U�?�C?2�f?��?�?�&1�Gj�>���=���>���>�?�P	?g�>q�h>.qM>��n=�'R�����z�{t=m���F�=�dC>R)5>ҍ�</YN=(tJ=?�:=D��Y ����<T�����;�6�=� >��>�?-�?�Hȼ^�ǽX"�my���=Χ����<��w��$h�ȟ�=lX�<���>S2.?%6�>�/"�����?���ݾ>��>@G?%�m?.8E?h�>�D=>z��[U�4���ә�>�R�>�����=D�~����%~>1?��'�z!�=|˙?��o?��*?�4y�V󟾬��U7���Q��o'����>��>��>��Ѿ2Z^�wЎ�6}���nU�HażQ����r�B"�>�>u�I������0#=��#>��==w
?>�Ħ=^�ٽ�ԣ>}y�>�
?��=><�����	�F5+�H�1?_i��陽��mC�:R��9;���l�= ��<��=w?Y����.o�n����P�c��>�\�?���?KX?���=*<�+>���=��=��&�2.z��K�=&.>�~�>�tE>�2�'�t�����j>�uh>�^@�����|����z����(R�C���5���a>�#��%[�;7�>R�<=�:���6dB>����|��F�G%�e����V�wL��T�?~S?�n�>E,>�I�.�#�ޢ���.��]���{��`�cř=���s���V�q�iz����پ�1þ�Z���$�>�$\�����\}�`�'��W^�ӟA>*|.?Gľ�h��H���d=��,>�A�<M���R��Ls��z`
�U>W?-�8?�:뾊�� �5&>��?�n�>�&>�������Gf�>�4?�-?T5ļ@��k���Ι�Fһ?��?�=?[���U]�q�$�� ��~?��?Q��>�%�����?��h��>
~�?`S?�{�2��ڂ6�s��>�i?�76�k�G>AA?�y`>������B����l��`*�� �=��,��ؚ���5�2RD�-�pN>{z�>zu޽����>$�龲�N�|7H�n~����J�<�4?��P�>3zh>_�>�~(�����i����V���L?�b�?�IS?�38?�����"n��3	�=�>1��>A�=���ޞ>��>�w辊\r���"�??�?��?0Z?�um��fȿ
���KI}�����ieټ�?���=N>�Q��X�=�>m>�I�=H �>`�>�w+>2`�=��=���>D\�=�2x��,��������gw����m�ɾ}�J�������_��U�E���N5B�\�Ƚ'�ݽ^���;��O?���T��$X>�-?/c�>Z�?W¢>�Z=��C�������0����ù��mY׾s徧B׾ah���<]�`7�ܳ�}����a?�D�:ũ7>��?�cd�V>���>�`�=���=�2>��A>G>J�=v�=!h�=,[�=CÓ=���>���߭f�Ń�U]��-;d��>�|F?�{C>�B��~��:۾�`.���.�>��4?��z>l���j���BE�>"���jK��8Z�]&\�(x�>�2?
�>5�+>>	���0��V���X ?{��>�Jv>Qw��_٬���>��> �Ӿ��	>�?y>\s?F�w?(,4?�=�H�>�r>�;�>u؜=	�;>qU>Hv�>��?e�.?i�(?�Y�>�ж=�yL�,����W~=U�/�	�4��uؽnd%�����7�;���1�{=ȳi=�o[�A�=hT�=�:+:���&=�	?	'?͚>��>;i;� YA���-��[�e�M>adS<�֫>�U�>���>�I�>���>��>T
���ž৺����>�v%>>}\��cb��n���=�">�7?�*?��Ͻ>�����U:�f�>&��>P�1?1�>���=������࿚K��[ I�Igþq��=�T�=�LV<�����?�,�>����>P6e>-��;�Q�Vq�=!�>¼;�w�>��>L���כ>��N>�~>H��7JM>#�p�R`>��">�H=��I��Hнڧ��M�?�ӳ�=Z���N�=�?�(?& ��E&�<R�P�؍羽P���[>[�>��>�u�>0y�=���__�U_I��X���?��m?K��>:���O�<��A��s*�O�>�A�>}�D>H��T>�����> �=`Ԋ>R�?&��><%н�I�!KR�b�f�>��>iJŽ�G�?��j?�[ži�ֻ�=�ӬW��E�&[}�v�佱d��顩�z6��� ��¾��پ	��R�B>N��>��?��Y�(>�>x������Az����2����=���>��=��7�ɾ����x�=Q%�=�K��� h>��=���>z/?M?�^?Y��>`K�><���eQ�>#�6=~P�>���>�f?>C�>P��>�9>�>��A�� ͼh���a��'�=����/Ku=�9l>�K.>L�/���,=��=ŧ�<ߥ��)A�<9h=d�=/z=��
>���=Jd>R�?���>�a���%ٽY�������^>��>�µ>)��=v#ٽwD��"�ӽ��>�4?z��>�p�9}��/��#����>��>1\=?,�+?/�=j�8��K��`�=���@�>G�[>9)��� �&���_��d�>fΦ>��:�y�=�8�?ʅ?:H?��n>������,��]�K��=��l�ȓ�>D��>��>�Ѿl�9�����`�l��S���n��ȵ�:�>d�>nu_���U<�4:�T3=�>C�>D��=k�q���a�˔�>h��>�?���>�"�0%.�^L���?���=����e��=�	�=���=M��� Z��&b�XҘ>49߾x����f��������Ի?�~�?��??��@�E�����o<VS%>ɽ�iC��0� �[>L�>i�>��[>���:�1��=�7p�>�f>i\�\����ϽAze��d����8�M��)���+\�RwE�hf�ڂ�>�2޾��=���u��>s1����ҽ�C
�2����H�y����(����?���?�5��پ��T���.���lW=p�'���.l�LR>g����#���P���@���	�jW�褴��v�>�>����11��qM#����v�>~�3?Yw��&ڴ�>&��>~�)>�6+=-Q�%\�������
��R?t_D?��\e���F�i�>�?0k�>F�>��_�����Z��>�(%?<�9?~!޺����y����<����?pA�?	8?>󞾄KN�8N>�p���3�><�?+�>��I�=�8���Ms�>ow?�DU?�W��l��P.�%�?�?%�����>���>��>��O=�9Ѿ+�lv��T�l�>��2��8I�S޵��[��)���X?>��s>��:c�(�Y��>M|���׾�z�I����<�4��"x�>M/ ���.<�.>���=r1��Q����'����J?���?,�:?��?v�����%���;�P!1>�	�>D?�>!�5�P�`���>杠>鈸��su�Ux0� 
?�u�?%Q�??�4?�2���ѿ�撿�w����7��=D�=`�C>�{<=HG�=IL�>�]o>�Nu=<#>��>c>�x�=�R]=J�=�>u0y���.�*����,��m�`�S�#��羳�M����n�>�C��j
��Z������i7�!�ǽm������<�[K<��ڽ��x>�k6?	�?{�>�d�>K�;�˯��Q��!��.�5�[yᾜﾛ��/���@Ҿ��3���N;O+�!Qҽ�Չ�n?gt�=��1=np�>Q�(���=��>ˡ�=��=f�>=��=�S�=��D��Ʈ=��M>O>�|;>Xع>6"�<}ZC�p�y�C�������>�-A?��>�ǽYcݾ�̾�I��,�>�WC?~1�>�	�	��4�tG�>r�X}D��rZ�c|����>��?�(>��K>�GB�J,3��S%=9�L>ɠ�>[�>��-=��_����>w��>.ܾ�-=8��>.� ?#m[?p3/?s�>���>��N>�C�>�L>bH>��K>�x>�v?�~*?d�?�U�>K��=t#���=�=��#�����v�8�Y�<���J�7<a%����o�q6�<�Qn<�=��;��x��:��=��?F3"?R�>��>c+�� "\�O0���ս���=5��I�B>�:>��>�>�>�k�>�\y>#�=XԾ�������>��K=��A���k������U>>n�>o�c?>0?�w��ý���U+�=? !?��]?ڼ<?�$>�L��~��=���c���m^�!:��%�:�PUH�1��=a�=��)_?$Z2>G�����>�F>�4>kZ.������>_9H>�	�>�>=9_�u��=�O>>��="JY�.a
>e�;a;�3c��t�=y�>�������$-D=n(=��M���Z� ?��0?" ��U>X�Ž�� �:e��c�=���>�b�>���=�3��i��避�	_������K??��?c������#��=~�g�X_˽1�u>u�t>)>��:.�B�M�E���;�ð>�Q�>��>ce�=s�1��}r����Z�a>�ė=g��=卞?䛁?���W�(>��߾ɥV��P�G#+��^�=���=[D����"��.F��*��߾��v<���=g��>��?�;�Tܟ���������rY�X�ڼ<��>�$�>� >m8�G��=Gx+��6������# ���0�I�>Ӯ�=o@�>jo?8�?τV?�1?���>Te����> ��=�h�>���>?�6? ��>VY/>��O>���<�@�3�����@��m�=��ݻ�Y�=W�><�j>*�]��;�$=<�ͻ�<��	��r
=���j��)[�=T��=�~>Ӧ?�D�>��>JA<�C��/� ��:p>a�>��>��?=��>��;���k��>~F?j��>e�E�:��|I����,�>m�?�P?--,?p$�>�L;[;�('�2V��N_�>��>�f��8�Z����ɾ�� >@��>��]�=e�> �s?N�S?�N ?1+ʽ�p��?e�t��Hsm���.�f��>+h�>6ۙ=6�ľ�r8��}��HQ����*��<�I����=8>��=ݲ=��_=���=RGA=՗��r潟����FP��m�>|�>���>Q��>���=W����Ҿ?@oV>XZҾX������1;�����ܶ����>�f
��%��懖�#���� Y�C�?VM�?\yQ?3f:�3�b���<�ʼmD>��3��]�p�Y=�A�>��5>�4J�U����ފ��{1>��>^��wHH��8��ۍ�N ����k��i�'���5Q��K����X��>��<k)�=�'1�L�>?>8���\�p���¾y�ɾ�/ֽ��?]�`?��=�^z������$�{�����=�G��ڋ���o���=z���o�qV��-����𾡆 �h��bC�>�0r��j����z�=��W�=d�>�+?Չ�����7��P�=�_�>P%g>VՃ�L��	���fI��KO?k-? ���澼��C���Y?}��>�P1=�Q��GJ���`>�G?�,?�P,>"����̖�����ZD�?lD�?	�.?����a=	���=��$���v?f`1?|=�>���@����Ѿ��>��?R�K?����m���.7����>M�j?����>}i?��>܎>� ��;&���te��R�>0N�=�}���ΐ���K���y�>��>��%�ު���>��Ѿ	�	�����z�mDb���S<�}�>E����=��^>�^�=�����A����{����N?��?�=?�m%?�r���������y=���>�&�>�{�'��
�>��M>���M�r������?��?%��?3�A? ���ڱпܟ����/V���=0C�m�>_�=M=��>�R>�e>��w>]Η>=>fY�=_�=�VE>���>�y}��,�&��.t���L�~�4�P��o������ �<O$Ծu$���ƹ��l�Ð��a�˽�.^�C`o��)�}��7��>��!?HO ?��%?zn�>�M�<>{��+I��8��'�	>�VW��m���d����b�x�����:���.y��>C�\�⾎��>���=��>�?*/>�{{>��F>�bw2>AL�>@1�=̢�=a�;n�>%��>��>�S>�N�>����X���y�1]a�_¥��WH>��?ּ=
T����B����d��
��>�$2?A�>�"��%w���ud�>u�߽aւ��(׽����̅�>��>��G=�.鼭$�����9���H>�M�>x �>@�O��٦�Z�9��_�>��>�ᾣ���>c�?�A?�o)?_�=�S�><��=�^>�͘=	!�>�_�>�e�>�%?^�?5�?KR?!��=nK�ġ�=Մ}=Zz5��8�:։ݻo�=���r��;�?�<�܅=M�*>��<���=�
<��&��H�<�����>�X(?���>�k�>{��*�}�6��96����=H<ĽD��>�8�>Sl�>�?�>q;�>�VV>�ɟ=d�������>�>P&Z�-���*,����=#��>Q)T?y�:?��j=��x��(߽w�<ǯ�>�)?��.?ȷ>��==��3c���Ͽ|g/���3��&_�Z��=�'�1t=��G<���>�
>��C>�+>ś>�>|u�<J�0<��=>m=�1�>'��>B|������q�=��->9�G�'.�<Ɵ�<���:�N�����;^�9<�ґ���P�O��@�<�Ȑ2��O�<��?��?�
e��-E>)�|�"��6��7*>Y�>�o�>,��=h-m=�\1�)��\nb�!�:���B?�˒?��5�����B>0lS��َ�I{�>ƍ�>o�=5(Y�����_�{�k�H>R�>���>ks>�}�K�E��2`�a�˾��>n}�<��>O�?��p?�����ü^��6�Z����`LF��X,<���&9��B���a��=�#�o���*�����>Ɓ�?���e��=]�%��%��|ip��潭��>Al�>��>-_;�C >�K�Y�j{�k������?��=��U=A��>�/"?u%?=j?��$?4��>�U形��>I�m=�H�>���>��?���>J/�>�R>�>B���Y������۹��$�=��!��#
>��h>��<>�A�=��;<K��=�=�8=7:R;˫U<?���	�<��">_�L>{v.>hq	?cB�>lT�=II=�#��N�̼m�X>`a�:�m>hk�<�����V�׼�M�>??�!?^������_ �Mb��t>�>;��>`B?��X?�>���f�+�a��EMƾ���>�/�>k%�� 3�|�!�����]~>T��>^�S�T8>�%�? 	X?2?��w
9���\�	.�S	�<��w���>H>x�n>:�ϾP|<��΅�����~�b���<�g$��3E�='��=��Z=�",>�7=�mn>�_/>��Q=i <�O=K�׼�\>;�>Ԥ0?���>d���I*�Odž�H+?�$'��o��RO�����D�����>*�@>#`�=}��>��k$��4㤿��&�XY�>o��?���?��?I�¾�a��T��T͒<������x����}�>d	>�)�>�о>Ĩ�cE�j̄��@�>���>��)<�`���ǡ�c�8<���G��W��S�M�������Ȑ���l">\�3>�>�?���o�>_�>ą
=6y�Q�y�|���T�M�����?.�J?ܓ�mD�=ш�JN��#̾խ+�Ϟ��	�G�c"վ�;����/�`7��uґ��詾�B̾׿��9ĩ��1�>I�_��_��?d~��q'��x9�><>R�/?�%þ�3��Ж�IO~=px/>ֺ	=�$龬݊��ԙ��	�v�W?1y9?"��o4��:C�o�>�^
??��>� $>5������9�>��1?&-?�U���U��Ec��r�?��?�]??�i��9�����MK����>{S�>�?w�-��Qgо� �>4q?�Y?��Q=x�]�e�+�/�>
ܒ?����+>(>?�j�>�oZ�����C���ښ�����}R=�[!<sэ�F{���V{<��>\~�>��E����Y��>M|���׾�z�I����<�4��"x�>M/ ���.<�.>���=r1��Q����'����J?���?,�:?��?v�����%���;�P!1>�	�>D?�>!�5�P�`���>杠>鈸��su�Ux0� 
?�u�?%Q�??�4?�2���ѿ�撿�w����7��=D�=`�C>�{<=HG�=IL�>�]o>�Nu=<#>��>c>�x�=�R]=J�=�>u0y���.�*����,��m�`�S�#��羳�M����n�>�C��j
��Z������i7�!�ǽm������<�[K<��ڽ��x>�k6?	�?{�>�d�>K�;�˯��Q��!��.�5�[yᾜﾛ��/���@Ҿ��3���N;O+�!Qҽ�Չ�n?gt�=��1=np�>Q�(���=��>ˡ�=��=f�>=��=�S�=��D��Ʈ=��M>O>�|;>Xع>6"�<}ZC�p�y�C�������>�-A?��>�ǽYcݾ�̾�I��,�>�WC?~1�>�	�	��4�tG�>r�X}D��rZ�c|����>��?�(>��K>�GB�J,3��S%=9�L>ɠ�>[�>��-=��_����>w��>.ܾ�-=8��>.� ?#m[?p3/?s�>���>��N>�C�>�L>bH>��K>�x>�v?�~*?d�?�U�>K��=t#���=�=��#�����v�8�Y�<���J�7<a%����o�q6�<�Qn<�=��;��x��:��=��?F3"?R�>��>c+�� "\�O0���ս���=5��I�B>�:>��>�>�>�k�>�\y>#�=XԾ�������>��K=��A���k������U>>n�>o�c?>0?�w��ý���U+�=? !?��]?ڼ<?�$>�L��~��=���c���m^�!:��%�:�PUH�1��=a�=��)_?$Z2>G�����>�F>�4>kZ.������>_9H>�	�>�>=9_�u��=�O>>��="JY�.a
>e�;a;�3c��t�=y�>�������$-D=n(=��M���Z� ?��0?" ��U>X�Ž�� �:e��c�=���>�b�>���=�3��i��避�	_������K??��?c������#��=~�g�X_˽1�u>u�t>)>��:.�B�M�E���;�ð>�Q�>��>ce�=s�1��}r����Z�a>�ė=g��=卞?䛁?���W�(>��߾ɥV��P�G#+��^�=���=[D����"��.F��*��߾��v<���=g��>��?�;�Tܟ���������rY�X�ڼ<��>�$�>� >m8�G��=Gx+��6������# ���0�I�>Ӯ�=o@�>jo?8�?τV?�1?���>Te����> ��=�h�>���>?�6? ��>VY/>��O>���<�@�3�����@��m�=��ݻ�Y�=W�><�j>*�]��;�$=<�ͻ�<��	��r
=���j��)[�=T��=�~>Ӧ?�D�>��>JA<�C��/� ��:p>a�>��>��?=��>��;���k��>~F?j��>e�E�:��|I����,�>m�?�P?--,?p$�>�L;[;�('�2V��N_�>��>�f��8�Z����ɾ�� >@��>��]�=e�> �s?N�S?�N ?1+ʽ�p��?e�t��Hsm���.�f��>+h�>6ۙ=6�ľ�r8��}��HQ����*��<�I����=8>��=ݲ=��_=���=RGA=՗��r潟����FP��m�>|�>���>Q��>���=W����Ҿ?@oV>XZҾX������1;�����ܶ����>�f
��%��懖�#���� Y�C�?VM�?\yQ?3f:�3�b���<�ʼmD>��3��]�p�Y=�A�>��5>�4J�U����ފ��{1>��>^��wHH��8��ۍ�N ����k��i�'���5Q��K����X��>��<k)�=�'1�L�>?>8���\�p���¾y�ɾ�/ֽ��?]�`?��=�^z������$�{�����=�G��ڋ���o���=z���o�qV��-����𾡆 �h��bC�>�0r��j����z�=��W�=d�>�+?Չ�����7��P�=�_�>P%g>VՃ�L��	���fI��KO?k-? ���澼��C���Y?}��>�P1=�Q��GJ���`>�G?�,?�P,>"����̖�����ZD�?lD�?	�.?����a=	���=��$���v?f`1?|=�>���@����Ѿ��>��?R�K?����m���.7����>M�j?����>}i?��>܎>� ��;&���te��R�>0N�=�}���ΐ���K���y�>��>��%�ު���>>����~0/�="&�����X�=e��>�o����z>4a�=�z=�/��ݑ�����Qgq�X�$?���?\gp?:?��ܾ�{���1�<��%>���>�c,>x�*�<m��͊�>&��>�u�����&���b?���?���?�H?|g�����yߐ�x���J�����>�&�>����R_>]�
�8B�=�,=�>+<���>R��>k>�!�>}�|>4>c{�1&� ���~���j�jb��v5���ʾl��~;����ڽy�Q�Q9�Q����$��_�<���刻��S��g�=~W/?B=�>T&�>��d>���=���Q��*޽N$���H�H��������ƾ5�¾7 ��1x������\���-?��=�;�>l4�><�=ȤM>�ߏ=��>aD�=���<��>C��>N>,��>�\<��R>�g����> �=������x���.���:��輞�C?��7������~.��kɾ�d��W��>�	?f,x>�����sP~����>�X	��K����8�(�>Ў�><��=u�;<�&�<L����&�J\�=經>�>)�ϼ5ډ�X����=@��>*P��6b>���=8CF?Lp?��(?�9�=ٝ(>���>���>���=�8�>�˃>02�>8�?��?8?b�>V��=.�����=,�ɽ�\��f};_�B��>��E�n�=�׍��ƛ=G�=�iG��*@=�奼k���A+>!��=T%	?	�??�y�<�	&?�Ǉ= u	�H����_q<�*>&b$?yI?���>��=؞�>�>?
<|"$������>[J�>XjO�d)������	�>���>�F)?�@?5W��.�ھ�:�<���>R��>D�>?f+?��?���13���S���X¿��0����㑾�x�>`��>�}q�>�IT�6�>�d�=ش�k4�>#��>U��=pм>/ѽ���>0��>r
>�+�|�>8?;IN��=�%=quK<��= �ؼqkνf�H����0�9��h���=�e�=$k?O�?̭k<�J�t�i�|=�si��!��>�y�>���>7P�>z��=)(�p�^��zF�<_i�P�>e?�~?��H����=��ƽ3�-��|�>�7�>P��=�'o�W��������<���>�
?z�>T[����T��	c�:��F{>/�(>�@��e��?�q�?�%��0lľ�&������M���>-�Z����D۾�7Q��]�!�	��BL�&fJ>tG>D�>�jy?�羡A�>@ﵾ�`���;��*ԗ�WoG>࿧�i�V?+��>�ߙ�Rq��4���G����q����=��v>2��=���>��?q�>�jm?�	?+9�>�Q��bH�>B
)>�j�>>��>b�?�(	?�?Ƚ�>|Y�>N9�=�e��
� �v���Y=�B!��;�=
>u�L>Uױ�3#H��b=�J�=D`���`��=`9�<O�t=�u�=�t$>l�>^�?Pl?�[6�|9ʾxǻ>-RQ�,w[���=��>,�=HX�q�=�	?��?��W?a=?�d�>���b�H�ᔱ�|�ڹ�p?�q�>j�>�v���(b>��Ȉ��l]>jf>�߽p�����)��n�K�L��;>;�>5>�>h�U?�-F?�u*?���kH'�hHo����S��E}�=(�U>P=>�T�����һF������i������;=��w��=_���o=F��>cL|>G�=<��=���DJ����<�&=��>��>�C?[�&>Z�=A�ܾ�$�)�I?𗡾j�E�oо(l���>p�<>-�m�? ����}�	��C=�e��>���?���?�=d?C�C�����\>MSV>�>��.<q�>����Jc����3>,�=�|y�������;�]>Q7y>�ɽ�ʾ�/侠�H��C����Y���-:Ծ[a��_⸾_*�{ά<`W,�?������GO�0ŀ��=����J���������E�ͼ�?_-�?#!�=�T�Ũ��%h�ы�I��>!O�`���к��Ҁ�m�K<�#+��T�=.����(�/_�׼$�!b�>s�K�,w��Dl�G�H��RԾ���>F�`?TL�������7~���>�7>D���Ֆ�Ր����7Q?��;?�����νPl/<��轴��>��>��e=P7���s�=cz�=1�?v0?:�Ҿ�>��[����]����?i��?.}E?�vW��'�_,����!�>��?l�>Q7��G��u�#�,3�>4�C?'Γ>1������'���>��q?��I�LB>\�	?"�>�w���`���"C���R�<�0r>V(U���$�7f���Ѷ���j=yA�>f�e>0�1�@����� ?�ܾӃ����>�V�����=�D?l�7�q8���®������_��+����}�r�<�U:?�?j�8?�<?T��I�9�U鱾�R9>��?�Ľ=���z>)�?�f������	���?n��?"��?�R�?�>b��~ѿ�ѕ�����o5�� ��=!�i>�->"�U��o,=[>N>zu>X3c�@0�=��>�o�>\lM>.z%>l�W>X�U>n����i&�|������\16����n���m��������߸ľ�o���\�b�[��ϼ����m���۽@����hX�*�U>�-?v˸>1Nz>)J,>�^y�򚌾>��:�^���#�<���N�����幾���f��C9�����7.��c(?���=i�C=�P�>t,��?>0"�>�|�=�;%>�W�>R��B}>b�4>��J>��>���>R|�=�+�>'9)>�ڃ�\x���6(��tn��j3�KC&?���;��9x3���оS֒���>Á?2�A>�)�%����=��Te�>����iA��*��H������>N��>#���xj�+����n��r.�e�=>`�>1�>N��6�j�ђ)�a 1=�ۢ>�'ܾ��I��۔>ְJ?d�w?���>�R>I�?�6>3wH>�<>K�>��>�c5>ʨ?Q�b?�|?�[�>g�;>cs�_��=��p�G��y�=����o"=��Y���=Tf=rh>���=AH=X�)>c>=_F���%��Q��:5?!�S?�>a�>W;��;�m�d1z��w�=�Y>>��W=ER�>k;?���>|�>�>�o�UE�y�־u�龟��>p~�>��B��ޠ�z�X>Tm�>�r�=T��>W:?K�]�FhҾ�7� �>���>(�?��-?9k�>������r���qo��I�(��R8��<=R�X>�6���~�(���i$�>�7�>Y�Ͻܓ�<�:�>��>�6��-�m=2�>���=�}�>N+0>�h�:P��<}���(�E�-;�2�=�C��Z�C��Xս��T=��<�b;"��#��9��G���Q�A���)?�%?��>��>����v6e����RK
?�Q�>�$?�.�>���>ǝU���L��E���$�L�]>��u?�L�>���>�I��K�F>���>�T�Zƽ��ټ���=�L���>̳.?*?�
�>�������B���}2�v??T��=��0�]י?�"D?��������9�2z?�Z@6�������-ʾe����1���4�����#�-팾HA/>�C�>nɠ?����TJ�<ߡ��z:����h���\����Q�=�^�>h�>AD,���ؾt�K����׋��ꞔ�}�>xԆ�2**>�+�>�4J?5��?�iA?|�>x�>=�c?�ܜ>}��>�z>^�R?�-�>@af>Z1>���>�Y���>q�3��8����=¶�=��Q��ڼ�ж=�a>� �M"��������������	b��i�;;Y<><�>��>×?��Q?:J�Q���9��w��=��\>8o/��L�<3�&���T��$o�>�-?��?�`?z	�cl=�%�2�t����t�=��W?�E?���>5�>�ؘ=�圾<X��4�>�H>��r:`���������@��p%!>}A�>.W�=+��>꤄?��!?�?�ݽcK�?�~����J%������!s}>{[�>��¼g�߾��5����������5�$�g9��P���>=�	�=/�����`>;r>�@�=+���r�Z���ka�;]5�>N&�>���>7R>���<�Ҿ���>xb?����ʾ;jξdcE�tzg�ҩ�>�V�>�,Ѿ�9>���ij��FA���$O����>���?�ǿ?�s?��E���?��m>��½N�=�bP��1�w����t½��>���=����tȡ���>�?s��>���Fܾ������#=<����@^�,I�V$����c��*׾�K����=�P�����=9}����	�H܇�C�#���8���,�C��T�}�k#O�m�?�}?W#��#}�<a^(�e�[�v��q�>�7�+0��efǾ���'��=Ծ�{��t�ھ�(�i����>��b�J���>~�$�/���dSB>��'?�ξ!Iо:M%�*����4>;��=?����%��
̕��>����^?��3?��R�Ѿ�n����3>�0?�>���=�ϟ����05�>��5?uQ8?F �<�ٌ�P�����;���?w�?�}@?tP�F�A�������y�?��
?S�>�D��rlѾ�s�oL?d�9?���>ܪ�����l�>��\?�N�'�b>b
�>c��>A�����L������q��\�5>�#�!����`�]�9�Ҡ=�Ԟ>��s>e�\��t����>>����~0/�="&�����X�=e��>�o����z>4a�=�z=�/��ݑ�����Qgq�X�$?���?\gp?:?��ܾ�{���1�<��%>���>�c,>x�*�<m��͊�>&��>�u�����&���b?���?���?�H?|g�����yߐ�x���J�����>�&�>����R_>]�
�8B�=�,=�>+<���>R��>k>�!�>}�|>4>c{�1&� ���~���j�jb��v5���ʾl��~;����ڽy�Q�Q9�Q����$��_�<���刻��S��g�=~W/?B=�>T&�>��d>���=���Q��*޽N$���H�H��������ƾ5�¾7 ��1x������\���-?��=�;�>l4�><�=ȤM>�ߏ=��>aD�=���<��>C��>N>,��>�\<��R>�g����> �=������x���.���:��輞�C?��7������~.��kɾ�d��W��>�	?f,x>�����sP~����>�X	��K����8�(�>Ў�><��=u�;<�&�<L����&�J\�=經>�>)�ϼ5ډ�X����=@��>*P��6b>���=8CF?Lp?��(?�9�=ٝ(>���>���>���=�8�>�˃>02�>8�?��?8?b�>V��=.�����=,�ɽ�\��f};_�B��>��E�n�=�׍��ƛ=G�=�iG��*@=�奼k���A+>!��=T%	?	�??�y�<�	&?�Ǉ= u	�H����_q<�*>&b$?yI?���>��=؞�>�>?
<|"$������>[J�>XjO�d)������	�>���>�F)?�@?5W��.�ھ�:�<���>R��>D�>?f+?��?���13���S���X¿��0����㑾�x�>`��>�}q�>�IT�6�>�d�=ش�k4�>#��>U��=pм>/ѽ���>0��>r
>�+�|�>8?;IN��=�%=quK<��= �ؼqkνf�H����0�9��h���=�e�=$k?O�?̭k<�J�t�i�|=�si��!��>�y�>���>7P�>z��=)(�p�^��zF�<_i�P�>e?�~?��H����=��ƽ3�-��|�>�7�>P��=�'o�W��������<���>�
?z�>T[����T��	c�:��F{>/�(>�@��e��?�q�?�%��0lľ�&������M���>-�Z����D۾�7Q��]�!�	��BL�&fJ>tG>D�>�jy?�羡A�>@ﵾ�`���;��*ԗ�WoG>࿧�i�V?+��>�ߙ�Rq��4���G����q����=��v>2��=���>��?q�>�jm?�	?+9�>�Q��bH�>B
)>�j�>>��>b�?�(	?�?Ƚ�>|Y�>N9�=�e��
� �v���Y=�B!��;�=
>u�L>Uױ�3#H��b=�J�=D`���`��=`9�<O�t=�u�=�t$>l�>^�?Pl?�[6�|9ʾxǻ>-RQ�,w[���=��>,�=HX�q�=�	?��?��W?a=?�d�>���b�H�ᔱ�|�ڹ�p?�q�>j�>�v���(b>��Ȉ��l]>jf>�߽p�����)��n�K�L��;>;�>5>�>h�U?�-F?�u*?���kH'�hHo����S��E}�=(�U>P=>�T�����һF������i������;=��w��=_���o=F��>cL|>G�=<��=���DJ����<�&=��>��>�C?[�&>Z�=A�ܾ�$�)�I?𗡾j�E�oо(l���>p�<>-�m�? ����}�	��C=�e��>���?���?�=d?C�C�����\>MSV>�>��.<q�>����Jc����3>,�=�|y�������;�]>Q7y>�ɽ�ʾ�/侠�H��C����Y���-:Ծ[a��_⸾_*�{ά<`W,�?������GO�0ŀ��=����J���������E�ͼ�?_-�?#!�=�T�Ũ��%h�ы�I��>!O�`���к��Ҁ�m�K<�#+��T�=.����(�/_�׼$�!b�>s�K�,w��Dl�G�H��RԾ���>F�`?TL�������7~���>�7>D���Ֆ�Ր����7Q?��;?�����νPl/<��轴��>��>��e=P7���s�=cz�=1�?v0?:�Ҿ�>��[����]����?i��?.}E?�vW��'�_,����!�>��?l�>Q7��G��u�#�,3�>4�C?'Γ>1������'���>��q?��I�LB>\�	?"�>�w���`���"C���R�<�0r>V(U���$�7f���Ѷ���j=yA�>f�e>0�1�@����[�>��ƾ��a��L[�^��XH�,�=0�>�ɾ����.>8�=?-�Gk��Eځ�����N6?ݢ?��9?T8?����'ɾs�>��ǽ�?�>�� >E�.=fv�>��>��"��#^�>��LH?��?E�?��`?N>I�AGӿ��+���������=!%�=��>>��޽�ɭ=��K=�Ø��W=�w�>l��>o>;x>n�T>͛<>z�.>g�����#��ʤ�,ْ��[B�� ���wg��{	��y�����ȴ���H�������#Г�y�G�e���T>�M�i��Y=�I?1�?��->�A?�wp=�3�����G��q�"�ß����)ҾrPC�Q����'�=?=��L��F�b�ў&�5��>�q�=*c����>B�P����=�>V�.��K>Xŀ>��>o.>��N>��:>$�=�41>�I/>���>A�=F���ك�dr<��^���s>��3?7�X�iѐ��(�j޾���xBa>���>�G>n�$�󳎿"�d�k�>LpU��u���p��8/���c>`��>��=q���wÓ�$�)�n�>�c�>0u>��<�<l����[S>8 �>&վW >
_�>��!?#�y?��0?�!�=�κ>#kb>�8�>���=l�=>:�M>�Ќ>a�?D�:?:C/?
��>嚵=�u�ۯ=Ҕ(='K�N'u��Ͻ�����#Z���߼]^=GH�=���<�)�=�M=4�#��򅺝�&=�Z?m?,��>W�?�� =Z�����.�jZ���R���C����>M�[==:?'�K?e�>j	>�b��N��|�Ʀ�>��=(E��78��Ĺ��X�=�A�>t́? ?WrF���
�ю��n]��>�/�>%�@?��>R�?<l�������˿�0�#E(��+��j�=�s6� y��G�>�/�>��l>-�=?,�=��W;y�:>��8=�ʺ=��g=e���E>�>Y(���[�<��|>��4��[8=����=�c=�R<`�v�x� ;�2{����J�e���h<L�<>�h�G���?��L?%J��&0�������.��<_�H?O�3?H��>y�C?t��>����*~����7��<λ>	/�?m��>z�`�7�X>�Dٽ<��rT?E�>��)�e>��s= %���iS��3?j8)?��w>u���7������@� ��-�>\'�=����%�?;�h?A�������e�(h[��v������b罣*��	榾W���K�����8:�ѿs>1��>�KZ?c�����=�ݽl��y����߾�E5�W�4��"?���5k>,L�=�!��e��B˾���=�!?�փ=���>� ?�?��b?�q?��?�;�?��=���>�<�>�?- ?!X�>��~>�>a� =��.�y��pŊ�}�<v������=��>0�'>��d<s�"=z@4=���<��>�6O���{�<5�7<�=c�=��=T�>�?�2�>`E1�3�^>�4V��l����o>���<4=?��� ��Ծܹ�@`�=*�?�/A?L[?�e7>w�ھkP���Q���5>�/S?VU?�S�>�+=�A���C'�;W>kf��ps>����E"��C��N������>�`�>)�Խ�\�>���?�#?�C�>�U�>����hW�!	��l����/=n�>���>Y	�>����>I�z�����P)2���L>���>nJ>�j�"� ���F>��J>qq�>��� ��,p>�/<��:���>y��>j$?�H}>UU>i��t�2�� ;?�=���	�Q�y��'����=s��>���>��g:��>Y̽�r��;���X1����>M��?Z��?�l?�^��*" ��i:����>y�:$�8�Q��� �p>n�k>�:D>y�}>͠�*B��on�=R>>��>���8R���T g�/�/=�ி)&R�_#Ǿ����(�5�پ�ڶ�
���f
��G��|͒���׼*0��0;�H�:����ް���̾��ľ���?Z۝?���ƫ���,�t�0����W���w��~�������j$�ϫþ%���Ӿ!��ٹ4��#���/_�>��X������5}�V�&�X��-68>G�,?�rǾ+˸�����t=l�#>���<�T��a֚�^��V?>;?
�羇����s�'>Ǹ?b��>s�$>���������B�>D`0?r�,?�X�9��%����R���?���?�j:?I�����1�[~��z׼;��>j��>= �>Ww��(�ʾ�tؽ~+
?�cA?l�>���Q͉���(�;e�>Z0`?�pm��ˀ>0�>Z?�>@ώI�r����<6��K5��f�>��;��C�JM=��h�w��=Bt�>�<~>|���}���� ?�ܾӃ����>�V�����=�D?l�7�q8���®������_��+����}�r�<�U:?�?j�8?�<?T��I�9�U鱾�R9>��?�Ľ=���z>)�?�f������	���?n��?"��?�R�?�>b��~ѿ�ѕ�����o5�� ��=!�i>�->"�U��o,=[>N>zu>X3c�@0�=��>�o�>\lM>.z%>l�W>X�U>n����i&�|������\16����n���m��������߸ľ�o���\�b�[��ϼ����m���۽@����hX�*�U>�-?v˸>1Nz>)J,>�^y�򚌾>��:�^���#�<���N�����幾���f��C9�����7.��c(?���=i�C=�P�>t,��?>0"�>�|�=�;%>�W�>R��B}>b�4>��J>��>���>R|�=�+�>'9)>�ڃ�\x���6(��tn��j3�KC&?���;��9x3���оS֒���>Á?2�A>�)�%����=��Te�>����iA��*��H������>N��>#���xj�+����n��r.�e�=>`�>1�>N��6�j�ђ)�a 1=�ۢ>�'ܾ��I��۔>ְJ?d�w?���>�R>I�?�6>3wH>�<>K�>��>�c5>ʨ?Q�b?�|?�[�>g�;>cs�_��=��p�G��y�=����o"=��Y���=Tf=rh>���=AH=X�)>c>=_F���%��Q��:5?!�S?�>a�>W;��;�m�d1z��w�=�Y>>��W=ER�>k;?���>|�>�>�o�UE�y�־u�龟��>p~�>��B��ޠ�z�X>Tm�>�r�=T��>W:?K�]�FhҾ�7� �>���>(�?��-?9k�>������r���qo��I�(��R8��<=R�X>�6���~�(���i$�>�7�>Y�Ͻܓ�<�:�>��>�6��-�m=2�>���=�}�>N+0>�h�:P��<}���(�E�-;�2�=�C��Z�C��Xս��T=��<�b;"��#��9��G���Q�A���)?�%?��>��>����v6e����RK
?�Q�>�$?�.�>���>ǝU���L��E���$�L�]>��u?�L�>���>�I��K�F>���>�T�Zƽ��ټ���=�L���>̳.?*?�
�>�������B���}2�v??T��=��0�]י?�"D?��������9�2z?�Z@6�������-ʾe����1���4�����#�-팾HA/>�C�>nɠ?����TJ�<ߡ��z:����h���\����Q�=�^�>h�>AD,���ؾt�K����׋��ꞔ�}�>xԆ�2**>�+�>�4J?5��?�iA?|�>x�>=�c?�ܜ>}��>�z>^�R?�-�>@af>Z1>���>�Y���>q�3��8����=¶�=��Q��ڼ�ж=�a>� �M"��������������	b��i�;;Y<><�>��>×?��Q?:J�Q���9��w��=��\>8o/��L�<3�&���T��$o�>�-?��?�`?z	�cl=�%�2�t����t�=��W?�E?���>5�>�ؘ=�圾<X��4�>�H>��r:`���������@��p%!>}A�>.W�=+��>꤄?��!?�?�ݽcK�?�~����J%������!s}>{[�>��¼g�߾��5����������5�$�g9��P���>=�	�=/�����`>;r>�@�=+���r�Z���ka�;]5�>N&�>���>7R>���<�Ҿ���>xb?����ʾ;jξdcE�tzg�ҩ�>�V�>�,Ѿ�9>���ij��FA���$O����>���?�ǿ?�s?��E���?��m>��½N�=�bP��1�w����t½��>���=����tȡ���>�?s��>���Fܾ������#=<����@^�,I�V$����c��*׾�K����=�P�����=9}����	�H܇�C�#���8���,�C��T�}�k#O�m�?�}?W#��#}�<a^(�e�[�v��q�>�7�+0��efǾ���'��=Ծ�{��t�ھ�(�i����>��b�J���>~�$�/���dSB>��'?�ξ!Iо:M%�*����4>;��=?����%��
̕��>����^?��3?��R�Ѿ�n����3>�0?�>���=�ϟ����05�>��5?uQ8?F �<�ٌ�P�����;���?w�?�}@?tP�F�A�������y�?��
?S�>�D��rlѾ�s�oL?d�9?���>ܪ�����l�>��\?�N�'�b>b
�>c��>A�����L������q��\�5>�#�!����`�]�9�Ҡ=�Ԟ>��s>e�\��t�����>H*�JlN���G�2�������<�<?7󾚟
>�g>�>��(��猿�i�����2L?�H�?aSS?ƃ8?Y����0ﾻP���=�;�>k��>��=j��eq�>���>h�/s�`<��y?u��?�n�?̈Y?f�m�7?���F������`-���[�Z�=�nY>��9�AN"=#�<�6�=e��=*�>��>�>�n=>��>���>� �>��~��>��E��:���) 7��a"��8��
ؽ�d���4���!��t:�d���vA�����O� n��������=���� (9>�>qU�>�ZP>�c�>w�>֊T�5��WO�� �"��#'�9~��wо����t��u��Y��Ay���w��Qj��{�>蛩=DO>���>�ኽMk>v�>l�L=1�B>/*><=�=��+>�s>�xs>Fjv>��g>�n�J�>��=�I���9}����p��
<�;C�4?�տ���m�KL,��餾q�۾~�
>)#*?��\> �4������WV�>gw��~7ξ��E�}�E��F�>�κ>	4�<o����̾#�n7rk���e>塢=��=|��.�־����"н���>	�����=y��>�|?C?QC;?���=Jp?��>*2�><:>R��>��J>M2�>�%I?;R??�p=?�>: >.O���)�<�n�>����A�O�½{%�<�位h!>إ����=��>�)��ռj�ƽ&�=�k�='^���>�>?�?m?���Nj��t��_ҫ>/�n����>�"�>�mO?i4?�0?�Q�>�r->���8۾S>���=�2O��$��T�>G�>��R>]
*?��U?���SP7��3(>��h>�3�>�z?�I?� ?ػ�>}�U>�����ƿ"签S�����>.�c<�no����>xe�ٟ�>�LҾ� �>XD��Be>��y�HС=(cY>+P>]]�>��>�>�"�=�R>u�>�<R�+��=6*�>TU���>v漽=�J>aO�^q��^6��fR=�K���������?%?����P�=�{Q��x�ֹ���c�>uT�>'��>̩?=:	>�ȾQ_D���*������?On?m?�>� �ǩ=� l=�$�<,/�>�3�>���=�S��j�Q4����d�d0�>�w!?A��>�Ҿ��;j�%�n�"3�⿑>�η=�kV��T{?g8?��ݾ~*�'�_�2�w�P�q���O߾�����5�+Y�24���;�D��q��5c�>⑾?"[�]��㧾�����������S>N\*�_>�<H���������[;�'�'��s���6��ڙ>>U��>=�*?�.?l0u?�8?�?��h��=?���=���>�}�>,+?D;A?f�>o��>�`?� �>O>>a�޽r6~��� �J���{<KFo>��>�7�=&�o=�>�R�=lν5<K�$�S=���oԻ��<��>s��<X�?�k?� ���r�=�D�;	��j|�=3��=)�>���+Kݽ��D� j�>K��>�5? 	?�>Z�����߾�iھ$2#='5�>��-?���>���$p=�;޾�	f�!��=��>)2���.w�@V��R����ݽ�ӡ>�*�>��>��>B�?��V?�hL>�eھsm�A�^��e��3�"�۾�B~>�h���)'�ܪ��nr����Q�X6���-�;���b=��f>��#>�Z�=�>�i5>���<X����D���I�>b�=>�K�>�]?P>?4�>�>p>�q���	����G?|-�����m���;r;��]�>D�>>
;	��?'���5~�UD����<��_�>�a�?���?k�^?i8V�/���? t>I
P>Q�>F��<I�]��~����Ž�q?>��=@c���8��c.��R�A>)E>@��o���w��)+��Q��bZ�1�	�8������#��U۾x5�>WKm�Q��>�9��[;��ؾ��l�]�<�����~�̷���숾β�?�T�?*J�N�e�~�)�W�5��*&�[��� ���H�<���;D��<Nо�h��%�����U�4��x%��F�>�?E��W�����3�#��q{���=�=	?Cz �4;_�3��Q��=0.)�rYK�k4ξ~���MY����&�o�"?�P?�޾$U��!7��%2=�?/��>:��q֖���<�+�>�4�>�0?��3�U���ю�����UY�?в�?��P?]�Ǉ@�t�*��8߾<��>�k?v�>D*
�1eZ�2&߽�o�>9��>�&-�ԃ�iŊ���Z����>�m? ������>b�?\��>WT־�ꇾ%�)>��۾)ֽ���=��ɻ'�I��8������&�ۺ�>�R>�����z�&k�>?���'�H��D�L�޾{�)�H�Ѽ��?����l>��>�`$>IM@�����c!|�����>?�|�?��B?.)>?�uǾ��ܾy5��5r<A_�>��N>L��;"޽<E�>���>	� ���v�r	�X2?�m�?���?��B?�}�H�տ�c��PԾ1DﾫI=w{>s](>'�=E�>�>I���$��=_�>F�>ߜD>ѯn>���>ڟ>��+>�ބ�b ��e��ME��eu/����(��8�e?��|�H�ȩ4��Zj�)Ex������w<����E�����Y�C<�I���] >`�>B�>�t]>�>t0>��V����l��i�X�~վBz澰	��҅V�f���(���0��?�u���:�>Ig=��>���>�5�j[B>�u�>�!�=8�6>� U>F>�HI>��l>mA>�2>.�}>���=Є�>�W>�����s��@���$�=GL��
�>��oi�����=徫);��i;�%�=
�=�K�����󰜿�7�>���=�<��d=$�)$4>>|�>�w[�Dg�ӗ���v�0�	��g�>��=��#�ݽ����#��SV���>'���݅>���>p�>QO�?��d?�= ?Zc��]�>V[���x>`R>�e�=��3?�V?�v{?Ē4?�d:=�x#��艽�Go�����:xk=��7��5;1��*�=��ݺ�J�;�9eJ�7A��8�ν�� >��3=&h/�،�>�HG?��?pS
?��x�+�+���?�þ�ٌ=�����?�ˡ>�J�>'�?�$�>�A�>y.�=����.k�ˁR>8�>b&q�4��h@�=r$>EW�>_�?��Z?��~���=��=�@���>
�?нP?�W�>�<�>Q�>���I�Կ3���u�{>�u+�.�"��K�>(8�w��>����*w�>Z��V�r�ʇ�>�o�=Q!\>�[�<>�n>��> �=z�<}�E>rk>�S�;<�H=U�=K�}���=����[_=�U��I=���=�^��og�Ҕ�<�=rD?�;?����r�UFf������ا���>��>	��>�~�>���=C���8R��U=��a8����>�i?7 ?(�6���=�ON����;�ʶ>�t�> �>�&=����E����r<Ph�>��?�K�>�����W��so���
��.�>���=�T��Ll�?�K?���}�սE�
��4�����S��E<Uv����ؾ!�e�A[�2��\� ��@�uӚ=���>z�?���=R_�=�n���ch��o?$��45>cc�4xq>�F������+(��/7��P,��ظ���q��`C>�ZI>ʿ�>u�?�j'?��?y�?�5?�l���+?���R.�>qŌ>:l2?��?���>],�>�O�>%1w>є/>�~�J����n>���=���<�&�>��>��q�q/F��3>���:�����ɽ(���F6����%=�Y�=�KF>��>��?�?����?��mؽ���zr=~6�=��D>1Q��)aŽ�%���f>�/�>b�+?�U�>�֒=�Ͼp��'s���ǹ��?��9? ��>���=��=�y���yR��j=��->nǊ�������5��<Ƿ����>��>�G>�D�>�ˑ?��i?l�?�����^s�����=�0����>L����r�>�>��/�����_x���)P�łI�<�/���=��=�R�=r{�>��>��=�2�,4�=/k&>n�>�T�>�H?ar?��?���>H�[>s+��$�ҾY0@?�㡾#{��ĳ�:��0 ƽ)49obG>/���#?��\�q�� ��]�A����>2�?��?-�J?wa�����=�>���=*�D=Jd�ω����Q����N>J(�:�H���#���m�=� *>(P>ؿ��m羍��ઽ�A��~�F�3��#˾��H>��������9�>�}��.?�>(	0���v>�5ξ�N��ܦ	>e��&�e�u��_L�"�?E,g?��>I�/ל�5��+�^������k�v<�)����'� ��j�
3���J�	�꾌Q��v�ɉ�>HW{��(���Jr��M!�����;�=�N/?����U���{��ۊ<���=Q ��W�Ǿ4b}��\��;�5�T�&?[7?<���K{�<q>p?��>Z(>�GɾoA�bk�>�,?�N
?�(�岓���������B�?��?��>?��X�|�@�hs�ڜ6�;�?�2
?/��>�<��d
ѾN0׽$?��/?�P�>_��I�������>�N?��K��!{>��>'R�><ؽ^��B���YM��S��M32>-��9mU�p�o�"�T�0S=�{�>�e>�/N�UV���v�>�S��IN���H�|�	����&��<��>S����m>Âc>��>�Q'�V����Q�����`�I?�|�?ŧT?��5?x����澎��@�~=oT�>�ϭ>A�=�	�1u�>���>��澥kr��H���?���?���?^�W?��l�#0׿;ۡ�������ܾj5�=��X>cQ>��=L�=��<Q(��J�k��Q>诱>�/�>�>�m>���=SRs>Q���j�$�Ț�L!��o�4����Wh��/޽h���!�{����+�t-���j�;�٤��ٽi]F��P8=�gJ�$Ԉ>��>�.�>W>�8�>��>y#��C��F}���j�n�>���������Z��_)���o����=N�=�#�a��@��>o��4�>b�>���!��>̽�>#�=Ŝ�>��>�S�=�u�>�X�>ݻ�=^{g>G>���<0j�>:��=;�������Ώq�bC��<M?;��@�>�@���`�ľ��Ľ2�?��z>ֺV�����1�� ?
?�@�ۣݾ�uS��B��p<>dW�>���=&b���z�*S#=��K������>BX>�J߽����j��G_=b��>����w�<-u�>6ѹ>r�R?|3X?]>�?��1>Q��>_� >�M<?��>��>��?/�B?B??F��>���=�b(��G������GK�����a�=/��;���;���Қ	>(��/x*�`�^>.n!>F����<��=}v�>1W?��?%g?�J�=�u��pO��y���E�>oq�=`�)?���>|?C�?��$?��>"p�>�h���&��>�>��#>L�S���s�YW�>1��>��4��YB?�)G?�G�Ҿj�=�)>!W>�L�>̣	?��>�G�=� M>Z���B�Ͽ���g�����>|��=��9�H�}>\K�
3�>/�Ͼ�=�>�/>uj�>N��>E`>�k�>j��=�aW>��>��=�?>�0"�g�8;��">���=��=�R�$`�<�q���#�=�=��=��{�A*m�tU���9=m#3�Y8?��?"��=���<��ʾ������A�\�=�:>��f>;d�>�F�+"�&�V�H�`�� ��B�p>�ej?kY?�A���jV>�䨽�L=�U�>+�?�V^>���%���3�|ø=A2�>��?���>0�ؽX:��la���(��ox> ��=���c��?�&P?�uپ)�Ѿ�n�n�2�|�*�
������V���C�����J�o �����m2�}�Y>�B�>��??�<Gi$>�Ny����դ��E$���Լp%�z��<��Y�ס��b����%1�����H[��գ���>��=�\4>��?�?F?�?9�=?תL�	$?��=��?�i�>��?�Z?6�>�n�>6�>����/�-7]��f�&:��J1=a������=�n2>��Y>;�K��j�<���=\E>=���a������ɽ1ޤ=v�V>z?�=��>�<?�@=���>sj)=e���vZ= �	=�?�4��*;�;X�w� ?'�>a]0?� &?t3�>p�ھ� �2���K���%?�;?fP�>ߎ!=r��>v��f�����=ׁ>�;½��lQ��䂾Ò��z��>���>Ҩ��ܐ>��?��;?���>-�y�<4$��WN�u�?�$�7���ꤱ=rT��������$a���~��6P��K��[�=��1�zv���Ԇ�'�>-�����W�^>Zj�=��$>%�=���>�=>�@�>�z>�71?Z�>�WN>A���-�	�I?�����c�	ݠ�'zо�>���>{�<>l����?���9�}�����>=�k��>���?���? ;d?V�C��>���\>9SV>��>ג1<��>�Z��_��0�3>���=\Sy���#�;�]>�Oy>�ɽ;�ʾi:侕�H�k��� *U�����r��>O`�3N���>�Ǐ��g>� 5�Rwu>!Q�=L<D�*�>���f����Ǿ3ݔ?���?���풽��QF�(|����7����{"���Ͼ?����Ѿ��;��������°Y�M�.�l���	?��������x�����Si/>��)>,?0� �R�$��0��)ꆽ��ս9�C�~�����8򴿪�<��3?�V+?�o��i�RD�=�����?v�?­�,����z=�w$>��>/cT?�&>P�������7Y>��?�'�?�^?����13�&:�� �yk�>`i$?�`>�� ��%3��^@����>:?ƫ�	>�B���%+�aZ?pax?6 �����>9�5?�P�>b��F�q�=+���Ǽg�=�
	����Tƞ�c���S�=H�>�y�>�j�o��Q��>�&�%%O�zC�����,����<	��>�v���w�=,d>B��=H-*��o����8����B?U%�?�jS?�F/?l꾖�����f�=�6�>�y�>�a�=/���q�>��>�ܾ��g������?�x�?1��?10V?�h��Lſy����X��<�ɾԖD>�Ʊ=ש%>Gn�=�]2>��=x;=�e�=�!�>#��>۴�>N��>�Ő>�0>@>���[ �k(���ȕ����]��Be�d���$4���W��w�}�����,n =L,ڼK��2Y����ĽQA��Z����t�=&�>�T�>���>�>���=����� �����4þW淾�O���龩�����d�d�-��l��e���F�rr���>ߙ��-m>X��>H�����=G-�>ٽ+>$r>?`)>���=Pp>��Q>)�n>�܈>��4>��K=\~,>18����e�sr��M���#��o��@cS?߼��c�+�b�V�'��ֲ�B=>2�?՞f>-Y2����a�{���?՚ռCȾ���[�;�G>^�>rYB��:<��<�a=�NX��_�=՘>�$:��f;����Ľ�>�t�>G���V>Diq>�ˊ>kx�?(�c?I:^=�@�>mE�>��?����n��>���>�>IR?�8K?+�%?�?�>N�=�{Ѿrȼ;�<16нV���Y���=u��G<��|�=���Gq%>�E}=�A =
&>�7}��ڽ~��=�/;f�>�K?�?ұ?�tb�gX����2����m�>��=�0!?�6?��[?��0?��?�b�>�D�=�ٽ���/�{��>��)>�77�ck����=��S>C�.�k?V�I? D��*�p��:�v>�^U�>�:?p0D?��>�G�=D=����ؿ7JF�pY<�`(�S}=��T�<E��<���T�8�Z��%�̼\ s>���>��>��>]�>S>1�+>6��>֛�>�%>p�ӽ��޽~�<<}D�=�5�*���3!�L�'= U�e#�=v�����,~��4�V�0� <f?��?���B4�V�־"۾��>��>8/>L#�>X��>�҂�"���?r���Q��H��H^�>�o?�?���eA>�����b�R�?��?�?�>M� >WS�d���&|>�'�>�0?J�?s ��^�!�����4�Uq�>>�='�<ip�?̗S?�?�0i��r@��O?��� ƽ����!<���ϼ��u���:�)�������H>S;�>���?<��&>U��j���삿������Ծ��X>�0>��ؾz�Ⱦ��2�g�߾�������y>�1�=���>�+<?��X?��?0'?��;?[Q����J?��`>�R;?��+>n�?\�B?=/"?"&-?��7?���Z��a��[^����=H;�=k =�}�>,*�>	�I��,�1>U��=U�ɽ[��p���o�x^n�?�:�3.�=�>�?��&?�R���P`:���y��Y=ܥ�=��{>�$*���0�g�<o>s>��?��/?���>̆�=1�ھR��آ��Q&�=̜?zi5?h��>��<�2�=4D��m�����=��k>lA`���|��־�\���%��.W�>Ԭ~>,�=�en>4�?д:?m��>L���Ƃ⾼	?���O�#L>��B�?�Y;G��,�.8��]A��}����:�5 ��O=�!
��:<L�q��A>a7X=?޻�#|>�)Ž鼋>��>��9>�A.>��>m^�>g�,?�أ>�)>��j� �,�w�I?����-i��렾�oо3U���>n�<>N��?R��2�}��
���F=����>���?���?�<d?��C��&�I�\>IV>��>�5/<��>��7���3>�=�sy�v���$�;E]>�Ky>r�ɽ��ʾ�0��H�J����fI��ｖJ+�!˪����,�־@�>+%����=��-�^;	>�������S�=�������M�-�޾�Ǎ?�pn?LS>�~l=�Ac��(���&HH>+G��Kg=�k!��D佤:�����(��:˾	�)��>I�)�R�?v����=��N!��T�V� �+���-�i�?�l��\�<H20�c^�=s=�4ꐾ�侵ox�Q@��Qo�b?8�H?�����O�8�Iܞ<�`#?�?��3=K���A����>��>zn�>�<���	¤��*[>G�?��?	�j?a-����X�#O��9\�>4A�>YL�>��+�2�d�󏾋D=�d�>�^@�~�*��\���^F�și?
��?m莾���>��?b��>$O
������r=�x����e��ޣ�4������:Y��ڻ���y ��\�>�"½���/�þOM�>X����N�v�H��X��R���<�?mL���8>P2h>��>U7(��,��0Ɖ������K?���?��S?��7?b]���4������G�=_3�>_��>�K�=�
��'�>���>8I���q�F��<�?��?�{�?��Y?hm�P�Ͽ�똿��ͭƾ�j�=�~5>$�>�/;��zA>Ѧ�<��=��!��c4>���>��>�4�>��>�r>|� >�h��|�"�/������<�(g�'�q���~S�gGy��a�%%��:%ؾI}����'�Փ��m���
�����:p�p>D�?��>��>� z>���=	���Fྖ&�k���������J���]�v�V(ܽ6�k�-��آ��Q������>Y=+�j>{�>����|�=��>�!�u>��L>�KF>D�(>�2�=�� >�[>�>��e=!�d>���<�O��lqz���	�[��k��WF?xw��T9�uM��Z���ӾO�>��?}�D>?1:�Y�����~���>�bK<9<��>
�<�+�O.i>��>�#>�I���=��9����ѽ�d¹���=Um�=T�F�=�ʾe����>�=��r>s���.$�ާ�=c/+?�rd?K8?{�8>��=�s>�;%>��]>���>�E>uٗ>���>��"?�81?�?b�>Hþ�_�>(~>J�.��3T��쟼f�/��2�=K1t�ńN�_E����F��?�=ic�=j�!>�Ƽ���?@=?ͽ??�?�����i���Q�����|�=�A|=�+"?s��>O��>�7	?��?\j�>F��=���H=���>��6>-MI�g����|�>�'�>�L=;z{?�[n?6��d畾qX6>���=8�?�<?�{C?��!?��>���9)���п.�(�{�7�4�=2k�;�,#>�q>Q�k=�d=�y�Cf>��v�>S�>��>
�z>8�P>� >6�?#1>�)Z=iC/>�x2>�4�;<�Q�>�+;�#�	>����>�(��UX�𫨽���"���
�➽�Y?�!?�Ŗ�{��� ۾��8�T���h=��z>'��>�?�l���d׾_<Y��]F��,T��=v>��l?ݻ ?a+ɾ�2>*�4�:��С?���>�6�>gP*>�λ2�	�
N�>Sl�>�?��?Y�(��6T��s,�5��y��>8.�=���'�?ޥV?f`��s+#�3�]�<�sL�7�2�\�=��¾N�;�g�LV����4���,��&~*>��>;ڨ?l��8�=�p_�CC��2G���x��ꆀ>M�����>Cz]>jv��X��6�wc��ϕ�������>�@�=�]�>� ?}?ɸd?��)?�"?�*!���.?��=��?Ye�>a*?u�#?�W?��>�?���=	���pP$��=���I�= 蟼8_�=H�[>�S>gү�!����h;�[�=xŽ�������6��<#��<z΄=���=��I>.,?OM7?�n�=m��<[�=��A�Ŀ߽��y>��?o?�=�X�z!�=.a�>$�&?�D9?&�-?	��>�Ă��N������ =�v�>؞"?��>]e>�w>��=0��q�<'�>]�2=�r'�v^��+����ǽ��>[Ҝ>ڨ�>���>�c{?ļC? B?3ℾg?ؾ�:]��C�`$>�$����=���Vb>�x$��t��tj����6Y�#✼�{�<ю�%�V=x��>�4�*{ֽ'�>}�!�EU���>�8=�@8��+�>��>h�?=�/>h	��ǘ��L,��nI?�U��a~�����ξ��&��@>/�=>"����?�����|�Y西��<��s�>9\�?���?�d?�'D�Ft��^>FOW>e�>�|(<�?�d��II��uU2>4W�=�oy�3��AF�;]	_>��x>�ɽ�˾B7�:�O�b���/]�׀����;�.>���u��66[>���ث>H�6�D�>�罾\s�=д�=��Z=[�r��ʾ��ξB*�?} t?�'�<���������h�s���������Ů��g�j�Hi���o���&#��~a��`C�ީ�?z�>"<\�c����r�P		�����~P$?wU��H�+���y�=�,����'��N������OB<"�?@7*?�?�g+���娽��S�_@?D?�b��J;���f��>�d�>�]?�O���'��������;���?eq�?�#D?C+:���=�#7����?#?���=���T��|½+�W>�,?���bS&�2�}���7�1�8?��}?mu�8�o>7�.?�ϥ>dۂ��w߽���=0�ɾL��<p�>J�-<uQ�셵;�?L��J>��?�О>�������~.�>�!����q�%W��{����4��}˽�A?['��O>ѽf�n>�s�>d0�GO��������X�W@?���?��?��J?�xپ���}2>zK��R�>U��>����a��Z>ǐ?��
����C�f��>���?Z�?�7'?ӿ��
MԿ�����pľ�M徻{>F?�:B~>���M��=�>El�#�}��⺍�>�A�>���>���>NO�= ��>�����%����yIP���!�w� ��a�\Y
��Ǚ��0�~GԾ�ξ$%�\�=T��=%:�����*�DY�@D�=���>Y_�>��?eW�>��V> �"�*�P�8�iDy<V��<ɾ�徸[7�T�7���߲�������ok���!�uL0?��==<=��?s�E�m�C����>߀>u�>}��>rp�<]�=�0�>e�J>ȇ�=G�>�>���>4Q=E����$}��o��C�׾6�A��U�?����Dl�X�����D��`G��S�>�+
�愿5���5����Jo>������>`1׽�OA�M"?>��>Na����K>�@þm
�=ϻ�=�O%>�
>����0��ݾRb��V�>CgO�Js@>��>V>?|�q?��2?׏�����>�Yz=5�=��"�\ވ>l��>�ʠ=a/2?�M?��?��?m��=>,ʽ�	����.������Q�jEμ?=���T�]�(����Pƽ���W��;\��=J�0>f�=�!�=��T=���>biy?�A?S]%?W0۽�y�/���BG��G����>iE?�C?���>+}�>���>Z^�>-,�=��z����Z�h>���=�v/��@"���>4��>�<>&��>M?�4E��៾d5=��O==�m>u@�>�f?�t�>|�>���>�8�L��.X!��V=�yO/�c8｡C�=�e1��N[��)�gtJ�@g���;��?�2/?�$�>(�>��>O��>k)�>)�Y>��<+��=���=�=�U�:%�����!��Z"����d�=�-���3���~��鳼uD9>�E\�w?�1?.�E>�9>'jP�����ھ�7>E��>�`?�O?�l>�v��z6��t��^>���>ƒb?�*?d�%�D��<�7�8А�Ru�>�S�>�j�>�l>H�	>�q��m�;G��> � ?2�>���'��_�Y����e|�>�>۷��L�?؄f?b65���<-��{�g�?�a�w>��=ك�=d��ʠJ�r���־1F�i�)�- ����>�-�?���3�>Ӿ�˺�jJ����S�.�����>�(?T� >�N�=�(������tľB����v�>�= �^><�>�@
?�(7?��k?>�)?^Y?Z���G@?�>B(�>l�=Q?V�?�|�>��R=3�>\#����>�CȽDʄ��Jӻ�o=�aC>�kA>�u>�\Z�>3ټ�	=�Qν�١=d�7Tz�ގF=�!>�f=�l)= l�=z��>��?��Km���(�C�(���� r>�:>�Wʽ�[���Ic=�SH>���>k�"?�l�>I��)l��1޾-���^�A?>b5?P��>���=�?>�u�S獾�G�=-ي>��׺�D^�����Ⱦ�,̽ʮ�>�s>)��=���>�?^>?�@?$S �&,��T�)���݊=K�@>�r�>}�> �'>񋽾�0���x�SLN�t��"{\<N;��F_��Q<��|=Y,�>ٝ]={��=
ַ<d���"6�\��𽑳�>���>m�?��t>�"�=����ͭ���I?�v��F �˪��3�ϾX�P>�u<>k-��H?��#�}�p饿��<�^'�>t��?���?d?��B����s�\>đU>�>�y$<
h>�3l�����4>7�=�y�\������;�\>ڏz>XYǽ� ʾ����PH�ط�B�����(�����f�/���z��jE�<�݉�S5q����8 ܾ�z����`Nd�>�T��������W�{��q�?n��?�a���E�ַ'�0����N4?2���ʾ���a�<�􍾈����F�4u���`�@�H� ��7��>���Ds��Ë����"�D����#>�??_�i����$�?��>	��=�������s�Y���s�8��	?� ?dx�7q5�Vj˽�4�>���>9�>�\>��=��	y��?+K?�.	?����63��6�h���=ۮ?^�?%:?�.;�vRC�|e�� н�l�>F?�:�>5���ѳ̾�E��f
?�q3?߬>BY�w@���%�N��>��F?/'?��7@>c��>%�>?9齽򜾩����U���ֻDkT>�/�:�-��|U���
�Ue�=[{�>P�<>�[�aͯ���j>����K�%a\�}�������m��'?��þC���K(=�ݓ>��������s��_��}�I?η�?z�#?��G?�龺���"pؽ��N=���>��>� g=-����q>M�>�7߾�%e�/��A?��?� �?�2?����i���p��
��״��>�Ac��>�j��y>��=����!=7�>I�w>.�[>T�A>d�n>�q>��;>u!���W��������C�G��(>�����@�:��ӪҾ��9��k����q�O��ٽ�'��o�3#���[.���*�G�>�>�>EQ?�v0��>��H���E�C8D�1�2�IU&��\�gd���|����}Q6������e���	���~��>Rx�=Q_~>���>���=Z"��s>J0!;���=+�>�f�=t>�>z_��sD�>�N�>��=ef�=�3|>>�����������=�-����� ��?6e����>��Z�%n�'|�%3��PO?�^�>`2�=���a����?󱖽�o����=����<��>�!?����8��^-=�X{=Cd����_<G3�>J(�>f9'��_4�!���^�>��(?]������K?���>sSq?zE�>�����?�?���>8�����=��>f>B�?�^5?ѳ??���>(0�=���`o�s�;)ڇ=�J�=�<�9���N =vY��#��[�=�m�;��ռ!�=|�=�����߼m8�f��>�$W?FZ?�c�>�(�@C�؇U�~�,�.Z=X��=�6�>���>Œ,??�c�>�#1>�<�Ϝ���Ͼ��>��L>�:H�*�]�����(��<�>S>��Q?�@5?��q�he:��$�<m�f�&ֆ>OB�>3�?tt�>懍>T��;����lӿ�$���!�"ソ�U�ԃ�;i�<��M��U�7e�-�g����Q�<��\>��>��p>}E>��>=3>�R�>_GG>M��=��=ݽ�;�t;`F�)�M=���ߒG<{�P��S�� Ƽ����1���!�I���>�.�
^ټ�?�r"?g=�=��=lC��	'
��Fa�j��>�|�>�8?���>��h>Ǿ�A��	I� l�|�?#�c?��?
:�L	�='Fy��ҽ�6.>�8�>��,>ڹ���@�P�;�l=>��=A�>o�>�J��]��([�7D���3�>�����C>���?��!? N0�^2-��|+�Ds��hA���>�I��/��������;:i���u-�;̾F.�D��>�լ?���s>���L���%e������}�g�>>c?B�ټz�G=�N���l���'������ѽ�04=�[0>g�u>�??K�2?{Wv?vD?���>�Xp�Q��>�J�=�Y�>���>�E/?K�?ԡ�>\N�>�j�>�7>7FM>�)�:F����=J�Ľ��л�6�;�H>��=�>(<�2K���>fC4��ؽ	��<�����=a�>�.>�v
?�?"?���!$ͼ�7��N�����<���=��O>؁����f���=b�i>��>�,?���>��=c	پO|⾸����h�=(�?�~(?B��>����=ñ���s����=7=[>]1��	���^�4ȵ����QU�>�0�>���=(�_>�~?{�B?G ?���/���s��j*�'���*��M`�>�o�>���=�oݾ��4�xUt�rv_��0��s1��*J�2�%=
��=z>�IM>�j�=	�>ZD=�Ү�uнLt�<=2�u��>�/�>�?�]>-ћ=����a���I?e���h;�\����Ͼ=���>Z�<>:����?�
�?�}�f񥿎�<�2��>�y�?I��?�Xd??mC��8��}\>)�U>�>�=<5�=��P��!��^�1>�d�=2z�,T����;�h]>L�x>J�ǽ׀ʾQ侾\J��鿿�8�����(��Z꘾ι�2��m� =Y�A�T*^�rP���=ϟ�D=N���ɽ2�v�:!G�Ŷg��l���FP?F�\?��s=�j��b�O�kG�l�T��=�u�������d��{c\�4�p�_���ʾ��"�W��\�F�=��>䄗����MT���eD�2-o<-��>�4?�}Ⱦ^�߾�������P�=!�<��p�G���#å�B����:?F(?bb��+V�@m�vd�<)��>L��>ey��f4�;�ۼn�>pD,?�/?��O��̠�����ҽ���?��?:�4?������)����&4;���>�r<?v�>��m�a)о~���i
?[�?5f�=^������*L�g��>8X?Dߝ�f�>�@?/@�>v�n�.���*����=�΀�>:�Ͻ$�?<uw���hվI=r=9>�S�>�]������~.�>�!����q�%W��{����4��}˽�A?['��O>ѽf�n>�s�>d0�GO��������X�W@?���?��?��J?�xپ���}2>zK��R�>U��>����a��Z>ǐ?��
����C�f��>���?Z�?�7'?ӿ��
MԿ�����pľ�M徻{>F?�:B~>���M��=�>El�#�}��⺍�>�A�>���>���>NO�= ��>�����%����yIP���!�w� ��a�\Y
��Ǚ��0�~GԾ�ξ$%�\�=T��=%:�����*�DY�@D�=���>Y_�>��?eW�>��V> �"�*�P�8�iDy<V��<ɾ�徸[7�T�7���߲�������ok���!�uL0?��==<=��?s�E�m�C����>߀>u�>}��>rp�<]�=�0�>e�J>ȇ�=G�>�>���>4Q=E����$}��o��C�׾6�A��U�?����Dl�X�����D��`G��S�>�+
�愿5���5����Jo>������>`1׽�OA�M"?>��>Na����K>�@þm
�=ϻ�=�O%>�
>����0��ݾRb��V�>CgO�Js@>��>V>?|�q?��2?׏�����>�Yz=5�=��"�\ވ>l��>�ʠ=a/2?�M?��?��?m��=>,ʽ�	����.������Q�jEμ?=���T�]�(����Pƽ���W��;\��=J�0>f�=�!�=��T=���>biy?�A?S]%?W0۽�y�/���BG��G����>iE?�C?���>+}�>���>Z^�>-,�=��z����Z�h>���=�v/��@"���>4��>�<>&��>M?�4E��៾d5=��O==�m>u@�>�f?�t�>|�>���>�8�L��.X!��V=�yO/�c8｡C�=�e1��N[��)�gtJ�@g���;��?�2/?�$�>(�>��>O��>k)�>)�Y>��<+��=���=�=�U�:%�����!��Z"����d�=�-���3���~��鳼uD9>�E\�w?�1?.�E>�9>'jP�����ھ�7>E��>�`?�O?�l>�v��z6��t��^>���>ƒb?�*?d�%�D��<�7�8А�Ru�>�S�>�j�>�l>H�	>�q��m�;G��> � ?2�>���'��_�Y����e|�>�>۷��L�?؄f?b65���<-��{�g�?�a�w>��=ك�=d��ʠJ�r���־1F�i�)�- ����>�-�?���3�>Ӿ�˺�jJ����S�.�����>�(?T� >�N�=�(������tľB����v�>�= �^><�>�@
?�(7?��k?>�)?^Y?Z���G@?�>B(�>l�=Q?V�?�|�>��R=3�>\#����>�CȽDʄ��Jӻ�o=�aC>�kA>�u>�\Z�>3ټ�	=�Qν�١=d�7Tz�ގF=�!>�f=�l)= l�=z��>��?��Km���(�C�(���� r>�:>�Wʽ�[���Ic=�SH>���>k�"?�l�>I��)l��1޾-���^�A?>b5?P��>���=�?>�u�S獾�G�=-ي>��׺�D^�����Ⱦ�,̽ʮ�>�s>)��=���>�?^>?�@?$S �&,��T�)���݊=K�@>�r�>}�> �'>񋽾�0���x�SLN�t��"{\<N;��F_��Q<��|=Y,�>ٝ]={��=
ַ<d���"6�\��𽑳�>���>m�?��t>�"�=����ͭ���I?�v��F �˪��3�ϾX�P>�u<>k-��H?��#�}�p饿��<�^'�>t��?���?d?��B����s�\>đU>�>�y$<
h>�3l�����4>7�=�y�\������;�\>ڏz>XYǽ� ʾ����PH�ط�B�����(�����f�/���z��jE�<�݉�S5q����8 ܾ�z����`Nd�>�T��������W�{��q�?n��?�a���E�ַ'�0����N4?2���ʾ���a�<�􍾈����F�4u���`�@�H� ��7��>���Ds��Ë����"�D����#>�??_�i����$�?��>	��=�������s�Y���s�8��	?� ?dx�7q5�Vj˽�4�>���>9�>�\>��=��	y��?+K?�.	?����63��6�h���=ۮ?^�?%:?�.;�vRC�|e�� н�l�>F?�:�>5���ѳ̾�E��f
?�q3?߬>BY�w@���%�N��>��F?/'?��7@>c��>%�>?9齽򜾩����U���ֻDkT>�/�:�-��|U���
�Ue�=[{�>P�<>�[�aͯ��'�>�&龳�Q�	�O���
�? =��'�<�=?�c߾�[�=4\:>Ŕ@>.�$��d��CG{�vR��3?$_�?�G?��6?ʾ�d���~<�A*>�E�>:�>S�*=x<�(��>]��>	k�c�k������>��?M�?�;,?�jt��ѿx͕�ֱ������	>�"�=�� >���nK> }��A+��%�����=s�>�9k>앻>��>�,�>�dQ>D�������l���%���D�c�%�7��A��Ҡ��Ķ�l�%�/狾{s���ནځ=��ǽ�ׁ�]�8��S�m�����=��t>
�0>!?q��>Ur�>�`��7�`��Jw�<(�o�w)$���(/��]Ѿ��h�G��ՙ�<w�ٽoE
��?����.*>�8�>�q���>�d=-u�<��9>�#;>O�N>㵡>���>c�>1D�>>A>��ٯ�>�|1�[���Uw��H>�����l����Z8?f{~<��ߺ��Ծ?\�>��=�#�>XIl>$4�.x�\����?�>2ǽ	)_��E��*�b��X�>�?�ȥ���̽���Q�#�;ˡ�X�<'��>9s�a��<\��}M�f3(>J�>ӆ�S�>���>�I=?&[g?X�?q����?^��>�l2<��!>p>��>�=.�?\p\?�WH?�8 ?��>d��gC��l=>=�j��=�ڱ<E����Ձ��
��X���R5;X�Z��l�=7>22�<)��bij=�]�=��>cc?�A7?�?��7�f��C���x��K��r�>y�:?��?v�%?��>�T�>t�>�C>�>��4F�j�X>��!>��C�23C>��=��0>�OU?:�6?-"K�܍ݽo�ͽ�R>T�>���=d��>�h?Rׂ><��>���T����Y.��W��b%���ٽ��7�m�>XHH>v���_��.����5��1�=�g?|p>�#�=��_>�-O>� ?�>贈=���%����ǽ��^�O>�;�\o=3hO���=���=��ѽ���a��x��A�=8�d�U�?X�?�HQ=�&=����"������}��>4I�>�-?���>C~z>)U��3U���G��ڇ��?�9?о?V ���=���B!���>E��>�:>xG�=H����p����<E*T>���><#�>��v���:�$�Y�����֗>xɎ=(�ݽފ?��T?�/�4�������"n�i�7����=%���*�+���=�������-��c|�0$��x�Ž�ӹ>���?@�ݽϲ�>�;���B��UE��%���?�f�e>SB?��K>�j�Z&�T6���g��#���g��l�����=�v�>��&?��3?�l?��(? ?�r���	?�*=rj�>#��>=�%?�?T?0E�>M6�>�t�>���=�3=-�佣Ƃ��?��y>qO�=kW$>�M�>ք+�Zh>;|>�jJ�B��=IƽgD�����='Ȃ�o׼=��=_�v=�?#&?%]���bN����� Z�B)�;Q�=D"A>�����Q�]ϊ<�,r>�'?�r-?@��>�Π=;
پ3��u��ME�=��?^&0?�W�>ć��n��=Hk��Ti�rG�=1�?>�@'��J��	��@���=�8W�>�/�>WH�=�dd>_�~?�DB?B.#?����,�|�v�ʷ.�`Of�L��;�-�>f��>1�=K�־��0��l���`�d4�Q隽8�G�RCd=�5�=�u>٣L>/�x=RS�=��f=�=��#�ʽ{U=R慼n4�>��>�c?�No>���=�5������I?Ϊ��<��)��f<оO���>s=>����i?��e|}��4R=��n�>\�?I��?�Fd?�gD������[>�T>G�>�2.<�=��`��L���4>?��=�jy������s;�*]>��x>��ǽ]˾]��K�O� �����V��}�������?㦾�"����=��D�)�z���޾l�@S��Q�6�5�
=#P0��8o�|�.�8S��
�?�fo?QQ��G��A\1��^���� =�\U��R�?\��	�۽��a�b㬾TP���׾n�.������%��>5,þ�Đ��m�|�X�I�����>��"?����?Ǿ�Q�\y�����=���<��3
�P������?N?�8?�E���⩽8f��a��^�>P1�>#U�`,��#e=�üGX=?Q,?!���񢇿o�����=��?���?q�J?�Ԛ���/�p
��^ǾiF�>��)?z�~>Tn��\���٫�4R?�`?-�f=�W!��l���:3�o��>�ve?������>X��>���>�b�=����ڴG�ٷ��{0���>�Z=��(��N��~o�����=�H^>�N�>�w�����~.�>�!����q�%W��{����4��}˽�A?['��O>ѽf�n>�s�>d0�GO��������X�W@?���?��?��J?�xپ���}2>zK��R�>U��>����a��Z>ǐ?��
����C�f��>���?Z�?�7'?ӿ��
MԿ�����pľ�M徻{>F?�:B~>���M��=�>El�#�}��⺍�>�A�>���>���>NO�= ��>�����%����yIP���!�w� ��a�\Y
��Ǚ��0�~GԾ�ξ$%�\�=T��=%:�����*�DY�@D�=���>Y_�>��?eW�>��V> �"�*�P�8�iDy<V��<ɾ�徸[7�T�7���߲�������ok���!�uL0?��==<=��?s�E�m�C����>߀>u�>}��>rp�<]�=�0�>e�J>ȇ�=G�>�>���>4Q=E����$}��o��C�׾6�A��U�?����Dl�X�����D��`G��S�>�+
�愿5���5����Jo>������>`1׽�OA�M"?>��>Na����K>�@þm
�=ϻ�=�O%>�
>����0��ݾRb��V�>CgO�Js@>��>V>?|�q?��2?׏�����>�Yz=5�=��"�\ވ>l��>�ʠ=a/2?�M?��?��?m��=>,ʽ�	����.������Q�jEμ?=���T�]�(����Pƽ���W��;\��=J�0>f�=�!�=��T=���>biy?�A?S]%?W0۽�y�/���BG��G����>iE?�C?���>+}�>���>Z^�>-,�=��z����Z�h>���=�v/��@"���>4��>�<>&��>M?�4E��៾d5=��O==�m>u@�>�f?�t�>|�>���>�8�L��.X!��V=�yO/�c8｡C�=�e1��N[��)�gtJ�@g���;��?�2/?�$�>(�>��>O��>k)�>)�Y>��<+��=���=�=�U�:%�����!��Z"����d�=�-���3���~��鳼uD9>�E\�w?�1?.�E>�9>'jP�����ھ�7>E��>�`?�O?�l>�v��z6��t��^>���>ƒb?�*?d�%�D��<�7�8А�Ru�>�S�>�j�>�l>H�	>�q��m�;G��> � ?2�>���'��_�Y����e|�>�>۷��L�?؄f?b65���<-��{�g�?�a�w>��=ك�=d��ʠJ�r���־1F�i�)�- ����>�-�?���3�>Ӿ�˺�jJ����S�.�����>�(?T� >�N�=�(������tľB����v�>�= �^><�>�@
?�(7?��k?>�)?^Y?Z���G@?�>B(�>l�=Q?V�?�|�>��R=3�>\#����>�CȽDʄ��Jӻ�o=�aC>�kA>�u>�\Z�>3ټ�	=�Qν�١=d�7Tz�ގF=�!>�f=�l)= l�=z��>��?��Km���(�C�(���� r>�:>�Wʽ�[���Ic=�SH>���>k�"?�l�>I��)l��1޾-���^�A?>b5?P��>���=�?>�u�S獾�G�=-ي>��׺�D^�����Ⱦ�,̽ʮ�>�s>)��=���>�?^>?�@?$S �&,��T�)���݊=K�@>�r�>}�> �'>񋽾�0���x�SLN�t��"{\<N;��F_��Q<��|=Y,�>ٝ]={��=
ַ<d���"6�\��𽑳�>���>m�?��t>�"�=����ͭ���I?�v��F �˪��3�ϾX�P>�u<>k-��H?��#�}�p饿��<�^'�>t��?���?d?��B����s�\>đU>�>�y$<
h>�3l�����4>7�=�y�\������;�\>ڏz>XYǽ� ʾ����PH�ط�B�����(�����f�/���z��jE�<�݉�S5q����8 ܾ�z����`Nd�>�T��������W�{��q�?n��?�a���E�ַ'�0����N4?2���ʾ���a�<�􍾈����F�4u���`�@�H� ��7��>���Ds��Ë����"�D����#>�??_�i����$�?��>	��=�������s�Y���s�8��	?� ?dx�7q5�Vj˽�4�>���>9�>�\>��=��	y��?+K?�.	?����63��6�h���=ۮ?^�?%:?�.;�vRC�|e�� н�l�>F?�:�>5���ѳ̾�E��f
?�q3?߬>BY�w@���%�N��>��F?/'?��7@>c��>%�>?9齽򜾩����U���ֻDkT>�/�:�-��|U���
�Ue�=[{�>P�<>�[�aͯ�Z�>���V�L��H��/�fp+���<	�>�����>bR>x� >��(�H��L��Z$��C?<��?�;T?^20?����y}��=�=ۆ�>gɟ>�1P=��rղ>v4�>�s �J�o������,?���?0��?O�Q?<�m��A׿e��/n������q>��=j�>��	�Fx!>��5��
N�6���[G>��>i��>���>�ђ>��i>H>�_��� �<�������^!�D�a���G��59��(~�a��s1������е*<�kA�@$��&u������zȽ{k��Wm>�ޗ>��i>�Ys>���>)*>e���G?E��'6��gξ�L�:��Qn���>�����H[�NDX�0�ܼ�H�m$�w�/?B��e��=�?ǣ�w9�>@7Q>%ͽv��<q�>�ܮ>>�>�:�>�Wx>���>���>�r=�&\>%�B=_����~�;K/�m�8$<��??�ZH�����Ƙ;�S@ξ����Ut>`�?*iN>�'(�(����y����>�żL�S��h ��oN�	�z>�f�>fF�=�/��~6?�]a��yҽ��=�>q�>���2���˹�F�=k�>C	 ����>dP�=F�>�!�?��?i��=]f�>���>�.�>8!�=q�>��>�ߧ>d?"=&?�2?W��>شf=�=z�Ɉüą�>׽�w�=r�=��2��V<!�C��G>���=N�=���']�=U&!>�D�����=J���L ?��0?9��>m0�>�'�����C������d>Z�>�?�u>
?H�)?�O�>�=�>�)�=J�˾�R�a��>G��=��J���j���_��<>��>�_?�So?��=#��<����C����=��>z�.?�B/?S#�>��@����y�ɿ^oJ��p*���6>���!˻+��,��=����6ҏ�n����>���>CS�>�e�>��!>��	>�e,>��>��\>9�>���y%=ۊ{����;%Yd>&��=��Z���Y��A>d����6����ؼ$��At3��1����p�?�'?F��=R:;%ݘ�P.˾�{����>62.?.�!?Y
?�m�������c�<�������?#?��c?T�>P����<Ɯ��3=�<c1�>>��>k>��#�遾����7��g�>�!?�w`>8��L�����[�C&?,��=دν݂�?P�\?�-$�GB3�n=�\d���b��=<�=�ӽ�-b�����/��9پT��6� �G�=r��>co�?�'J��|>�p˾%��������C>�����=��?���=�E������������;� H;�K1=��>���>�=?��w?)��?�Xh?��0?��g���>���>�� ?�<��V��>��?2�?V�>��?�U�=ho?��֑���ѽ���j�)<�'�>!qb>��l>U��<�c=in�<��=�7d=���=��u>���.D�=:>�Q�=��=g�?�X+?.�P= �6��8H�y[-�������=�L�=dރ�F�5"�)�>�-�>��@?ф�>&0�=���;����L���k�>r�4?��?�ߋ>0ˢ>�.־8�þ�|�=�4(>��I��~������r����"I�>�<�>ъ�=�Պ>�?vJ?sl	?���g�uנ���I�����Y��=��>ٽ�>3�=�n��-޾���]B���P���/�,�W�<=���<h.�����>��=�9����=X;� ��W��� � ƨ>;3�>�.?7נ>>��=~9����FI?�`������֏��C�˻q�DT>�@�>�=;B?�w;��~������28�!u�>(��?E!�?�{g?�t��\ݽ�O>
�e>L�>�`��y(�[�N��A�5Vf>!��=�V���u�������z�=�3S>C����'��žH�v=�t��KOX�`þT�ɾ����G�_7������	M�O�����,�CQ����Pk���7��۽/Y������j�پ�׍?o9v?���<eL��5"��4��ž؊>>v׾�bi����t%�9������G߾c�%��Q�w���	���>�70��U�������[��?l���l>T�{?���n.�Q��E.�>�������$&��|��u짿ni�=�f?
�M?7D��������B!	�ћ?N?|�.>�7��y�r����>��B?7�,?��<࿧�����V"�\��?��?��F?A���^FY��(�ޏ��b9>'4?�T?qþ�:��ξbI?��?؃��S1��\
��X8_���(?g"�?0�e��~>w�)?���>�ҽ�����wd[�����	+=�?��3�s��;㡾4->��>r�M>[h���ᾆ��>Â���M�)H�_ �U�����<�� ?y���$�
>c>J�>ĭ(����Vb��t
��J?A�?�T?.�6?�C���*��d����= ��>d_�>��=�1����>�S�>0�gp����#?�^�?ґ�?�W?�fm�gcؿף��5׾�Ϲ��/>i�=�A(>�����<zܮ�N�>��=�/>B��>m�>�ݘ>��A>(��>��V>|T��~��������� �V�Ch#���F�;���6�x�fu� �-�s����L=�E���*���=���Խ���=����m���?<6[><1a=P�^>��->oG��j��v0��羗, ���|����x�/���$aa����@�=Ql����͠�>�h�;1F>Lq.?^����>�?��s���^>#l4>���>� 
?��>L�>�M�>�7�>W�,=��=ؼ=�{�e����Y,��6پ�p��a?���Q���u��/��C��U\>P3�>��=�	J����k����?��K=����[��FV��f�>��>PA/=�m4�ǒ ��T��ĉ��4;G�3>J��=g]	���n1���u�=�J?�L���I�T?wL?ilo?�aM?�e�7��>��?S<�>�A�DU�>Hup<
��>"?օ^?P&>?��>`��=	1�/r<̐�����뉽�H�T��=�tH>ǌ������[��G3=	)�����=�I����!�Uu>jT�>R�Y?x�?�T�>s���%�I���e��$��}z>�=w�>_�]>�?_�?��>i�g>������&�{�2��>��>�e���_�ߤ4>a>F%�>��U?T0?s/���Bܾc>�>��,>�!)?$�C?��x>JW=�������-{Կ��1��;��H��8ٽq�<=������`9���N��+�;�߇�.]�>;�>J*s>��E>M�I>z>�]�>�x}>���=�:��^�U�9�̽|۰�^�X>��j=l11=�sa�W�E<���,	�<=Q۽�O"���}� ��J����?{m?/�'��x����f�N���֝�����>Xl�>U?�>���>�U�=�5���U��\A���F�jS�>�Mh?׽�>d?9���=߷-���>:���>Q7�>��>�`��2��(��5��<���>��?�^�>S)�<[�G\o�Y�
��J�>`��#¾���?�<I?���(H���G�3�W��x�<1�=�}L>vW˾��L��(
���F�pz����.v�ئQ>~m�>���?�ͽ�l�>�F2�]"��������ckz��h1>ec?�l�=sEp�4�C���)�̾������a���0���>���>1;�>�h/?��]?*�%?2d?�����	?�T�>��?Da#�3B!?�S;>���>c	�>xA?Q�L>	Z�B��ȴ��M|j�a��;Yu�>���>5�v>��0�)G ����=v�'>$f�=�Ӎ���k;�\=��=�N='XS>�h>��?~ /?�f>qV=[��%CP���w�V��;᫉>�XY�?��,��m�>�S?q�V?A��>��\=j ���=��оҩ�.j?��D?5a�>�Rq>�Z�>Y,Ⱦ����N�@=��>��6�_	����᾵��Z_Q���>vo�>Ȁ'>+�K>T!w?ϳS?��?�����^J�FC��D�C�/�A�.	�=�յ>��5>�{�=Z	���3L�3?n�QjI��=�i�ν�m;����=���=m�f<��<>������=]u�=�����(�����e0�y��>�P�>VM/?��s>�;�=K��v���I?Z���j��ؠ��aоO����>	�<>
��>�?o��d�}�T���D=����>Y��?x��?�;d?��C�B�2�\>0V>c�>��-<`�>�A��-��$�3>���=*qy����w�;
�\>�'y>/�ɽ��ʾ�/���G���̿O�U����3�%��q4�Ս��V⾘��>5�%�孾tO�:�>�}	�C��=�pg���c��'����������?"��?�UI>&B��m?�����Z�W��=� Ѿ{\־�e
�r��}���t쾃ʾ���4�y���d�!�=���Y>�(�Z
�����*u7�\�8��Bk>��l?�;���:�9M����>b�;���=�"�Z꠿�����I۽�a6?�<?��ž�龆}=��&���&?��?�%-=N����1>��>:�C?�/?�5
��!��q��e���P�?ٟ�?��'? ���>�?������\��>;?*��>�l��%��1�����J?�u�>m�"���L�����"I�O,?�i�?�v���=��:?#M�>8�|����!8����*9-�T;?�x��$����^
��_�!q��+ �>�}�>t9��>R��f�>ƶ����Q��N�4��h{#��6�;�h�>d<뾫��=էX>�D'>W|�V���<���G���BL?���?w�N?�4A?[j羨����q��7^���i�>�y�>��/>fn漉��>|z�>s:��������HD?���??/�?6�N?��f���芢���پ~8>Z�=��=�4��K��tB���5=˨����Y>M�>�{>l@�>"tu>�A�>ۨ�>�B���"�Y���;��@1K���:�+i>��譾k�'��Hj��B��'8������'�=����k��GN��*�	z>b~��A����T4��De>�c>�5�==�=�	w��a�?���:���.4S���/�3�辦﫾��5���ؽ���Θ��H_�n�ɔ<?*L�����=���>�J#=S@�>���>�H=z2�=�A�>�A>Ȓ�>��>M3>���>[s>�)�=���<΁�ֆ�0	���.?��ة��I�c�c?�5n����i�b
о5��ey�<ɼ�>ƹk>�+�Bb��qw?��j�>���=8B���	�ɷ��pd5>���>�7S>�r=EQ������$"�=)��=���>�i<>yq��F�վ_�~�>=d?K��nS�=_kR>Q?%�?XGD?�!	>I0�>�g�>� ?di�=� �>F��=��>6�!?,_?��n?Z�?>�-=t���4=�!�ͯ����(����@���Rݽ�j�=�!>.v>�@)=o��=�>nH�|�=z=�=FN?�Y?�	?��?��5�0�Ed���� X�>d�'>��>q��>�?C��>O`?�_4>�$��2��ޞC���>���=�;�}�Y�4��=J��>n+�>bJT?�O?r��9)֌��j6=���=+i�=�6�>�d+?�f?��z>�e�=�����ɿ�I�HX��r���3)��A�V��'a`=8�D��Ζ��>i�@>��>���=��>���>0ғ>��>Xu�>K�F>��<�����:[�=�&¼3I�<$j����竏��(�=]�>!�ѽ���W���j=0;��ǎ$���?�=?1�&�-�d��[�E�7����A�>�u�>��>Y��>�p�=�y��HV��:�^�:���>w�g?� �>��5�l�=����� ::ܼ>ڦ�>��0>��J���,�
!��0�=�h�>��?-��>;��T�Y�Q�i���_�>�2�=�NL��S�?{nN?��8��yc���M�޾V�f���5>3�=:�X��w���X_���[��������⃟�5X>���>:��?�g��b��>��N�ʿ����a�(�xH��>}}$?d�=�<��t��gz�Um �$��!¾�$�=��>�0�>'?*0M?��}?�eI?�J1?��`���>�,�>�[�>g�=�l9?�Z�>e}?"��>[��>�Q�=��e����2}�1�ǽ�&��K��=��L>�76>�-�;h,>σ4=�m���5��!���>�Q˼��ֺ$3_=N�8>PRX>٭?�??I�>��>����uh�j����қ<t�g>]Q=P)��=�>�I?Q�H?���>��=��#��Y��þ��3�AY�>��@?^#�>ƎG>��K>L;�T�|�(>�M>�˸��G.��N���Ώ��e����>,��>�7m>c�>��?E\?M�?#���Fh�Mߍ�s�T��b��>��>K�>>��#��[��苿Vs�}�n�L籾���J��=¸7=��=�:? 7<>L	>�y=���=yEG�O�e#��^>OZ�>�I?��>��R>�F���JI��H?x ���������&Ѿ&��`�>�:>s� �/�?̡���~��.����=��#�>���?���?h�c?��C��� �=^>� R>�
>%A�<�`A��$�J��a18>v�=�y������6�;�#a>�hv>��ѽ�Mʾ�k⾱�T��Q�g�:پ��'��A���i���q��ӹ>�>�;:������9��x�Ծ�뎾@��'==�Z	��Ľx���?z9O?/�X;e��=�'��R�޾<	��M6�>
	|�悾����:l���/>��1����>ɾ�ib���!��a�%��>��=����c����Oc��`M�> �?�B ��\5�fB��I�>٪Z���>�o�Q���Xص�e��=<?E�.?���5����z�#�A��>E�?mS�=잾VE�=��>b[/?z7?,�=�`�����[Լ+_�?y��?�w:?�敻o�2�"%�SΤ���2>��?� ?(�@�ǾZt��QC?V�?�x~>@�C�æ�� g��f�>8,t?�����=��(?�Ƚ>�_��ك��S��nt"����Ƣ�>�.=<�����hx�٢}��Z�>��>�S���Ĝ�B��>1����I��#E�& ��w�R��<���>=J���>�	\>sJ>K^)�Į���������lG?�1�?�aV?9�6?z{ ��=о�s��(R9=Z'�>��>T+�=����>��>��پ�eq��"�{?&��?�#�?DLU?�$l�Q;տ�����zǾw]׾d�L=�j>���>Uݼ��U>�w>���<����<}�br�>�>���>�,>�$>�}>�i��,��N������9�G�2�C�����ņ���p�B�!��������������!�r��Z�$����r̾(�ѽ/~�>��><��>���>��~>j����]���<��Ǿ!&��E���~ ��������@}�ڃy�M�>낯��+�3=?��ѽV�{>&�?�����^>��>�!���C���e><�H���f<$��>�`�>���>Y>�������=A0=I+}��ϒ�b`�0 ����н�OK?�
�"���b�����B�ؾafj>B��>��K>�hE�c��N@z��k�>�d0=�x��i�t�Ҝ��f|>a �>�}.>�j������;�Y�.�����e>5ޣ=3�'��Ǎ�ã��p�=D&?t�6�=>J��>��$?��?׋*?�Ȁ�� ?�׳>�)�>˶�=�>sT�>!;�>v".?��e?�A1?q^_>+S;>�v%��Lb�����/��:�	=���=�����<�Ȏ�;"�>=��=dI>���=�:��j���a�g��TT<J��9���>tBG?���>8��>��S�z�?�G�R�N�-��q|����S��>ı?�?�Q?qN?�/u>�Y��`�9%���>]��=B�Q�f�]��g>g<�>0]�>�'?@?]��=�"��8�=� >��?��?ބ?�[	?��#>�z����
��տ!)�A�*�rh��/�`��<�=��� <��_<�H�liX�dY�biW>�>�>4x�>R?>M)>oD>�x�>��E>��=�X�=���=-���!�ӽ�D�=�缸旽le��*U�<]/�<���0��S�@�퉽p$����O�B/?��?*<)�a�+��Q���z���?��~,�>�9�>}��>}T�>ľ�=
���3�S��C���T���>��d?JK?$\�s�=��<J�d;�X�>i�>�>�����M�nĔ�Eg0�?��>�?|;�>�Xӽ�E�ug���5u�>X�>=r�m��֜?��V?��(������fG��Ic�߰��Z=��V������پ[�o�CX-����S�R��F>| �>�#�?�鑾���>��F����y��v�k�=�AJ=�G1?#�.>�Y��k" ���5�ea���Kݾ*��f>Ԣ>��>���>!�%?��Z?R�*?�U?�[ �i�?��>���>>Q3>�n?�s(?/�?��>v�?�')>6���,��^E_�s�R;}�=��=��^>��>%�l=���r�l��>=���ʼKm������ ܼ�,��gR�=�>˻?+#?��t=�4!=ȑ�=Xq4�,�����������>%��n7�i?�>!3:?� R?��?�&">L���#��oȾ�;:D�?�F$?���>7`+>.�r<������=��8>s��=ߓ����ʾ��<���U<Y��>���>rŞ>	k>ϊ?J�M?A1?�S��t�a������2��G�U��) �>� �>��I>v͛�+A��6�6��_��G��41��U��L�=�a(;�K�~��>��X=�3�=�a>�f����A�@A˼X<!�>�y?X�M?���>���=pھ�9�;�I?�џ�P��`���о�N�2�>5j=>*����?T�
�d�}�!᥿�<��?�> Y�?5��?]fd?X�C�ę���\> �U>��>k)<se=�0���s}�T7>/D�=�v���x��:��]>�Lx>��̽��ʾZ����<�&1̿�:o���l�_�0~���Os۾�>��:Yj��%�G��⩾�����{�dPP��.,���ξA%�%���{�?��?�	_>� ��3ྸ'��@2�.��=kҀ�����򾵠X<@"�8x����V��n�xO��K	�s,>,$!��U���؟��ݾۮB��f�=��~?]Vپ�G��"��$T>:�8��ʏ����M��}§��ƒ��C?�H?�ԾO�����=��8t ?���>U >�D���6�<z?�5?!.?s-����쟱�T�=�%�?���?/�(?'"��m�o���ھ����0>L�/??�	���$Qm>P�?Y�>M�ǻ��x��դ�#=�ki<??�?�*s�!�#>t�-?�8?NL���ʛ��c�=ܑ��P>>�x7?O:�<5NԽ� ��7�a�K>�?�1�>V����r��>�]־t�>�<�z^�&���wQ=�}�>wi��>��=���>�>�n �ԯ��!�4�;�fz=?�ܪ?�!V?`�&?{��V�\��,8>=��>��u>���=]�)��y�>z�>�=���~��p��`|?�&�?j��?ަK?Gp�~�տ�|���@�����D=.Ŗ=XZ-=@�[�(�K>w;�=m0���	���+�<�M�>[a�>��q>?�G>c�	>}/l>m����P�1��t1��o�2��r�i5:�7�����ݹ�n��Po��Q���#�<�ڵ�`��4���
���Ǥ�]�B���<^��>���>g�y>��o>V>�~N�� ;�n��[���E���+�:O����߾K��q�G�gVZ��S�/�5�S�=��v?).>t>7b�>����=xx=!�>ؓ�=O?���==k>�;�>q��>;b>OQ_>�2�<�\�>��>�1R�i6j���:����Vs?4��=�.�
���o^�߁۾&��=C�>;T>I�1�������� ?#�P>~3��v�ҾC��M#�=i��>�%�=\�$�V{��֚��K<�� d�=Ꚇ>�J�=�3��칾���<�_=p�>a��+<I����>^݅?��?ap?�S��z��=�!�>*��>��(���+? �>T�>*F4?�^?�=M?��>LΆ:b�=�0�=��=��C(;0n��E㟽�ᄽϾ����<PM#>Δw>��k>.�B>�>ƞv=��[��C��3	?��N?��?�
?sey�2WD�+�U����6���w�����'?.��>��s>C��>`Aw>\��=�x�������+��x�>��>��M��R���@���j!�QG>4�{?���?$�����%��b�k&`>���>�?�$�>��=����Q���C���q;��y�Y䁾��=�Jn���2�bR�=ܝ�1����:��e^��;�>AF�>�L�>j�4>i:�<�ӊ>���>{nm>!�>�d]=׳H�P�<�=u�F�Q�!�=�{�=�&���������}���<��=��;�'�,?�.?OoѼ�L6=�V����;�1��f�>>?���>º�>E�������'���S#�Զ_�4�?�?�?��=�:�ǻ��C��@�����>�n�>��>;��*.��JV�����l�>��?�_�=zU�S&��W�<����>+W9>�ॾ2��?
��?��?� ���l����z�
��T?��o>�`>�uA�?i�'�:�����R����<�h>���>��?$���#�{>��N���&�������!>Y�=��>�\">�{�떅���(��KԾ!���_낽r]�=�%X>�P>:�>��?��o?4�=?�W?&�@���>�6�=,y�>��'>�=?mԶ>0M�>\?�:�>� `=��D<��ҽ�T�ڱ(<��=\�o>(T�=��>�0�<H�����t<��P�j߱�����3��6����S�=0�]��I�=�>��?\d%?��=�}>������Tt�;fM=�<�=֥#�������=��?V1?V�>��O=(w�t�?�E:龺>̽(�?L?��>mʓ>0��>
: �B\ʾ��=�<>�C6�򡊾{V��p���#���y}>��{>��>���>�҂?��K?43?������K��<��/$�������Y�>tU�>Θ�>эݾŢ>���{�T�d�ޡ5�3H7������`��u;">��*>(�>�Y�>`�;���=��E�I��>�>ߕ���=���>5�?�A�>)��>����"��J�I?3����J��R���Ѿ��>��;>:��?�� ���|�O�����<��Z�>;��?`��?Y�d?��C�K@�z1^>��Q>zr>ɇG<+�E�����N���C>�~�=6%��o|��p�L;"�M>1�q>
Ƚ#�Ǿw�޾��?������؀��Jξe.�������jc��A��?���Ʋ�`����x��|��h�=WR�;P4^�s^����ݾw/�?�l?m"�=rg����!���Z0��X��>X�=D���ݐ��[��mh��闾���:�!7"��,�Fh+�Y	�>��s>����H����@D��/�h>�җ?ni�'=^���L��(�>�ܱ���<ux�̪�(��#xo=gP?N�(?�Tʾ��������<�u	?#�>�|�=����v1�����>���>MX?�|Q����i��j���i�?�(�?�DP?��=o76�i��I����f>=� ?!��>�EL��y�C@ھuKP?9pC?�~q>k��Q��{1V�v��>:I�?|�"õ=�W?O??�Ⱦ�Ԇ�q;�=��'����=�	?�2��~��B>ข�/��=�}�>>�>.ž��@��??��V�v���<�;��->��>p�?��d�:����>���>�!�N�f��������DlO?��?c.|?!��>=�V�M��ǰ�W�d�z�`�� ?�)Y=TŬ�z��>3��>S��)������ڶ>�Q�?s��?�?S����п֞����Ѿ�$���>>�ޡ<��H>����`�2=Jb�'*Ͻ9�2����=R��><ZS>a�Z>3pV>
�8>��>�n��7(�҉�������\4�M���k�Xl��3
�4ؘ�̲�EH��Yq���%Ż�+���i��GZ$������z!`��%>�9�>��>�?��>�p�>%eO>r*�����_=�>�v����`�����鯾�O��=��Ͻ�J�|Y��5>?�i�<)��<K��>N �c�>�;@>�ȁ>_+깤�>tl^>[�>(t�>�1�>�d�=��{>�M�=-��>ܐ�=X6��Ӝ��Z%4��P�Ť���&T?���J5R�ۀN���ƾS���P>}?��@>h�&�񈚿���Ǌ?Bᆼ����B��@
�k��>���>tv9>>:.�פ,��3����y��=G��>f>�=�*p�A���k#�X�=�3�>5����R�=�;>r�1?��y?�<?;B�>�[a>���>�l=`|=L2�>Pѵ>e*?U�E?��?"��>m�C=��s�4��=6JF>]���j{ѽ����
�����s�D艽w��=ǐ~>��=줫=�C�����{ҿ<���<�z�>y�A?�h�>;Q�>������:��KG�]|y�:'�<0D�=G��>���>��?�i�>e�?W-P>��'���/���.���>?��>�	{�8����`߽��>�`>��?�Ye?W��<��Ӿ�8=_��e�?W��>�H{?��>Y��=V ������NĿ��!�x�̾ �<d�ҽ��<B;����&���M��Xھ�����5=x�>I��>��>/1C>,>I�*>GB�><*>X��=�v���9h�[�=�g��%�<6�$=�"->n�ս��<�C<�M:�ߵn��M�����w㝽�˽��X?�?EW�6<��C���s�/TX�q�>e�	>�7�> ;�>~���#��%o�!j[�w����>�>[AX?J�>=dɾ�wG>�K^���(�T�;?�m�>���;ߓ���ӽ�Q����P�B�F>�K?X��=m����R�����A��Gi>D�>������?�]6?=)�s'����.�58�Y�>�(�>�|.�!��T��;M�=������K�F�o�\RY>���>N�?�>P� �����i��ue����蓗>T7�:;�?0@�=��F���G�Hy����,W��#I�>]_�=Ț.>�D?E�?݉�?��?�8[?����6?���v�>&�=��>-Z@?!�[?Ƃ?��?F�.>�~ �-��-�ш�=�5>1e=�p�<0v�=y�L>���=���<�:":�F�������2<�s	=m�۽��;`��;>83=ޯ?�BG?h`x�^�ھgC���b>�'�=�>�=���> �n>O��҅�|�(��e?t4?v�=?�5n>eV��&�	��Ͼ�"�<L��>�L?,��>D��=+}l>N*�M���=y R>��2��Ś�9ا��n�O0[���Y>�)�>��1>���>d��?��i?�1�>!�l��O���f��t�D��+>�K�=UY?z�+?9v ?�{�7�-�dZ�Lss�J�3��X���+�Ѝ�~��=��>5PF>�ш�.��=���4c��䨽jD=��=�0�>���>�(&?u�>�y>������ �J?Bo�.���澺��&��=��q>)J5>^l�<��8?��=^ol�%������#�>��?�:�?0P?��?�Geg�_�j>��>.�G>h�D>��|��.������<v��=�~8��`��  ~��h_=��G>s��ܮ�p���L������@�Af;����֙@�냽��Nܾ�	�<t�7��:>4�J�����7���K1��K�� �;�0m���Ӿ�l;Wӡ?o��?���=�a`�rS�� �s�7��#�>��۾����tϾ[���pL���9���þ'O�տ0��*@�?'��?P�d��D��̙u���$�瞞>ֻ2=�4}?��� ��Z>$�;��>>ɻ>���:�����M��������X?� X?�#�A)6�ʤ>���=ި6?�?�&=v��/���!a%?�(?A[#?��=����[���m��;�?ǫ�?X�N?{����Y������^K���?N�?#�>����$�9z�˫?��6?8Y�>	��P����(�� ?ڼ|?l�E��LK>W�>ӈ�>��-�h���� =����Lѿ�J�0>�9�=\eJ��͙��H�|��<��>fb�>pꖽ:��Z��>)���x�pb-��@)�I�o��g�=6�>#����F�)��>i>�!-�Wx��<�� J���;7?�u�?��v?;�?</�����f�����9G����>����B��T��>?�
?�.�q������+q>���?�%�?��7?ĉ��x�ݿ��XW�������.>"/�=q�=��>�@�=�ف���x=��߀�=�9>/�K>n��>�I>��>Ã�=Т~��G�6���5���h1��a���(��h�Q���*Җ�4��_��Sƾ�i��<��W��HIn�'���_<����ev=��d>Ť�>~.�>t͔��|>>�W>��O�B����!���8�3���?�~-��ھ��@��>�B�����Z:���,?tX�==�=�?OҐ����=Ċ�>�6>B�3����>�=x�>i3�>5:�>>�G>�FO>ל"=�v�>���=�jd��d��D�>�w8R�f�?�L�D?W�����	��!r�9�+��)����>N?�S�>�A1��ꝿ���PZ?Sk]�,~ʾ~�3�1@����>	�>���;��>!=r���ݔ���<��x>.��=a��g�:��X#��h==mW�>s�оY� >��>�},?��u?)�:?�х=3L�>_�M>Gk�>Ώ�=��R>�c>n�>�T?�|<?�C.?�I�>
�=��g���<g�L=`�2�v,a�����?�����:��<	�����|=�4d=�j�I�A=�a�<0�.��zĻL�=ĸ�>@�J?pb�>?Q�>�M
��m7���E�����f��>��2�e�>��?��?M��>�1�>���>>�b����$��>?���=T,��M������ˊ
?�|?�IQ?-^E?)�<�Kξ8�E>�$�=�CT?&�'?�v?�)�>
K>hl���%z˿�6�G��;����\Ƚg9�rF�"����ȉ��==5�<�J>�%N>B�j>��=��>�SZ>��?u�Z>��@=>�����&=��F��u��>L�^=�W(>���:t>0��X)�=���o����P��q#$<��	?)?������Z���ɾ�>��꾂�ӽ���>2RK?n�>��޾Q�5�l,;�M�`�hs���=���?k�8?k�!���+>��=��$p>��>>��<�&>��e>�v%>��罺8>���>��_?]ך>���=��V�O0m���ڦ�>ܳ�=������?|mC?n=+�d�d��$��e?��{>�ˈ�;2���ȭ�������A���A�u��P�ɾx]����=V*�>l&�?����m���x�1Ƙ�aэ�锾��<Ui��|4�>٘=3T澻Lɾ�E4��L4��Y��~"�>�Q�>��ؽ�i��d�s?�!v?�&z?-.�>G|?�vv���>8v�A(?�{~>Q�#?�;?7�W?W/?d�?�5>zA�5T��!᯾TR�~x���e=/�=�
�<�	w=�V�=ٍ�<бa<��>���O��߼pȶ��ʽ̯<_�>�'?��Y?�(��ߞ��~=4��>?9�=7uW�+:�>�X�>rgt��.ؽk��>��6?��G?_j;?�3�>�KԾ{R� ����>="%?ӏ5?�Z�>ȇɽ��=�'ľ��Qս0�>Ү[�{.����پϳ��?�#�>�;�>���=ǘr>�mw?'�?8�.?N�o���������[;=:Y���V�>ȹ�>�L{>8[�����|g���]�~�B��Ec����T>�X�<�3޼ށ?犢=�"��M��_]Z��y����т ��>�>1E?x�>\�=�V��#%�"�H?���91�#3����p���,0>�#>�Y��z ?�.5����ٔ�� �B�aW~>)X�?Jn�?EOd?����Y�@ђ>�`�>E��=H;=n����n����q�s�=�k >vt���W�� �	�T��=��=>�l��1�׾
������
��t]_���ս����K�@�w�Ⱦ~㾮�?>�C��"μ~�;�@B�=�욾Xҽ	�$��h������H��9��Cܘ?3du?�z=9�y��4����Z*��o�=abѾ��8���D�0��u����Ͼ���Μھ�'+���D��,��>�>& þ����Q��?� ����>A����?�疾_)����2�y �><�=>?���x~ ��2��ԗ�����`�m?��M?wk�46 �4�c>r�=ڳ?�G?�=�sm���??8%?+���t���ߛ��a�;A1�?��?��D?ȣ{��{N�p�k@��Z
?4?5}�>m���*kܾ����ދ?�1?!��>��a������#�?�Il?43I�Y�j>G��>z��>\��R����
<	���P���P*>!�P=A�<�q}��f�7�E�Q<��>MS�>8�-�y�1�?G�$��z��5�804�r*>U{�� �>�� �;����i>���>qmT��g��Z���堾{cG?6I�?��q?"K�>D�/�+!u�q�C���rH��P?x�W��K����=�kL?�2*��W��jd2���>H-�?�k@L?�o��1�޿Ҹ������؞��^>�V�=A9>>��J�]�Z=�*��B�L����>���>ɾl> ��>� [>٢3>�/>���u�����d}��)�4�8��Z�������"/|���������Z���n����Ƚ��l�������W>�Йþ���=��~>���>���>��>�m�>> �p����C5c�]ݾ� �� ������FD���
��(滓�>�6���?�<e�<=Î�>�7���f`�O@?0n_>HA)=�ŝ>t�q>��>~ZK>�+i>�u�<�uH>uY>�@]>�� >�Ӈ�!;��u���m�P����3�t?
(ս䉾!�F������B���r>jj�>+,�>w�"�E񞿐0h��i0?�w��/!�H�Y�=I��?��>�ׅ>�m4>�뭽8|�=c�������f��=�ܴ>�8���N�J��e7[���Ͻ�j�>[�־�$�=! �>�D(?	�u?��7?�R�=ܽ�><Uc>N8�>���= aT>�?V>ls�>�?)�9?��/?���>�ص=Tjd�V�
=�>=�:���9��ů�k��h��<�#�e�Y=��t=`nn��H=Ó9=�÷��j�;�� =�X?Q�=?V��>� �>1ӡ�ʵU�*�A�6�T�똞>���=Q�>tt?DX?.)?3��>a�=����ߺ�b��z�>A|>��� V��R�ǽ���>��1>�,K?�J3?~->bB����c~>w�O?P�??��k?��>��e<;h��2�Zο�!Ӿ��(�K<<~��[<q��>�!�&����d��:غcH�=�cU>�;�>�IB>��=���=
3�=��>�I>�l�=���;���J`,�������=�������뀽�2�oн����飽e���G�4��:�ͽ�S�>�s??����Z��"7�>��#�����lg>���=�Y�>���>׃A��\���\��da�T�RM�>�9�?Κ#?:ʯ�fq�>��B���� ?|ih>)O^>v4���b>�4�� X����>Z�4?ڊ�>�!���$U��ƃ� ����>58�=/�{���?%�L?���6�Y���9��`E��-����=3xO���������e�D��2��O��΂ҽ9T~>ک�>���?�u �E?�����U�������L<l����>�K�>����'����Y�׾�D��� �?8�>�Ș>�r����(j? ׃?�V?���>H~?˘X�k�?F/9>��?�t�=ߋ5?Ȭ?�Lo?j�>K|?�Ʋ=�D���Q��_��� ���6�B�v=��C=��<�tq=��<i:��g�=
�=<��ZlN�RĜ��,;F����e=K�=@G?��e?�FQ�9��&��=�He>}o=~�=��?{�!?�]���n�?}:_?��K?�(8?Y]P>A�ϾFH��	�����y�>��Q?��>J]��3�>bƾ��B��'A���>��)���y�mgA��nӽ��> �>�T>�r>�:q?f�?�+
?T'�N�h�f�l�6�C�{�<���{�>��>�%=Hg����O�.6��rՃ�M�,�M�>�wm�O���w�<���>��:=>C�;]��>��k=#ci����Es�>NF�=��>?`�>8�L?���=��9>����7P2��,N?%�����.����f�V���{���a>��F>�*Ѿ� ?��W>Rj����1s�d��=�&�?�?Yj?7(<�T�۾�?|?�>�&X>�B�>���<rϽc%�=�w�=$�>�Kz���ϾՊ<5!�=�<k>DW�9?���`���G��
͸��N�,g��[V��P٘����򲄾�l�=�#��$N�9��鹾����M���ps[�aʹ�@���Q�-Е?�TQ?>١��nd�j(�ل��՟��Uk>Z��[��~����^���u�6����ݾl����s��x��	��(��>����p`����x��o�}�>��(��a?~�ξ4w��}bB����>� 7>9t!�a�����b��%o[���O?ma?\d/����ZPW=J��=��?`�> ���-��s����}>ZEL?�~�>;�j�9z��[?��:s*�`��?V��?�@?��O���A��;�����?T�
?D2�>�d���̾Kd���?CO9?���>{���ܢ����>�J\?�#N�Aa>W��>nd�>am��ᓾ�"��^�����ݗ5>�%��3�Vj���?��s�=�۠>Hhy>b�\��i�����>�k��%M��*��D������5?<��#z�=��>��.>ɏb��ሿ� ��,2�ӸR?%�?QOs?��>��<���j99��>�>"���̈�>� >��ͽ���>��0?���l��JW��9�b>[B�?���?[dD?W�u�>Gӿ�� ��������=%�=��>>��޽�ɭ=��K=�ɘ�DZ=�l�>��>o>D;x>z�T>ϛ<>��.>q�����#��ʤ�4ْ��[B�� ���wg��{	��y�����ȴ���G�������7Г�z�G�^���T>�	���,��=�w�>�?lz�>Ε�=A-�>�R�;�FD�1\� ������|��n��~���\���潩w��l� �;����?��f=�}Ž:��>l1н�W�=��>L�S=��=�r>Ⱥ>+�=@/�>�cO>Ճ�;�T>�[�=g�D>�|z>¥���:���������t���-?J�<U���o������/�Mu?Y� ?�R�>��5�����^�z��I#?:�D���m�m+�L��>H��>(�>Gs�b���𺒾�����@�=���>t��=L�=�d��[�[��Y�=	�>J־(��=h��>�_%?�Lv?=�7?�a=���>�BH>G�>�ɸ=8�K>@�Q>ci�>�+?{B6?�k.?�8�>���=��X�7%=�s4=0�D�4�G�׫�9���#�J����;p�P���.=1�9=4ڛ���7=��$=C����Cg<��!=��><XH?P�>Oʧ>��2���P��mK�B��%>D/����>m��>}6?�h�>��?��i>��s�3o��T�47�>��S>f�2�B���_���)�>>?>n� ?�l?fU���;{�<)xV=�o6?��>�us?jcs>;b�<�??�� ��ռ��RҾ8�⾦��=W���0꽤\`��-��aE<�<�;4����	���i�p�F>�P>c�>�뻈����?ey4>��#��9$�Ʃ!�����Jn���=9��>D0�>��=nO>�μS={½~�=&F(>&'>�'�"9+?�3�>�2��=�m����I��b�N���ҺgW�>��_?}�!?n���{$�����rg��c��\1�>���?�}!?��Ǿ�jE>_{>_�%>�D�>Ś5�G��>�K�=8|��D���b�>$l,?��!>@�I���T�<T��{SB�XE+>w��=���JK�?��M?��L�	'[�� +�>K�9���NI;s���;�O���޾�M7��@�]���?z�n
��6>OA�>�5�?(ތ���P��b��6����W��p�����x���o=)1�>Kv�<�tܾ��þ@}�"i���R_>X��>�$*����=6y?��o?\�,?L�?>z?���S3������>�P���4�>G3?�O?�7>��>J���Ӱ���������:�w�,�4��<�?>
�ȼCv����,��JŽh��=(7= ~���د;`Aýe�:��ڽ�E+=��=��?=�`?I<>b/��������28Z�"<�q?O�>�@=B���Xk>B`�=�q5?Q�@?��?���>�Ů�FB�����xp<S?��??���>��:�A��>�ʧ��ž���=�g>3���?�3�9����m<����>v{�>B�!>UV�>p�Z?�2�>��?آ�=�zk��o�)�ھ{q��ȥѽ��?��>���>Ù ��b�jo���d�R2��{�ݬȾ)0�;8U~=׾J>�r�>g7I�B�J��Z>_	��*�������"�ܦ>�{>ŀn?��>Y��=����s ��G?��r�0���@¾Ƃ��=:�W�;+=�e�9�V0?:ݼ�D���ô���1��I>�Ѷ?���?ˍ?:���	м=`L>��P���=5<$���3��[X>b7���-�>�>x[����<�8>��>2%�>Ӗ���оH���$�e�^����]��{�q ��,�X_��I�ǾkR�d=�T�{j��w���4�e�&��D��k
��F��짔�%����ҟ?o�<?k4�=�����#���4�*���t	�j����<B�74�ooѽ�;e�&K�W�x��%���9�/�)��پQ��>�#���ͤ�A���h(����>R�#=��Q?�[b�_䐾�"V�Ҵ�>ԟ?��ʙ׾�~k��������h�x?�mJ?�,�����V�x>�j���r ?P�?�/>�����E"����>h�G?W?GAξf���������aE�?��?w�O?uݙ�Y���%�m��?��>��>r�K�ݾ����5?(�=?�nv>�)��ي��1'�n?Ml�?Ivt�q�>���>�ؖ>|�ɽ� ����<�~���)���N">YX>�>I�z�ѾTk����ȽC��>���>m
ɽk�˾+�>�x���h5��B%��W�y���n=�����>�3��.&�=�@�>k�>��E��2�����E�u�!�?~>�?�)g?=Q�>�	Y��Ҿ�9�)�>:�Z>q�d>�,	=�Q���>�d
?J,���}���羋��>9S�?��?�%9?�x�JgٿHɩ�����'oh�ȉw=�$>�Nn>j����R��V�U=� ���
��4�,=[H�>;ݸ>wt�>�r�><Á>͚R>D����!"��.��7l��*V��i�"��p.�����<�c�B#��J׾a�辦YN�|[=����ܽ����y<���E��=
3�>��?���>��B=6 ?���=ʾL��KҾh9�=��r��G������g*�r��e��������(�#5?�O�<�{���?DH���dd<xT?�Q�==)�؝l>�^�>/��>��>�a�>�y <�_�>e��=��q>bL>��u�P�����������V���c?F�1�F���T�j��յw��o<>v��>�߬>yC�r���W;{�>�?nR��Ծ�[;�	�$��G?�~�>�/�>�.����>E׈�4�l����=���>�6]=L�ֽ>�ݾL��*oɼ-
�>�m��Y�> ��>�"?�7o?>?�o�<	��>D[�>;+�>���=D�y>MA~>���>R�?R'E?!�(?�p�>{��=�!p�lc=�@�=!h�}���o���$�м�M��lX<�j/���p=���=�1�yj�=	Ss=�a�������&=�/�>�41?Sv�>G��>[_b�g�<���`���.�;�;1+��jd>sP?�0?kN�>KG�>n7�>>lI�Y1���!�Ҏ�>�I>��N��h���UH����>��>�	^?g�S?3$H>�&�QX�=<"��/"A?�(?*�p?�F�>Kd~;S��%�	�2�߿9���ӵ�e$>b��t"<�{ܽ �y<9:�_A{��w�p�Q=;�>�w�>�(�>�S�>�.'>=��>�+�>�4�>߬g������=P2�}�N�է=��6>�������y^<�ܬ��g7��-��չ��KՀ�v鯽���)?C�3?�㈼HK��8�û����KV������%?7!?�J�> �|A�.h���n��m��ݾ�>v�?�4-?�?E��;�=�<.z�=0��=m5G>m�W>¡�ɤ��������=gj�>(�?��>���V@��`�����t�>�f�=�����o�?��U?�*J��;q���	�Ϻ$������=�:��d���O&�L�9�8��`_�Z�ƽ��z>���>O�?��LY
�V�,��ň��3�����@�=��:�\>7LV=���ۚ޾��&��,��3���S>	�>�>�}�>�y?�d7?ZLZ?zm ?��U?u֘��°>��t>�й>�-�>J�H?L7&?Q4?���>JB$?��:v�}��)���1�M=�b>-�^>�5�;Pl>ZZ=4��=�7����(;��<���<E��A�>��a=,ǎ=|*�=�0#>�?��9?y��<�|f����斂>G"q>�<&>���>�Aw�ov,��ެ>_�h?|�B?(W'?R�>4K��2�5�{����<�!�>��1?oВ>��<��>{����|`==��>K�w� <�H��2��ED���>�H�>�HS>H4d>#�_?�y7?��5?������B���_����h_��ka� ��>�.�>מ�<�W,��")���w��L�W���#=PV������:>���>�>�3μ�PK=��k>��
��d���=7M�=4�>z��=��6?gug>�r�>g����]�
5I?k<��ɔ�5ĥ�z)ľ��/�=�$>%��!�?����m��Y���&A=��m�>�i�?̀�?�nj?A�1�qc �]�d>Ԋ?>X�=ý�<�N$������ҽ
�G>e �=/7i�l��Q{<�l>��t>�pڽ�ѻ�$�׾�ar�����.�;�9�p�_qþ��+���׾Z�K=e;�=j����\�����=�y��b���O=\=��ʹʾ�疾��? ��?D��=Q���٣2�������Ǿ� p>�^\�y3��oѽa�޼�[����7�̾�9۾�1+�%�$������>7�K�e���)�w����d�>t��=,�e?ɂ��Ͼ�	뾸y>��>�X�oо��]���+.�o�9?�*?��v�ྒ̙=�V����>Ч	?�ԟ�*���pj5�a�>��*?5�?�7f�U�����$$�����?��?�=H?�CU���`�":��TL��m�>�`?f��>a{��b�꾆ͺ�<�?��1?�b>�)��a���:�~� ?�5�?��|��*�>30?D��>M�1�e#��N�=U��[ �挗>l��=��*���Ǿg�Z�ѽ��>^�>�	����?@*������-��Q����<��=$9?l�0�	
�MT�>[�?g�۾Y�N��<��:���z?5�?�h?:�0?+�@�R�>�>�>��`>Bxq>�䇾�����df=��>������_��i�N��>u��?�	�?��0?βt��aҿ�Ә��CO��C�H�>Y#K>�d>%�c��,=�ͼ��f�J�f8�=e�>��D>�o7>�:�=�$�=�\�=����M%��w��|oz���P�HL����n ���m�b�I���������{׾jj��Pq��5"�e���.H���ǥ���ʾ�!=W	�>}ze>���>]��=x�>=�se�ov�����$�� �T�&��5��e�z��z����rU��~F=T��� ?.�APH���y>�Q��W�=�mC>�`>�dx=���=��x����>XII>�<�=�!�>;�v;F!>i
�=���<�\d�ۡz��/�L��9�=*%.?�޴�p>ʾ�F����	��t��>CN�>�=J�;�잿�Y�0�>�sL�G�پHX���g�=vE�>�4?R��>.�^�,���D־�oQ��=��>Z)>H���0������֕>��?�$��%���0�>T)?��|?�@J?��>��M�=�*�>x��>c>{
�>%�����=V+D?VW?��D?�>&�<��<\�>�\�=�����[-=I6�:W�;N�>j->����=u >J��<h`�=��_=��r=���M2�;{��>�Q??�>�]�>{����n�
]V��.\�?9�>M�_2?fc]>m�?�E?�*�>�}!>!"+�C4�����2�>��>>8߂�{�����㼈�1?���>��0?��><T�.w �;4>�~�>��>L�?M7?�Z�>�T�<���Zk
��ҿ�	��VМ����M�S�{F������}�kV<sž�j�!�N<Y��>3B6>0�->��=Y��0��=���>��E>%��� -�=G!�=͒S=w�m<�2�=-��<�L�*'޽~��Z��*�����d���򇗻9C�<<<�?F*5?[3���_p����Q�,�ߞ��:%?zK�>̶7?J�?��<��q]��b�c��/X�>��l?zk�>�^4��A6>*Hn��+��.�K>�K�=�ۆ>;�>�:<B69����>G+�>��> ��>��f=������po��O�>���=�b��ǒ?7�C?4R�we���S?�h%9�a��%�:�� ?�Hش�����6��Z<������=n����0��?!�>�ϲ?���FN�=�?���:���:>i�x��=��J=p>�Ჽ|������B��5��� ��V�=�P�>T7�=Y ?�=^?z�>[�%?�)�>�?����;?� V=�s�>���>�A?z�'?t|?b��>JŊ;��L��=kA�M����%>��<�!~<m	�%'x=B:�:��<�	:>ٻ�lی���=�=�愾8�z�kϺ=;��<7;d>b$?��3?AG��F���>�!�I�>h?@>���>s�.�i`R<�ڇ>I��>�?��N?.B�>���y�;����]�����%&6?��/?I?�W����;����"+:>�e��t+�{6���	۾b*�<2�:�bc>��>+��=�||>�y�?�E;?}]<?��־?����"v�����>�l�>�>�X�>��~��㜾�徣<���d�>��s��>�y��S��<�p�>9��>��>��=_��H�Ŝ��T�ؾE��=Bֽ��>�t�>	��>�:�>�;R=E0̾�E��]?�m��Y6��U�=};����
>�1>
�	�����ԅ?6_��5�z`��nv�K�6>D��?�3�?���?���pF^��x�>��">'K>鯷�������<���l��>�*>wӆ����$X�<*�9��(>�%��Ӿ�;ƾ
^���mʿ{Fc�h���\�.��.K�u��5���ɾ"|���{S��p7�m����ξ�r��	)�I�V�2#پ�`��	˾`{?(j?[�1<�����= �3�Ͼ�iy� s�=�S���;��P�������̾)6Ǿ���{��������ׅ���{>�똾4�������i+;ْ*>�)�>".I?���V���:���,�O��=��>H��(������/�{�}?�4b?Ô�L�?����o5=��>��=�7B>Cy���D>�M?d�}?�Fb?T�=/P��UK���>c��?�p�?]??�]/��=���|K>��:�>8�?��>NX~�Wᵾ��ʽ<?��5?v	�>%<�/䆿T���3�>��`?�#L�GXJ>�<�>K�>�맽DÕ���*�X���N/X<w='>��ټ� ��Uo���K���>���>SJz>��w�TZ��xV?K���鑿����;Ծ�2>������?�5�&�<>;S�>�>��Ͼ0�x��􆿸����X?1��?@��?�S*?��ԾJæ�B]>Y�ս~�
?\Ь>Z+��(�޾��n=iw�>���}����IM���&?���?T� @o�P?U����$޿�Q��g��z��L��=�Z >���>���X�=3<8�h���<��I>g��>[��>�j�>�>�>D$�>���C:(��-��ǀ���)@�T �'�˾D�ս	��i������d��נ�ć�<�4	�8�;=�����;�=�Ͼ��q���B>��s>��;?iĹ=aƽ�6)���7۾��0a��$�U��� 4������{U�$������=�a��?��U��>��\>����b>���;!ձ>f�=%��>��M=�?��>���=6��>?�=5v�=�ȉ>�	>�k�(�w�Ȯ<���&�zy�=�gC?yey�C���@67����Ҕ�1�>��?���=H�:������;p��7�>��	y��Z]#����</?�>���>)�=���$�ǽ�ژ��� �=!>�?�>Q�r>1E�=���9"��z<�B�>` �^��=�*@>Pq'?>4u?�I$?�=�l�>U�>q�l>�/�=ӷ=>��@>���>�6?iC=?�X3?�0�>���=��M��í=f�=G&U��Ϫ�OD��]r�,Z޻2�;;Ȏ@��<�g<�k==�#�<�	#=��;�v�<2
=���>�:?L��>��>1G�:a9�� G������>��S�7_�>���>
�?���>�q�>�C,>%뢽��ѾI����>��?>�\��et�����^�~>�j>Z2F?��.?����Z_���]=Eu�=+)�>�*?�I)?B�>��$>�˶�c/���࿌;%�D	���˜��2��0�>�� =�ra�
�[������+�;���=E0�>ɝ�>b�>:}A>��=�~>�Z�>�J>���=W�I=���H���*�˽Ĺ�<���<!_��ӯ�ރ�$�H����@�d%��=�K<y�Eo�6�?3�J?�,�<a&�hM5��R����0G-?�*�>�Z�>T�?��14���E�0Ց�
ԏ�w��>��8?�>Ҝ�A�=�.���6`�I�=rl�=�n�>�ޙ>��J����T��>���>��?���>*L���T��|��� �p��>���=6��0�?�>?4¾ꂾ�J3�x3T�n��f��;O���Ɠ��C�?�
��16�
���.��������Ӽ���>�?i�e���3>�G��d��)9}��<־�{�=$���@8�>�ԣ�c�׾�Փ��5��Y��~W��؇�=�Ǵ>�&;>�P�>xAU?��?;�?Xw?B�?Or�l�h?�->Z>�|?�T?�8?v�)?%�>��$��OμfY~=���0�����=;>>��=�vb=t{>f$>���=͉�=%d�����LX�6��=���=��<�@=�EC>jY/>w_?�4?����]�j�u/�,�������b���'>m�5���@V2>W��>���>��?R��>��%��6���.ѾH*�=<t�>�?V�>gT~��/\����72X���*<���>�ɤ>�������ϾYG&<G/�>7��>�>=ފ�>KÀ?a�)?�m�>���nH�?�S�m~����>�jw>E�L?r�a>��K<�ݾA�:���[�	�M���D�?a��j4��%ͼ�w�=V)4>�6�>�(�>��>�B� �a������K���T.���>���>��?�� >��ý�*
�,:��&H?��\���?��� =%O�����>����P-޾if����>�y}�6��ٟ���肿!��>��?7��?`��?	��b��U�?;�>�:��C�%�	R���:���P���
?g����ϵ�=�"�����&�:��{�Ӿs�Ծuv��`ſw���A(���+�:#-��+-��ӽ7���}���9��b�^����)=rㅽ}s��޲����Oƾ?,��?�wE>��J��BξF��Yi�ǩ����g��%"�۰`��}��F�߾�ټ�����8-��V3��<�߸e>׫�������nj�B�����{�7c>x�4?'t�0�ý�Ͼ9��X][>���=�#���汿�ȕ���/��*�?�c?﷒�?��{�>��ҷ��??,N3>y>�m��f([>���>?��o?��ོ]����䴗<Ln�?�F�?��>?�C&�|+;�[u�$XN�(�>��
?z��>|	��~�þ�r����?m-1?���>0A�������ן�>c�W?1�A�j|^>���>j��>��� _E��؜��Pʽ�Gm>[��; 4�
�f�f�2����=�)�>�g>~�e��)��C�?�%9�Mm����<���D�ѿ�:x=�=��3?*�<���>wb�>�x^>�Ͼ�oX�����(����x?Wǧ?W�?�YD?T��	*	�w�>fE�=�Ʋ>B?ֽ̅�%��#�E>�)?kF��WC�JOE���3?�p�?jw�?Wa?�	���Iѿ*����#��G�X��>�Ԅ=��n<DG���$>\m	;�� � P˼f�">'��>Cn>�\q>G�*>�EN>nz�=�و��$�=��x~���1��N�(��	#��e���>��G �U��uVؾ8޽�O齞��y�b���w���,�hW-��������>�?�M?F�>��L���̾��4���7��
k�ۅf�ՕL���
��p_�B�Z��N����پ>�>��A��>C�ƾY�=��F>k��=�"�>�P��դ�=�$�>���>m�*>[J�>�[>��3>��>iA�=>�>p,�=��m��v`������$�����M�>�p?�꾿���N�,�p:��6ھ$I�>��	?�M<Fi����!N��>�>��"=\1;��g�ˢ�<B �>%��>8�f>�4���ͽUpҾ��j6�Ro;>�M;>���)����O�Lm�>+�>F�ݾ��=�<>%?�{?�&?B`�=���>W0�>�4�>��=�#.>�>L�>�r?T�??Y�-?��>[�=�ℾɧ�=��_=�*���]�S?�Q��G��'��F��r�=W&I=��p=�ny=n��=Aх<��1=5���O?��H?�d>1�>c˶��@;��3\����=�[����Y�<<&?Iz�>wp.?�S�>i+k>s��=*;��ʵ�+=�.�>R>�Ks�a2��U5�>l?�!p>.�-?���>2#�Zx.�� >���>�H�>�<?��1?P3>�q�>g���$��mӿ�$�3�!���P��݈;��<���M���7<�-����ј�<�\>B�>��p>�E>��>�<3>�R�>�HG>�ф=?�=|<�;�;��E��M=�
��BG<�P�ԍ��7&Ƽ3��������I���>��:��8ټ~�?ء8?�x�>f��!��=C�h��S	?�:�>�5�>W+�>ot�vQ��VD�Vo{�k��۠>�?R��>>�a�=�s���0
�1��>���>v2�>L�>��Z��ɏ���>'�?��?? A�>�]y��������J�/4�>h�=�ν�?��P?��^-x�,F8���N����<�Y=q50�[֠�Di޾��!��F5�a4���w�����B
;���>ղ?�Da�SE�=�ܾ�������n���ڌ=���;�_�>�2�=�Y`�र�2p'��R;��>�Z��=b+�>#J=e#�>�iY?��c>�>��!?�?>Ⱦj�L?&�t�4�>D$(?*�?g�4?��/?Kpa>�R�e	o��>����,P��7=>7C>,zv;@�^=��=�-�!�>��=�d_����ӂ��X�I<`�l=�!�=���=uM3=)��=L?y2?,�/9�{�;[�Ҽ~��wh�=�Km>;ڵ��)��9=w^�>Y��>3?��>zVr�2����Ҿʏ�����=��?��?���>���<
v=���Nu�nE�<���=��ӽ�p���*׾�r�I7��uP>(s>r��=RG�>tB?.?��2?���O�p�ے[��w���b=��6=� �>~W�>�u5>��Q��Y�0�z���?�J�J��M`;6I ���=u1>	X�>ip>���=�7��2��=CR��`*�����<� G��7e>�l>�;�>a@?>�N>K�ܾHx@���\?����%�R]�����:g>��! ��rB]�-L?�b��d`�<�b��By��>?>5�?�5�?*�?���Sv���<?�pk>P6>bW���-�'A���)��?ڊ"<��Ҵ�7j|��K5>�B���<S=����U��
�-5ٿْg���1=�<�o����ž�Q�qz�b겾MZ���J�1����뾏c�jU��{����E���R��Z��ea?9B?���=��ν���}ɾ�/�FE5>���E�0�
��������Yg�����g���-,5��?�ChB>'�ľ���]��(᡾z���x>��U?�3*���'��OB�x���<<�D=�Xþ�{���l���ƾ�;�?�g?Ѿj1X�㰽H%0>���>T{��[�]���C��>���>PJI?Y@Z?O���W~���-�A=���?z��?�:?���=�	5�'��e�۾��u>t�>�@?� �����ܧW>�'?��J?�_?C8�*w��G�tu�>ˤC?�P���,>N��>���>����d���h�=��󾠈>�a�>�0���V���;��|O>G�>l��>��	����>���Q�=wE�]5����A=��?���x:�=;m�>��=o�#����rW������O?��?�Q?�6?#6��I���"���;�=b��>L��>JS�=�/�:A�>I;�>�A߾�up�����?"��?���?��S?]�k��¿/���6��H��ԓ>���ΪQ>���^=�9=Q�,��=v�=�	�>��_>/�>s>�W�=ҫ�=�+���E�X-����*E �;05�"}�BL���-:�iG���m��Tk�����������lϽ�4������֛1��`����q=S�>-�>���>0�>���7����ɾ'���y�QdD��􊾪����f�Q#��%4�N���<M��!%�jm/?h��jd�>�Ǎ>�~�8�B>S�>�%���	<3�>����0R?���>u�>��~>JvR>|1�=�}}>��=,�������E�:�[�Q�ŵ�:7�C?�$Y�Jԙ��3�i�ݾW���!�>y�?Y�R>D�'�ã��-wx��\�>E|I�<�b��Mͽ���*�>X;�>�(�=bP�����Tw���㽄��=e�>+�>��h�(���B����={ �>��&�&P�!V>��E?nRd?�&X?.D,���<��>>yx�>��Y=H6>5@W>��=b\?M	_?=�>?+��>��>�� ��)5>b�>�ρ�"�p`>�e����G�Ѵ�=a�C��>g����ao���=�C�>�y>��B=�����?9�B?�>���>��þn�)��7��3��@�u>�������>Z6�>�b�>ES?A?�_>��,���$�4r!�Y�>O6>2K��D��O����> �>-�1?;<,?'���M�5�[>4��>	��>�"?N,?!�>��>i$2�k���Yӿ��#�F�!�2i|��T��XW;�=�9'M�ӄ:�`/�R���q�<��\>$��>Zp>\�E>G� >O3>�\�>BG>��=-��=��;��;�"D�WqC=�����><Y�S��z��P�Ѽﶘ������ G���9�������2b�>HN2?��ֽ%���g���3��D���F�>bk�>�G?��>�����%$��Oe�)�B��$#�P��>��L?눬>0!���,>�'U�Wּ�*�>�_Z>p{�<�Zq>�e=��p��R=�[>�g/?��??����x������ ��g�>��<{��5I�?	�8?*�׾v���^�)���Q����!"�<-)|�����2 �L�/�����@��:����]t����<���>���?����Z�=�	�B���&����ǽ5>$0>zN?	��Y�e���ԾS^3��ː���/��:�;�>�>�E?�[e?�'7>�e?c�3?CO�>*�Ļ�6M?�~ؾ��R?`J?p�>�
p?���>T>���z?ݾ�d�a��(�N>�%>%�->we�<�^>����LKm����=���ϴ��@��՛�v�=�]a=�Ǝ;�>�%>�+?��/?�����r=��ް�m���~���$>��>��[�q�M���%>-H�>9O?��D?��>���<�O ������X��=�?��?�m�>��=y˨=0mؾ��&�V�r=Z�>fKN=�[��پ���������>c�>9+
>�b�>ϼc?,�?|	a?2���#�U��[�k/���2$>w��=�?�)�>�p��
��\��.R�Vg\�+w4�$�=ӝ���]�)�~>(:�>�XY>.��=�R>�^����ٽ|����I�=(��TD>G@N>Y�?��>A�=�������CM?���=F��?����>+��>����ξL�?�����A�[�����x���>�V�?e��?�mm?Ⱥ�}Z�o?��M>�H.>2�����Д�P&�m	?_�>��þ�XO��AK�����1�>��s���>��$�ɽPIݿ�&\��@���T�7��8����&큾�ʾ�"+�ҕ��P���ھ��Խ½���Y$�����پ�!z?�Qz?�ߌ��P���#�;Ҳ��G����>�׾�*��
���w������/?������	�{�%��"�c���F�� �ž����Άn�DIr��>�=��>W�$?���� �f�	��]�����>[ԋ>6� �@Ӟ���ga���?�mt?���&S�*)�8�=��(?5��>�>��a�zL[>J��>�?1x]?���>�������B��<�,�?���?��2?���v-x��d�b�g=�I?��&?��>aƾ���#�V>mr�=s9?3?=?6�57���vľ��-?3Bl?:��.�=��?��>�c��2���ɨ>��޽�����u��O�>h�
��i���1���V�;��?7T!?�ѓ�z����?@*������-��Q����<��=$9?l�0�	
�MT�>[�?g�۾Y�N��<��:���z?5�?�h?:�0?+�@�R�>�>�>��`>Bxq>�䇾�����df=��>������_��i�N��>u��?�	�?��0?βt��aҿ�Ә��CO��C�H�>Y#K>�d>%�c��,=�ͼ��f�J�f8�=e�>��D>�o7>�:�=�$�=�\�=����M%��w��|oz���P�HL����n ���m�b�I���������{׾jj��Pq��5"�e���.H���ǥ���ʾ�!=W	�>}ze>���>]��=x�>=�se�ov�����$�� �T�&��5��e�z��z����rU��~F=T��� ?.�APH���y>�Q��W�=�mC>�`>�dx=���=��x����>XII>�<�=�!�>;�v;F!>i
�=���<�\d�ۡz��/�L��9�=*%.?�޴�p>ʾ�F����	��t��>CN�>�=J�;�잿�Y�0�>�sL�G�پHX���g�=vE�>�4?R��>.�^�,���D־�oQ��=��>Z)>H���0������֕>��?�$��%���0�>T)?��|?�@J?��>��M�=�*�>x��>c>{
�>%�����=V+D?VW?��D?�>&�<��<\�>�\�=�����[-=I6�:W�;N�>j->����=u >J��<h`�=��_=��r=���M2�;{��>�Q??�>�]�>{����n�
]V��.\�?9�>M�_2?fc]>m�?�E?�*�>�}!>!"+�C4�����2�>��>>8߂�{�����㼈�1?���>��0?��><T�.w �;4>�~�>��>L�?M7?�Z�>�T�<���Zk
��ҿ�	��VМ����M�S�{F������}�kV<sž�j�!�N<Y��>3B6>0�->��=Y��0��=���>��E>%��� -�=G!�=͒S=w�m<�2�=-��<�L�*'޽~��Z��*�����d���򇗻9C�<<<�?F*5?[3���_p����Q�,�ߞ��:%?zK�>̶7?J�?��<��q]��b�c��/X�>��l?zk�>�^4��A6>*Hn��+��.�K>�K�=�ۆ>;�>�:<B69����>G+�>��> ��>��f=������po��O�>���=�b��ǒ?7�C?4R�we���S?�h%9�a��%�:�� ?�Hش�����6��Z<������=n����0��?!�>�ϲ?���FN�=�?���:���:>i�x��=��J=p>�Ჽ|������B��5��� ��V�=�P�>T7�=Y ?�=^?z�>[�%?�)�>�?����;?� V=�s�>���>�A?z�'?t|?b��>JŊ;��L��=kA�M����%>��<�!~<m	�%'x=B:�:��<�	:>ٻ�lی���=�=�愾8�z�kϺ=;��<7;d>b$?��3?AG��F���>�!�I�>h?@>���>s�.�i`R<�ڇ>I��>�?��N?.B�>���y�;����]�����%&6?��/?I?�W����;����"+:>�e��t+�{6���	۾b*�<2�:�bc>��>+��=�||>�y�?�E;?}]<?��־?����"v�����>�l�>�>�X�>��~��㜾�徣<���d�>��s��>�y��S��<�p�>9��>��>��=_��H�Ŝ��T�ؾE��=Bֽ��>�t�>	��>�:�>�;R=E0̾�E��]?�m��Y6��U�=};����
>�1>
�	�����ԅ?6_��5�z`��nv�K�6>D��?�3�?���?���pF^��x�>��">'K>鯷�������<���l��>�*>wӆ����$X�<*�9��(>�%��Ӿ�;ƾ
^���mʿ{Fc�h���\�.��.K�u��5���ɾ"|���{S��p7�m����ξ�r��	)�I�V�2#پ�`��	˾`{?(j?[�1<�����= �3�Ͼ�iy� s�=�S���;��P�������̾)6Ǿ���{��������ׅ���{>�똾4�������i+;ْ*>�)�>".I?���V���:���,�O��=��>H��(������/�{�}?�4b?Ô�L�?����o5=��>��=�7B>Cy���D>�M?d�}?�Fb?T�=/P��UK���>c��?�p�?]??�]/��=���|K>��:�>8�?��>NX~�Wᵾ��ʽ<?��5?v	�>%<�/䆿T���3�>��`?�#L�GXJ>�<�>K�>�맽DÕ���*�X���N/X<w='>��ټ� ��Uo���K���>���>SJz>��w�TZ���7�>����M�	1B�����_8�o�=���>"a����>1�@>f#�=%L3��=r��a���Ģ��VK?�D�?�vG?1�j?9<�V�۾�ݽƜ	>�?�|>H��=� �=�ET>��>c��Ksd����вH?���?7�? M`?�#^� ؿ�a��eφ�**z���I�F��<��>���B>�<=!<���(��=�_q>��O>(Eg>�wK>m_�>0ړ>�@��ʷ�0���L-���tM�� &�nd���X�����i������V*�����yB�{~ ���n��׋���<b�>�踕�� ;>�{?;?]ı>�� >��s>�E����W�e]Ѿ�& ��봾����{辤�Ͼwⷾ.�S��C��&ٽ`�㾄�?��>� \=7c�>�4l���>���=0'�=��%>Y�!>��=X�W=��=�ق=�>X�>X�=ց#��+=�9�#���>�/����u��=1%}?xӈ�����^��M!��z����>#��>��G>�0�۳���4��r�>�ջ��fs�a�s<�{ >��u>�!�>�Aս��;{9���_�������<���=���<eNg;������m�*,�<9�>Lξ��=��l>�)?2t?3?�=��>�7a>Fے>���=��B>sH>ڈ>i�?h0:?h�.?b�>�l�=B`�>�=�H=��=�U�f�䩭��������~�<K9(�GN=Օo=�,�;�:=��7=㰦�L<pR=�o�>�G?�r�>W�>�₾� �������^����֬�#�	?�\>̏�>*>>�'�>� }>��=�\��拾#��>���>�P��)M����Y=���>��>��f?�W?{���s��<��=�3>���>c�;?�#?X��>"^��=վi���ÿÝ�U���\��ýQ1�2^5���w>D?>�������	�����=�>��,>T�p>��>.7>�>Kp>%c�=/���A��s�;�ˣ���=s�8�@I=��
�}j¼:�<�~����A������ت�ҫ��^3�>3�8?��
><�< �X��.��c�,��>��?"�>�,?@��)K��~p�l�C���>`:?�uX?�wc>O�?��%�4��>D��>��=�\�>��[>'x�l�����<�:	�ʡ�>&L?�ύ>�9v�	�K��x�R��l�>�ާ<<7��y1�?վ�?5���G�fJ��NJ�}�4�ZC=G4$�v�w��!��f�8�ɊC�Zw����ɾ��p�P�>}W�>��?�R�_�@���_����i����PW��8���	?�<=kM�޸a�����d����?���H��>bL�>�F�>�!>�Z�>&#S?�b�>��?X�߼ʊ�>b�.>�b?�C6?�>��>���>6o=?��=O�`�y�U> JL��~���=�(>>�I�O����O>�4J���H�(�b>�O�=�R�<,f˻��=L����TD��V�=�>�K+=`;?(r.?�f��9�n��<���5�� ��=&�>�.��@F
�B�&=;��=_'Y>�^+?��>��r>�O��
ܹ�Z���8R�>7%�>��?��$?��.�%��ߤ���<�h>��t>��
�ץ̾hW�h����[�d>�m�>��>Z|C>lCr?�E?d+?�2n��b�6BW�OKH�k����'���]>"E{>=��=l��28���q�c�2��0�p=	�j��o�;�>d2>�\>��>��Y>� �=�.)�����=S;<(�>c��>s��>G�>�0&�\ت�GB澞�E?�0��c"�Ǿ��-��?>L�ٻ� �=�=�>�>���9�!�����q-��@$?~��?� �?��7?��L�>8���˽} �=�a�>~>�0I>���hyĽ�a�>����,�6���qW>Zf�>|��>�#����ܾ]�J= 2ſ/3�IGy��>���&z�ݼh����=+����eb=𸣾�Q��AO��!-��1�Q����oދ�W]¾!�̾��?l?`�[=`C�fn�Q�I1E��gf>(���5�����5��\�2�������A����t��pU����}��>�Sھ}f��5L��Է�j�7>�x�=���>�xžX:<��5��ν�͛M>}y�>�;����y�{��/����N?��.?"�۾)�����ۇ>ӳ?��B>#T>��t�L��:��=��J?�j^?�B�=�2��
^���*�����?UҲ?�@Q?2�4��I��̘��-G=�!S?9?���>���մ�tU��[7?!��?�s@?��"�����y�@�D?�F0?�X���>���>�}�=]���ָ�?8 >R�Ͼ�E�@���醾?�	�I�� <�����b��>W�m>���$/e�{�>h��)�?�G�X��}׾֪�/��=�u�>�����>n�i>���>b (��|��W$��콇�M?�/�??��?�gr?�&�pN�����a>V\�>���=B�нc(��J�>I�? 
�͕r�v�� ?���?�0�?2CY?_N|�"�ӿ������V���D<�=?��=4�>Z�?.�=�k=��)=X�V=�T >���>�U>1�Y>�Y=>��:>�#*>�H���"��𥿜����T��� �:���s�=���cC���
��ቾ�ޢ��.����Ƚ�ō��M��7�a��
�Ҿ�3Z>�f�>��?I�>�5i>�C=7�!�R��k� ���͏���h�6|�2�Ⱦ�Ǿ���=��=:
ٽ��㾯�?&�c��]�=�>���=f�>��=l'<�L>,�=���=`�	>�h4�b�=ͤ�=�ܿ=�9>>��=�3x=�J���{�÷J�;䖾ŕ=��[?&4ͽ��_����\����S���N�>!G?�)�>7��f����t�n�>�q��pq�4z�m�=6��>d/�>ƃ�=��=R���½�����ؼL�J>ٱ�=�t��S�H#��8\s��.�>j�վ�=�#v>�-(?�Ev?v96?-�=��>*�b>q�>���=h�J>��Q>{��>�h?Up9?e1?W��>K*�=�^_��=]�?=G)@�,�[�e'���+弴 '�G^�<5�2�tC=ybs=ڹ<$O_=5�B=���Q4�;�4�<Ӫ�> )=?!a�>���>��3�zP���6�~C���=f9����>�&>�A�>� �>��>��>�AӼ���,O��8?i��=�P��hl�Uz���>��>�O`?�yy?C�Ծő�=iM�=4��=[�>��8?�#!?�e�>�%�ë���"
���ο	/�!��(��ւw��ۊ<�g:�� =�4�;�W����>#=�WV>9B�>��g>�=>Ũ.>ye5>��>o�D>MK=	�=�!����^�&���v�=��;��|�<���r���5弁�`��d~�v��L4�ؠ�yQڼ���>��?R�.>�4ʻ\��������j��>�z ?�Y	?ߛ>J�ɽ.x ��W�/K5�3���D?�VY?��]>q��P�����>�q�>��>��">l�=6���,2'�J>�򑾘��>C?M��=@�_�(cI�/�������}>�m�9�6��?��R?����F+��`�!�2<�\�'�:%>u���e�g�/�����,���-��4оW�ƾ	���ƙ:>ٮ�>�?�>�����;�u��xj��E�]�����>齌�?�V=�+�$�������_�0-���&�O�m>׺Լ�?":?��"?��?O\�>�A�>%E�?�?���<F�Q?7g?���>I��>5��=�s����$M��>�ž�Dh�(�r�ټP>�Q�=	{���=>R$4>�d;�DE�;K�N>�����{�iH��i��s���*GY=e�/=ױ*>�jP>غ?�?�d��͍��KS�ק���>��=��>�rŽ�t����=-�%=��>��?�O�>-7�=�};yW�Cd��۵>-�>
G?1�?������m�""��̅^� �>_!>sX��i�����̟��,���b>�w}>O2>p�>;�u?F�W?J�N?"K��"���6����WXͼ�W�=���>��>Ι�=��̾^*�,�V�+�V�!>#�(F�#���hϲ=��}>]��>_�`>�B0>¾��U�\����kO����>�H��.v�>u~>�j�>�B�=�������Hy�i�R?�q��@������ ʽD�@>�;��,>U�4>7��>��<!~�� �����<�v?"C�?t��?�\?�gI�s3���^�<��:>�L�=Z��=�<m�I =c��>m>�����(�K>���>��>�Ћ�m����t��+_���=п��*��¹�.��@j��	�žM��~>�?y���l=x����ང�'��Һ�m��t��B�z����������?�WB?��+<gx����0�he@� ���Ad�>.*���4=^,���
�בּ������������l
�5�J����ͫ>�c��|�\�i��H��f�=��>�C ?-3ھG��h�+��s���>���>�9^�ݒy��n��6�p�3�y?��/?|W�̨��r��(>+0�>���>d��<�_B��M�[5�==H?�Db?�����G���׼�1�?rp�?��V??��J�[��vɾ���m�/?f?�>ހ�2m��O��1>?�8�?\J>?7�þ�
����'	.?�2.?�����
?���>��{>�`���T����1=>�ؾ�B��	���4�=�P>����ф��0�sz�>��>c�+�Z�޾Uƣ>����D��BR�8;�����$�=D�>�# �"��>��>)�=��5� ������$0���E?2;�?.�x?��j?���D�����\>��	?��7>h�Q>8���>X��>����Aa���8�7?v6�?�+�?�t?�s��Kܿ�훿{���;p����Y=Q�=n�|=�O)��\G�P�\�u�P=-'�=���=��p>�<>HM6>�T�=8��=x̕=Q��R8��������8S�=��l���������Cy�Q��.F��Ɠþ���%8L���2�g�J�9ȶ�bq�ೠ�+|>���>B�	?��?���>��
>I���5o3��,������\뾼j����ƾZۼ�����޾���=��.>5��L���?2�$��o'=�>9�(3�>b�c><�=).�>@��>.]>">?>�B�=��#>]]>9m@9�>��<�.'=�RM��̇��g��P�gMU>�rC?v�3�Ŏ���#���{㞾�ܴ>�б>n�W>} ����y/���`�>!�ӽ������<!q<�Ӊ>���>uB��~�m;1�_��~������Y5��G�=�v>�6�����X��]x�=*X�>Y&ƾ���=A�k>�J%?KAo?Fr4?���=�e�>��i>?D�>��=�E>]�J>�~>n�
? 	7?@�,?ot�>	#�=!c`�G/}=i&�=��B��F���ܽP���W���
�<��5�ȕ=�=I<I�H="�z=]jݻ���;[O=	�?<?o��>'��>�����4�.�_�꼇>P=�_;�A>�>J�->�>�U[>��
?�.�>��2=w�	��0���I?�]>����V`��� ��=C�>m�Y?N~c?�Tn��$۽{�;��
>R~�>�l4?�&?���>�������w 
��ͿHC���%���	�|㢽?	���B�* ����D����ý�J\;�
O>� r>Rvh>�R)>��%>T}>��>8�V>��4=OI���{�{�R�Ἠ-�=�����}=K��X{��'~����]����Uw�H�̼�����	��� ?ۖ?��>��=@����|ƾ06;��?Z��=�?X��>
;,�������K�(�}*	��I?�L?��>�x���t�<��>��>9��>:�>q?4�)V=�_� �7H�*����>�?�q>0�^��PT��D���K����>m�=S�����?bOO?_�Ǿ��q�7��j'�3K����=��½�=��ޥ�-���"���ؾs*о|t�$�e>�?�l�?"m���k<Ñ׾����ˈU�fJ��=�>����(�?�==�8�Cϊ�dh���C���Z�%}�0�>�1�<O?:�S?L�I?��=?uq?{�>?�o�G�?��ݼ��_?%{?�?24f>+�=q�m=�b���S��,:�q�׽��9��M��x�=���=F�= �
=1����TC���$=��꽥c��Gl���=g���9z:�~�=�$'>U@�=.@?J?YlF���˺}�׽����ݦ�>�J>���>��<���#x�=��>�]�>�?�T�>j>�}��������*�>`��>�2�> 0?u�A���"���Ӿ;߯����=�S�>'gs��Zݾ%H.�����Rｩ�B>��>/5�>�WA>@]y?�1\?��2?0⽛���N���\S(��=s�>�
�>̓c=�m־-/�n�[�~N�M�2�(��Fuc�Pα=��>��$>"��=��A>RX>V5�g�=������n>���=B�>���>�#�>�>�	`�k���m��|�O?�=��*�(ѾB[2���=��h����>E;�>�Kg>���*������@�YG8?j��?�9�?C�?�X"�m���w��w��=K��=̲��">�Ԍ��{����ļ[>�f�����?k�="��>�B�>A�[�$ʾ�@����� `˿CL8�O
_�[�C��m����p�^�@7�=b.>�u�I=6�׾:�w�=���>-:LF�.۹�p�Q��6��R5龇�?�\�?i��P���"����1�Wa�>ܨ>V��W�
>���y��-�|�z����V������Rھ����D��9�_>b�������p���ؾ=ꔽˣ�=Y�T>�!��܈�-@��Q:��AW>w{�>3�6�e|r�����]�/�h?��!?H#߾����#> 4�>Z�>�b>.���;�������>!%K?�)m?�9�=h���G���Z�;��?�?��P?���c�5�o��Yκ�m(?���>;�\>P ��1���~Ҿ:�i?�E�?_�O?����E+쾡K6?RJ�>�m� �?�?HB�>��ؾ������=����֕=_`<3Z=�=	�ľ��������>\m>A����׺�כ�>���h?�ʶZ�N� �1���`�=8��>������s>�{�=}��=�.�V	��E���{i<�V?{��?EPC?��g?W�߾P+������8V>���>��>�|t>�ļJ�>B>��p]�_�Ͼ�)?L�?U��?�eV?n�_��׿f���i��2g����=��l�=D8<����>P��=�/u���ػ%�=(�;>Cp6>ο>Z�)>U�>�>oT���E�����b����/B���(�MA%���#�c�On4�]���;]�۾ǳ�?'��*ν�\>�a�м񴼞����eZ>��?�t?~!=��=CI�=+[�s(�~Ƚ��;nվy��/�	��侤|�@y=�>����K=5�9d?c	8=��;���>����a��=�C�>x?�<��x>��>�/='>>YQ�=�F>%+�=6�>�_>\��>T/�=j���h3s��/(��㻖!t=��X?�9;�{���d�þ����'l^>:\?�cn>��F��~����a���>�:��[���)�Yy!=`�>q�N>��0=�»�P>����j	��b/�ڜU>e��=(��=�>(�쎾��=���>P'þ���=?�c>U�$?,bs?�n*?�.=���>qC>>XN�>��e=I�B>s�j>���>�@?K53?Fy/?(N�>M۾=�c]�'b�<���=�M>��Wt��_����<�ø�����v����=B�$=(k��g�c=��=�����f㼾ˍ<s��>VjI?Ps>���><̧=��:������|�����h_��@�>��=�>�-?#??�ژ>�R���"`�=.�>�8{>�w���s��> S>ـ->��&?1O-?�.�<6�i�D��#�='��>�Y?���>��i>�?U<;�=�_�O���I��+��C�_�M#���_;��{��>�>f���
�T�\�F��P�<� ��2�=�Y�<�\>�>���>$<<�w�=�BU>\v���i3��v�=�)��/��斥<����n�Ҵ,�M�Ƽ��rC��8ʽ������O<�?�k?�w��Ku<0ݿ��	����;ݵ?��?u?&�'?���=�׾U*y���K���뾋��>;c?)�>)�<Q3��������ľ.��>q9�>|�)>�r�>�&�=T���j�>���>/�:?�x�>l�9�BMp��0���>��=��R�?֊F?c��GV����Vf��0�����~]����� ܖ��v�jn��P�<����/�<>�ʱ>��?�g��ռ0=��P��ԓ���m�������*>���4�>���[9+���`�䖊�맃���н��=n��>>	`�/>8?��d?2�[?6hA?1(? \�>�)��Z~�>ͱ�=!)[?���>���>��m>�ʝ>��&> ���*S�;s��~��>�<��u�=����3j>�lt>�H>)`; �s>��-����=��<� <�m<�Gw<��_=�^�=�:>��=�	?$�?L�u�\6�&��<�+S���)���`> �>�lݼ`����Z������>�)?y ?tr�='.�\������I>4?��5?9!�=�����0K>�cd��fоa+�>�O�;�cؽ5���x��ܾP��Ӫ�>�֯>0影�%>�C�?1�O?�Q?�CS��R�c�2���������}=g?��>	E�<�^�J(���N�^�\��B��c)�N����E�=�GV>Ĝ�>7�>܆>�m�<$�6����k(��n�=�$����>�*j>��>�Z>��i��殾���n�@?�˾+�*<оZՁ��=�g�=�M">5r!�Ɨ�>Р���y��ٝ�#����>z��?�p�?+�H?n%�4~�<İ��Q�N>��_>��=Pg>�hO�`2�.�>���=#���J��b�>R��>O��>92�l��h&���
��1���S�����'F��.H���_��獾ς�j�&c<�]ƾ��Y��H���,4���=�D�N�q����٦��U���`�?��Z?W�:<����d#�>��zo��z��;M�����Mu��,���t�d���Ӹ���Ҿ�#�_�
��Ͼ6�>>}�;���Iv�t=��o�>��ջL�?�ѾIˆ�@�-����{p�>d��>Ro�e�t��ɡ���;]E?`?6����Ӿ���;��>�D�>+,�>tp:>ة���}��rR>��Q?
G�?�a[>�M��ԅ���r���[�?.M�?��Y?�V1�C9!���㾅�>&(g?<D?�U�>2�z���(�Ey�����?(-�?��?�n
�m=����&1�>L���z��wK�>�F�>���=4E�ź۽5�=�zξUf��V����(C�Wg�>>�F�#�{�їS<y\�>��>�1��,���^o�>o���P���b��Ӿ�.����2=� �>~�
٧>~&>��f>D�<��Bv���FX���>?���?X�j?��`?ZF"�=���Zý���=��>Ǖ\>�;|w��xY>� ?Y&���g�w�"�^2%?N��?3��?�i?����ٿ�f���}������T�>�<��b> *�����s�����=|�=G�$>ˡ>Gw�=bnA>�b>��,>/��=���;�+���/���]��>�[MҾ��V���&���hq;�9b���Ǻ���)[���l�g�	B����X�����>���>��?���>o�	>�؀=��/���Ծ�R	��S��'��qϾ	� ���tg���ɰ���=p��=�͐����$c?n@��Wf�=���>:�G����=K��>Z0�<�Q�>�/��Y��=Wh<���=��_>I�.>I��;@�c�A��>�`S���w�.]h�)le�I�+>�e�>&S?z#>t暾ļ���I���ʽ���>�?��a=, �����萿q�>�R��)v��������=YƵ>��>.%>Ԥ�= ���:��aԽ��U=CA�>qG�>-��=�/���"F�ե����>0�׾�Q�=�Uu>��(?k?w?�m5?γ�=��>�a>0�>�=�=lL>�(S>���>+?�79?�1?o �>Yq�=	`��G=[=>=*>�OuU��ذ�����&��~�<�=��kI=AB�=��O<y-]=ױ/=݅ؼ̀�;A�==�>¿!?��>��n>��Z��=�V�V�ǽ��r۷={��k̍>쯇=�w�>%C>t��>���>��=��澱�p��c?H��=
���|��T��S�>$Ž>鮂?R�[?ା�}ؽ�oG>��`>H��> ?�*?澍>�<�Ak�[���ҿ�t#���"�$��]p�*L:<�	:��8��q�;�j8���8��<=r^>cx>�Xi>~�7>�>4D4>Mo�>�xG>'��=��=�ǻ��һ�^O�k�C=f���<<%N�l	Y��i�Ӕ��֌�3YW���k�l�,�2�P��?�?�K�=\�*�"�\�]�ھ���O��>&D�>�4?O��>Eܥ<�"��e��1�l���^?��c?�?�>���Mt�<ɇ>BT�>��N>k��>��L>A���+��q�7<쏕��?�?	�v>�"\���R�C��il�# �>���T�馭?Ev?׾���l�"�� O�,�3�`�>�ϡ�[��ԾZ�>�����oܾw5���!��Z�=&��>=�?�v;��w0�X��Pٌ��"F��;f��s%=�(�<O+�>kMj=�;���`�4龹ݥ�z�A�����55�>�I���?��-?K,]?��S?�?p�>n��W�?�H����k?���>�?8�r>W��=�\<��y��&H�2�Ҿ�@��/���I���K����z>XN>I�M=�^�=}�6>��=β�R� ��.V��(x��ȍ=x}�=�~=�׻=�,�>֯1?��
?%I����҈2�U��31X>A-�>�>b[M>���=��5>�p�=���>�?sM.>�0�>`���.����Y��>�J?{�?\��>3����m�¾VA��x�V>_�D>�'�Aܾ�4���ؾR���Io>ʻ>�>���=gMz?pW?�rG?'�f��!��~'��	�4�Z=чѽ�V�>e��>���=�z��e�*���N��ME�'&I�C~����&=>��>y��>R#t>��>�q�v�������0���ݐ=U�����>���>��>��=����蛾�
�".?%���B(�&�`�6>a�h=��ƾ7]�>j�/>4>����7����嘿��A���,?�3�?���?K�D?���i�<[���>�,>n�f<�
�=Uˑ=>�`=�t>V��=�#��Z��g�>�0�>Ԁ�>e>��ʾH����k��#οh�P�bdM�jC�����}l#�}�O��n���Ͼ�����z��\���q\���r�������Q�V������úh�U3�?�dd?$1e=���P9��n�_�ξp*�=���@=ͅ��h��H��'ڦ������4�"3��#�/�����">�d �3ي��Rn�����TM>�F
?�,Ͼ01%��%��;=!�Z>Ч�>�+��6�m�U���N�^��dy?oiD?�,ɾ�uʾ^���KI>� �>n��>�w>ᆾ%���>�YL?ۯ8?g7	>���?���=�v�?/�?^H?l��
EL��Bľ8����.?^!?и�>���	�6�Ѿ`!?O^�?ZF?v��ԩw�����?	�N?щ��M?�!?,�^>~T����Ⱦ@O���/���1�?7�=�K�,�>�~�n����1v�6n>mܮ>����.�����>���<�m;�Ȕ(��ꗾi��=tA�>���0OV>��>}��= =3�dxu���w���O�<�;?M.�?׿h?>�A?��Lž�?׾�o�=^�>�I�>sa�=��9��B8>�
�>�p����d���Ⱦׇ9?���?}�?f?��V�&�ؿB��ؘ�����	5�=� �<�N�=�&���j=���=-t��-���Y�=P=�>��>$�B>���=�b�=�'>"��H
!�K�j����B��C(�����ا�\��:yf�up�4���@e��k��80��k܋�nkl�	 �������>B;�>F�$?��c>O�=�>/���,�����i� �=�Ū��*��	����1.�M(��������=�������?���b�>Ѥ$>��a�A�н�;?M��<��s��9>��=�l�=M�=`��=�E�=۽�>��P>�&>�[�����=n�?�O�	����>A�J?n���`߽��9�����U=�>z�?�7>H�6�����m�o�a�>V�F���ܾ9߶=�:�����>��>�O>K���� ����2����=�.�>��>�$p�	�������D>�0�>ߜ��� �=��>�"?�_\?*?{�����>+��=U�B>�>2 �>��T>Ȕ>c��>��B?��8?���>Q��=�l����=;��=X?;��YZ�H+J���v�y�܀��eL���n�;l�=,v�<�W�=h��=���=��^����}	?�g?�S�>���>��q�9�)�?�V����QF0=�n�<�m'>�FR>}3?�_�>�>pb�>Ϋ�=���9.�p�>�>>\�k��#��g��J>�)?q}s?���>��u>�>��`}ܽ�"?�v�>��O?X �>A; >iAT���mӿ�$�7�!���P�'߈;��<�~�M��S�7g�-����?��<R�\>4�>[�p>kE>��>�<3>�R�>�HG>҄=!�={9�;�};��E���M=�	��BG<��P�C����$Ƽq������S�I� �>��9�39ټ���>�{?)��=r� ;d�C�^�Ծ�Q���>R~e>_��>`1�>���=��4�_���:����T��>m�P?H��>z����T>��%=Ъ��UW?��C>@�ԽC�=�h	�~���'�)�>�L$? �}>O�w�����\��@����>4�=�5��ό?-�e?�)�ڗ����
��C�Y��V�=:�ͽ�EW�������N�:�F���AT~��|>�I�>��?ӛ,�{L�������Ù�1���R���H�=��=��>��>>�T6�M��\���N�����o��=md�>�[R�N�?�XB?�7�>ދ?�+?��=�Y�x�J?�Dn�z�>��>H��="�"c>$�<�Q�=Ꝝ=�@%>�p���ޒ�T�/=}lQ=-W$<c�b=y�]=/l��ԽG�V�(v�=��%=r~ �Y�ϼ�4;=8*�<A��=�;�<���<r�?ڔ�>�Sž��S�݊�)�߼T�=[�=�� ���<�ٿ�v��=4L�>�?B�?�-�>��D>�W(�i��O�U?�>�+�>�F?��?�*����=_	���T�S>�a>M���U����
�J����=��=Y��>�_/>�<t=�,z?`qh?_?���=@�Ѓe�(����1�>��=E+�>��y>u+���#���<�:Sg�7E���-�4>M^�/Ń�C��=�26�1�p=]=P=�a�<}-]=9�=�*�=Q(�=��>5�>a��>*�*>��=� ���Ѿ�QC?��|, ����<��N�Y��>��>��z0?=m�Zt��ګ���k뾹-=?��?��?lVr?�@���4>>�
>�`��>�x~>08E���wV�>��I=�TľŽ�z��=F�Ƚ�M>�&Ľ��˾�YQ��"���t߿z�-��iۼmqp�����?&8�l������Ѿ��*��ꄾiCN�G����fo������Ⱦd
���09���۾]�?�	?#�,�����kC�����K����Ҵ>�׿��P���pʾm�t��D���s��t�>>־?��>���'ʾ�J�>���6+��gu��2�a�C>�Ն>��&?y½��r1��=�F��#r>�¥>��۽��b����E��7�1?��+?W�z���lF>=z>vB'?�l�>�F�;��%=Qk���[�<��o?�^?�?������-a��T�M=��?�̮?�a?l��4�]�w�J��9J��M?]#�>��>r�=� 2�����zf?�=�?j)?�վ22��O�Q��M?㿳>��4����>P��>W��><��H�� �н�亾�m�8q}<Y.�>O>�兾�6���=��v>)�>�6��-R�>Pq��9��@'���$��Z�GC>/��>XB$�vP�>��=j
r=-�A�Lzd�����[���C?��?S�a?��U?Q���J�*ɾ9�^=�G�> N�>��9>\ҝ� >(�g>o+־��W�@���G?i.�?��?��r?8�I���Կ.؏�����ݓ�ܯ7>���=
L�=,J��g���=i�=��(;w�1=�>�#>�=g�=���<�=Bʃ���$��ؤ��Z��9�2�����_�:�������|�Ӭ�0�ؾt"��O�.���ֆ߽6]l��W��xG������f\>LV?��>X6�>�r�<j)>e�����گ����b� L
�wT�[�X�Ǿ]t�d����Ũ�VN�V�y�{��k��>P�!=�/�=���><N̺V
>��>p����=d�+>r�=d�M> �P>y>Y��=+`�>��>	��>w��=GV}��rl��K�\P>�oT�=�P?o�?�}cT��-�0Z侨㴾�o>�>�>��>��)�����+E��s��>����ꢾcQ���2|�Pە>Du�>��=sꞽ
%�SS�yA-�"/�=��~>�"�=�>E=םi�G_����=���>��˾j�=(u>��%?,�t?+�5?��=ڣ�>_>��>���=�ZM>�uK>IM�>O?o6?�.?,#�>r�=
�[��j=��2=�C9���]�Ƣ���b̼�O ���k<$�!��F=?�n=P�D;�Zl=5=�3ɼ�4h�is =F�
?Y�?o��>?˾j���<��B�<@:=��i�KV�>���>���>Db?�	�>9o�=,�������.�8�>�W/>�f�	��hF����>?�"?q�y?S#�>a�>(�1#��눽���>�>��\?y�H���G�}��:����˰�\#�|F�9O�=�$W��*��CNQ�F}4�J*D=O�׽l'�=�6<�(ʽ��۽&�2>wc�=�0i=��>[��>	�>$��=���=�zڼ4t���=/�O>k�w���<����kl=�1�=��=�f˼�Ev=C��;���=�[@=��>>{3?��=_��=�紾���&�M����>2�>�?�?�k�ە����W�6&��`	�
��>;�6?Ų?��<�z�=p/���<A>�0>���=h:�=�߽d�J�X(>�=�>b�?%�V>��!�3���U����+��>��#=��ֽϗ?G/Y?�n�������dN�� �ף=%��Ҳ��L�¾�`�Y(+�R���h뾘�M�C�'>Z��>�U�?��j��x==*L��Xڕ�\rz��]�� r%=)G=�z�>�1>p�%���ْ
�ڝȾk����=��>���ʶ"?mGO?�k�>��?_z�>ĝ�=q>�2Q?�2->�i#?�E�>4m<����Qb�>a��>�@;|�Խѭ���\��������=�ǽ��>p>wS>���=*ފ>��F=�6=귣�b���8%<��缃�=/��[�=�+?��?H^ҽ�5	>�Z��@�<�g�=Y!ƽ���=(���3#��Xc�*~>���>�_?K8�>ܢ�>EI����ξX4得w(>e�?�?�A�>\'���;�� ����iʻ��=�ڈ�0e�o�{��L�# �>�6�>c#���4K>��}?�[?>�?���#/��|�����->��=t5�>�|^>3��q�#�!�d�Ź>� M��|�=�7�Z��<s@N=�g�=Ԧ�=��i=��>_)>L4���=**0>\��=��>L-�>��>�#P>�z��о�_��F7F?����
��k�F6�-+2����>�j>o����C?�Ɲ����:�����ʾ�$?���?�H�?u^q?D�����=x6$=c��av��u>�L�>C)���u�=q�>�P�x"������f�>�?��?@�ؖо_r���Q�^����FZ��� ���~������z"3�&�����TN�=�ݾ��1���Y����ݱʾ�^��rƾ΃Ӿ��/���?��L?�n{>�b`��I���	�oMQ��Y=E]� >���q��Ծ��j�;�����8~0�Me�����3�>�7��(4��R'��������>qO�=npY?/C�x(þ�?���8�X��>�B�>������{�u̔��y�>��\?J:+?�������|'�> ø>a�0?q+>�C(>
����:Q�<5>�Sq?��?�k������	���\��7ӱ?�3�?
�V?E�߾��}�G�9�����Bh?��>i�=<7���;��x��!t?��?^�?7����ؗ�=��T6?�C>��X�%??$�>[�7<����]̾5�3����-���;sQC>��=�#����������xܬ>2+�>�ؾ۾�4�>T��G�?���X��f���B�a�>{��>Ȼ����>�;>�f�=�O9��}u��ǂ��f�!-?�Ţ?<�`?c�K?�ھQz�������r�=���>]��>���=_ ��ې>�w>��%~�\7ܾ:?6d�?m��?+P=?4�J��տ{������������>U��:/�=�i��)��y�=O(�:��P%���,>6Ch>���>��!> ��=��
>Cʃ��r$�Z����Џ���A� ��S~�ᚷ��2�=�ڽE���ƾg�־;�ݽ�f꽞��<��"�h���y�1��̾���� ��>���>|�=����F�>��aGԾwN(>I�M�)]����=1��v�����'̇��Y��Q/>-x���8�>�6׽�{�=��>�>�=�P>~��>���=l�=<��=x_A=��>.>O#>�b3>V]�>�>3^�>f7�=(��*7q���>��O��u�>`?�{�7��ü��ý�����z>>v?P�9>(1#�����X��O�>7�u=Js��_���r��a>2�>$�=���9��<Lz��=�x�7�<�U>Y�=>�|�="�Z��� ���S�K��>DľL�=f�\>(u#?�q?L�-?�@�<���>��P>;�E>�͹=�R>�c>�1u>M?	�>?eA?���>(o�=��j���J<��<�%��I��q���j4�Xս���;.�ɉ=h�/=*��=�s=�F{<�:��<�x={2?�~?H��>i��>>���Q���O��9���x�q�N���>�n�>R�-?z�?���>��=
<;�E��Q���� �>�R.>�9L�i�4����;�>�U�>=�?'?!�qx=oj��x�=���>���>oY?��ɼ��>Q�>��	���¿����g�0�D]?�Sdp��dK�\���q���R�h>���}3K���$�B�C=��=Ù�>E|>�=X=Q�=:��>y=N@�=@��<��2ƾ���G���B>t?(>���=�s���=�D���p��J2��:��x�½<�������^?r�?�p��l��<t�߾�Y��{1�;��?n�>��?�?� �=ݤ���u���P��.%�| �>g)8?-=?GA��H��Y^�v�,��G�>C��>���>u�=��U>�ؾϧ3>��?�?ļ�>���+~�����>F�:=�!�ϩ�?�U\?���߀��R��OG�����cg=o��'	Z�?}���� ��6�0��*���'o�!	�=r�>�?:�~�P�Z=R��C嗿i�������d=n��=��>�ZG>Jj8�`����e^̾��H�KǴ<�_�>�"�<P?n�?!?�c?�S�>$Kֽ/|2��d�>��,�?nv�>	��=�>u�^x>�<�=s�> 3��Ps���S��!G���Q>={���{�=�10>�-�=�0� 0=�FV=r����/;�$��X��r�=�Ä=�>��=ȹ�=_?7� ?ov�A`>l4M�R��=��^><�}> �+=��ս��3�뫾�.�=��>z?�e?�h�>}�˾)�c��	���?Ź�>�!?Fa�>�$|�
���0%�V����W�>y���n�������o5�(p�㥣�]�?�?��=[>
ӏ?��7?9J?p�R�C�'���l�� ̾�3r=�+����?!#�>� �<�m���8�)xW�Fu9�q*�q�\��lT��(!=� >u��E�>�3=�鋽j���6b��D�P�{��=3�i>鏼>��?��">�'�=�����ھ�sB?�Ѿ�H�_�*�@��}c=&>O�C>�;.��-?8tr���}��u��$��z�?���?&g�?Y�8?��ü���=��S���ѽ���=�>��#>�~B��I>���>��=J�M��Ӿ��>���>��>���wt�����ƽfdÿM�[���+�=��SE��6J�.(�rzs�s����n�>٨J�� ��و�qF�a�BbK��&��4�vʹ�� �?�0?��=��>�H����վ�p��e
= �C��l�<ο2�!L��+ǽԏ�qO��4��ƻ�0�'�̾�d�>P�޾⁙�_�y����Z/>S�a�>�@?[?�[lL���6���x���>(�>GA=!~�}[����=��R?n�#?�����㾟`P>��>�H�>��>�Ig>���x	��"�=�:L?
��?�ym="��� g��'�%3�?V��? S?SX����H��*�6�=�� ?�/?*��>�)>Q�=�<@�A|(?!~?�_1?8*3�VᆿQMľ�
?}8?'��U��>=��>Ǵ>.?� r۽)il>z�2�sU<tsȽ_6>!R����u�=Ѻ�=�* ?��x>:�.��c���>=��5.��E��r�>�;��>�#�>�C����u>��6>��#=A�6�'!���k�� ��|gJ? ��?��C?c�F?�A��2��'����3>�)�>3��>��>}[ս+��>�>����k�u���᾿@?���?e��?!cF?b[�O*տ�x����i�3+���.><��=�>����w>Ж�=�ҽ�eͼ�*d=a�>0j.>+]�>A�>�R>Po>�����%�������y�5F��'-����ՔӾvP
�E�%�q�+����������a��3�'�=Qy�� �%������]����>��>��a>=M�>b�=&E>d&����׾}C~�<�}���߾�㾫7�ܙҾ�S���ǽ�g������<�f���?��u<��r=x��>��<e��<�$0>�$�=��">G'>+P>H(/>j� >��>�8�=OK>d�=�^�>H��="����}����.�#{����=�7??@c"��������SVپ�Z˾,�>�?YEL>�#��Λ�Mc��F�>�;�u����9=�Z]='�>ʲ�>�5W=�x�=�����u���½0>|:�>���>dd���Q��ɲT��H���>\�̾���=�>+�$?lIs?"�2?�٪=��>��o>�I�>�C�=^XJ>^-D>�>��?��3?��2?��>���=]��B=!A=|yN��`�vC���3��(A���<�X��v=��F=���6]=��==$�ʻ�	�<� =��?��> ?.�,?oMv<���KC��T��َ�2�M>��G>l>*>5�@?�?Sl�>m��>�Y��{P��m��l�>m\>.&6���9�^Ym>Ol�=i��>,q�?�x?��@>���m���-q�=+'�>ה?�3?���:�ғ=��>��a ��z����4޾��2��\z����=�b����`��7>�
8���w�a��<-��e�v�Z�>�޴�I�#=��I>�l�>�G`>	�&��?��U�A��
&��:X>/�$>(妽r��=i��=e��r�=�$�<V�>�OvT���-�g*t=:#�=?��'?Ə<$]^=�������iW��1!?���>WE�>��?!_�=�}a��iT�|����>&
S?L�>P��J��=~)*��f��Xx�>���>�jj=�(�=�u�o�$�BPR>9?�f�>}��>нbia�QP��~�>���>��<�;4���?�c^?������}w	�m�U����͆�=D�Ah�Gy��ts�8�<���׾~쾷�h����=�a�>)S�?��W�p+�=�F��\㕿�v��[��{�=�'�=���>�u�=i�j�ط������f���'�[:�<��>�����@#?�I?�%�>}��?�?��=pt>�>?S���:SN?K��>�*�=��>�Y��0`��H�Lo��l��e ����f=˱�;��>�F�=^>xsL��7=��#=�N.=<�|�<��{�<�l#=P�<��>k�>0�>��?;�?1���c�x>a������}��=�0���;<������:r>!ח>��G?�N�>��>����ľB#����=5�?��?�8��󩽬Y
��ܾ�/Q�.s�>��=�i����f��($���{�=�@�>���>�Y)=�h0>�^�?��D?��
?m��������s��p�=R=�� �>R�>I�����&���l���V���7�&i����L��ך<��
>8�=��>(��=b�>U�<���_#��x�<�����>=��>'?��>Z	:�����ᾇb-?\���r���]ξ�n;�W��ܝ>���=�E^��L$?������1���T�(�7��>`5�?yY�?m?����U ?>�x�=i�ǽ���;L�<[T=Fz>�i>S��>z]v=�hn�٧��=\J�>70�>��X�����G<�.;�I���0]����ge���^��m!����^��@�P��?�=��afo��4��)�W��j�
�Ҽ��='d��:���?�\?��%>ld�=��1�`.��þV���Z�
K[<����*T��3�������⚾�S�����H(�������>��ʾ;q��1�l�0�׾Ri�<F�>�X?��q���-�!�Y��>I��>s�?�	��2s��z�ǽ�[?p�=?�q$����S��=˿9>�K ?��=��>>�5�=��-a�ʇy?�ĉ?��H�%̒�R㪿d����¸?�ʤ?�uQ?zZھz�i�@'�1���PJ?h�U>�u�>�;_�rT?���}\V?G`k?�	?3�)�喐�iJ[; ~>�C7>�xi���?��?>�t>�Y~�#�7+����]����ة��P���}=�W��|���>�Ё>�>����+	�=�>lW��nT��0�֩�SF^����>���>p�1F�>���=P�=E�.�!��O���e�=4L?�[�?�(?��f?��������ݾN�<>k��>���>X�>�O{�H3�>�O�>��ϾxD���۾�{�>$��?6�?��^?��Q�aSӿ����v��~�����=ˠ�= k>>ȱ޽�ۮ=�rK=�7��no@�)x>K�>Y�n>�)x>�3T>�D<>u�.>����#�,ˤ�uϒ�ÄB���u��)�g�~�	��Px�s��h�����������󶽍�����G����3D=��G��.�>�۟>P �>�+�=�$<R�>M	�=�l��K���?x�
�о�˧������m���#O��[���P����O#�o����'?���]�l>0�r>����3�o��˷>�,;��e=��x>�=8�.�B>U>ט->@J4>`m{>�E��>��=��x��>u�6pR�t	����>��V?�y��������lc��9���n>���>��>�_�AҚ�������>��.����&w��k=���>�>�>۞c>�l?�|fQ��^D�$+���m=fz>�{>?�=�,����_���޽�:�>M�վ'�=��n>M�'?�su?�S4?h�=޹�>j�d>�p�>���=M>�lR><��>�?�<8?�b0?���>��=��c�%�8=~|*=�~C�+X�t���"?�?�*��*3<9��E�j=,�v=;Qv<�_b=��O=1�ؼ�<���<��?�5�>�ե>ЍH>| ��q�Q��{l�n�߾�q~��'�=	�>��"?қ1?�;8?���>1�����to���gɾ�r�>v�^=�v����̂J���~>��>AqF?���>������<��C:>��>���>�$?!�>�J>vuD��	��Ͽm��U��CR�%x��	&��<S'��"�U����6%�����8�<"�J>��v>P�c>[�5>r�>��+>v��>�00>�xc=t/�=G
< Կ���`���m=�������KU�*V��ԗ�&���1&��`c&�-nI����a��W�?u?�S=#�<����3$�E!�����>�'�>��>�x�>��I=!L���N���P���¾n��>�>?�?q�P�=�+��t�D2�<\��>ۚ>V>�Q4�������>,��>�?�6�>����>?���j��J����>2�2=ڧ�H�?�Mk?���B�þ�1���F��z�PJ�=s�6�8�x����C�#�B{"�N}̾C�����=���0>X/�>��?�o�����A�i��	��%�q�� '�h/>��<�т>���=��Ƚ���#4$�|��g����^F>3Y�>����?oo?:\?���?�['?�7�>bGS>���?1/�;+?��Z?�~h>v�i�;��>�ib>y�?�qྲྀP�����9ĭ��Kl=kb�=h>Al>�=�=໒���=�>jl=8���k#;=K��W=q�=fS'�4C�<��>/X?���>��������Bo�#�	���Q<fe�<��&��8���������H�=!)�>0��>q��>�I>[3��p�~��W/��g�>��?Ϡ9?h�?�� �sF��C�.�׽>�6>z-�>]c�<NM �Q1�[���rWv���>C:>L� >M�R>�?��A?7X?<_�Ӊ-�׿p��[ �Ug���3��>�E�>Ѝ_=Ǜᾌ�7��3o�9,[�!+�=����NN�U�<\��=�Z>FA>�ž=�8>�#=�ř�ȽϽLҺ�{.�Xʪ>���>2<?"K>��=櫨�"X��1]?��O�5�y<��d���P>�ʖ>Z�%=aKV��v6?�	D�_|���M������l?(��?�V�?��9?�<3��h�=K�1�?�L>x�3>���>#S<MݾK(ξ�[�>k�F�c���s���ޑ>��*?D'@?d<��E=+�e��Q��<��¿�<H�&Hu�pAF�+�a���������+�VV��λ5�C�\���K���p��q%��m�A�����ξ����?\�$?Pf`�����.N�ک�
PV��$�����>א��_�)�1�&��e��P�?���žE� �\���Z���H�>��������E	_�Dt��r\�=>=H��>Ç��e�,��d7� e^���}>ċ�>�d���n��͕�ˤ<�(n?�"?4�þr�Ǿ$��<���=m��>�O�>.^�>�P�c��c�$<12Q?�6z?��<r6���V��Ae뽈�?Հ�?�cN?����R���������>Ͻ�>���=B-���<�jվ5>Di?�b-?�-Ž�=W���-���$?�)m?苖�}��>z��>�SB=P��R}]��^�=��x=P͂��->��j��o
���T�������Z:���>;h/>J�Ӿ;�����>1��CO��gH�����C�ۖ}<%�?
���_g�=1Hi>۠>�y(���E�����L?��?��S?m7?s������u��V�=�}�> B�>Rӱ=�
�>�?�>����r����g?�i�?5��? Z?��l�Jaӿc��	,��w��UF4>��E<ͷ=�^��ݽI�3�]��=���=3X�=�c�>H�E>�s>��=Y>Zs[>8(��H�*�3+���X��������KT!���3�C�.���:��������ž��ܽm"T��ý�4����+�o�]='{��M�>�?�y�>{6�>)�.>{�>�	���
�R�e���N��ߘ�A4ﾕ�ξ������+��Vi�rW���Z��߀�m?�t=rC>9��>�"���=�׌>��=<*�=0�9>Ru>��?>��>��X>�(3>?�0>���=l#�>�Ol>C
���*��#�<�@�>5ؾ[�M?������>ԙ��D'8��ܾAʋ=L`�>?��=�v(�í��V}�!�?��>�5������ɑ����>�b�>��>�~���)�����1��<�������=�Z��X3�Y���:/=��>V�ܾK8�>:�?aV-?��o?�y?x9>4d�='>�h�>r��C>�Բ>��?�{X?�h?��o?MG�>��>�e��B����I>M6�B*��'�����<0\�h���b����]<$�)9�����#>d`i>��ż���=\�=1/�>?�E?�&?�v?,^� �^�*y���2�!Y=s[c=J�?���>�B�>R�>���>7�C>�I>�9�����`.�>i"e>xM�R�`��>��>��>�&]?|�>p�=]E�:C� �p=���>�4�>��?���>H�`>2��<����8kǿ��W��� ���-������T�Z��=�ʈ�1E���b�^��D�>!;�>�h�>J?u>�>\�o>."�>[U�>=�>.<REQ��`< I��iW=�86>��>�_�9�ǽ\n=u"�=���;)@X����jȽT�	���	?>�?��G�Xn���m��� ���V��=t�>y�>Ԝ�>Ē�>��>�� �+�Z���J����]�>~^?��?1?5��s=UN�<�~�<���>{��>�>�ᬽ�M��u���#W<.�>l�?丵>�1��$R�.^Z� ���g*�>�4$>���q�?�`j?��S�L�˾0��ӆ{�.f����Ԗ佫!�	�o���-��p��D�N��Ͼ3>,j�>���?�K��{no>�b��ᚿ]����D;�PJ=p��=�
?��>�t���Q�wS�+�S�����!)�9���dc>.��>��@?)'&?V�(?'��>�'?��;=��> =h=N�(?�a>�R�>>�
?i�?�k�>#�?�ڜ>b�K����s7���px�Ho\�iY>X<M>i�>K�=���=����T��h���v����<��q�=c��>)x>��=_�
?l%?J�}��Ұ��/D�W��6&�<��=lX>��2�ڬD�"L�;�q>�3�>��+?6�>��=��վL ��� �F.�==�?E.-?�n�>�w�<Z�=�[ܾ�q��p�=�_]>�=0�l��I�El��\��䩓>6l�>T��=�Z�>��w?=�?]O�>�C$���P�|b�eDJ�eN�>��V� �?g!�>�"2>Q���q�Y�u�u�k�~����2��뇾�/5�z�;>��><^�=�k`>��x>vS�=���=�h�������]�>��?�?F�a>˨�>��$�xȾ�`J?ԕ�����j�����Ǿ($�{q>�H>D����~ ?�z��C�P/���f;�L�>�?��?!i?+�7�l.���_>d�T>=�>Tk�;��M���_��^��V6>���=0t�к��-�t��M>��w>Wȷ�4��Q߾�oB�q����N���R�k|ԾB�}��>��� ���@ý�s�A��=����B��H��;*��@;�Au���k�]Ǿ]�Ⱦ���?�as?�9/<d`
�������%��r,(>G&Ծ���<�þ���=s�f�r�׾�ݾk۾�<�;�1�
?P�=�̑� ��9ྷ�>|ф>:cd?��D��mX�?Y�>���=o���v�s��Ӎ���۾#>x?��?S[���D��>�c�=��I;I��>u\�=
}��s�l�u?��]?;?�>��(_��,:������c�?t��?��=?�/t�8 �q� �����O�>k?��>]��� 뾴<���7?��]?�*&�gH�儗��1G���>���?�T��7��= �>���>ߧ�v��zT��Z�	�=-�=��=�w�>Ңƾ��x��׹=ֶ�>,I�>*g�Ċ����>�n��XL��kF��p��="�{Ĕ<S��>y���S�	>y�k>d�>�)�x�����������I?y��?��T?��8?�! ����Pٍ���R=;D�>��>+˥=�?��q�>`/�>=L�F�k�U��A�?�_�?� �?�W?'l��0ҿ[��_�^ʡ��0�=�u^=�>�*)�f��=G�<|�C��涽@�1>���>��w>YX�>�Le>�,�>7�=(݆��(�J��3���� C�Ǚ�ܪ��̼�+����������WvӾ�t��m#��2��@�ɀ��R��l#���fS>'u�>��>W>G=�i"��yU>�Qо����Ѿ}A��(��5���B�l�R�%�c����-�G7�=��!���4�B�?��>ǉ�'�>1��<&���]	�>��>��½���>�v>���>��E>K��>�(�>�'>W��=1�_>B#>kV���-��b�ʾp�B>
K���4�?�X־��;>�i��YM�������'��� ?���>(e(���������?P>j�m�b햾�t��wa�>��?SO^>�c��I潾 ���o7����o�=�BO=�=FZ���̾w'�=��>+�����X=�Q�>��B?��k?}�=?!n�=��?�:�>�N�>���=��>�5�>���>!e�>�zF?��1?�9�>C��=Os���/7���
= 	���v��l�e�����n�>�V��x��=��=�?>t(�=Z�X>�`ؽK�a�'��;ZL�>�99?v2?%��>���b�K��3��ɽٳ&>��G;u��>�?�->?�S ?���>�r>c]�<���vw�_2}>b?>W^?�x�R��=eY�>�3�>��b?&@1?���=�ѕ���P��c�=+V�=)�?��>��7?�e�>F	=�����进�0����1$��c�=�o����u�� �߇`=<�������CsF�Ο�>G��>S,M>�/�>���>�_�>E��>}�#>
��� �<��A> ��=��ֽx��>N7j��"3=�(˾0`�=)�Ƚ#8�<�? ����:�/�3��. =b�?��?zߞ���w�ۓW��B���+���N�>&�>,��>\&�>�@�=��*uR��;���C����>��h?W2?�:6�S��=�w��hv<�@�>��>_>~:��ٜ���E����=?�>u{?Y$�>�]�b�Y�Y>l���
�8{�>+'�=��n��?��e?�;��*ž���B��b`����ȍ����ꐮ�I��PFV�zw׾`7�s�^���|>_�>=A�?��F�|�=G]3����MΞ�����3�=,xJ����>,F�>��k�;����h!��W����о�f-�i|�=?�>��N>r��>O'?d�E?���>�}$?3�@���E?� >k�>?��>��?��?	?c�>^(?���>.�ý1��J�<�hN�;ȓR���>�>�I�=f|Z=�Q`=f���22�<�^�o�B���6�N�3�0��H��<ud;>�>R?x$?�C��߼ufk��3����<de>c�^>7z�hOR��\�<Nd�>�?B�/?�B�>���=>վx������l�==�?!M+?h�>��=���=֢��@�w��=S6>�y��cq��|��%�������k�>���>�>:�>�f?�>;?b��>UR�>n��*��7�F�<}���&��>qF>hEQ���Py��L�$Kz�̽9��Y�_^��G=>�Z>�>�W?>�R�=���=s�C>PW�=��O�6>�s���>%�?�:?���>-
�>R�I���(�}�I?B����q����YоУ�N>=>���?�1�h�}�:���J=����>���?5��?�5d? D���Y�\>�:V>�>��,<��>�9���N��)�3>���=��y����1�;-�\>�-y>$ɽ��ʾ?�1�H�e�ĿX|�5d��}��Xց��Y��	�_T+=VY�� ��=��@�-�[�����8�}<�5=ASc���C�G�žy�ؾ��?e �?�<j��X. �Z�z�@y>W`�� 0>�E�����=Az`��s�����Ž7�T A���&���>p�Z=���s��N�>���>ZB�>H�A?��	��jξ�F0�Y�ͽ��c���������� !��qƾ�LX?E$?�*��V�	��>ܰ�<�4�=�[�>/�t�1���5@���?�m�>�Fq?�7��S��r������ͺ?�d�?&O@?s���9��@��G^���>-�?*5�>CWǾ�侱Q�ܐ�>w�7?�W>��%������/�"��>��q?ၾH>s�?�><� ��̹��PڽE1���ϐ�M�>��&>��O�;6��:^j���6=*c�>��c>OPS�h�����>�2���N�v�H�/��������<�x?���q>Qi>->{�(�N��fԉ�$_���L?Ǔ�?V�S?�b8?Sg��%��l;���'�=��>P��>�^�=��ў>���>�g��qr��W�?�G�?g��?xJZ?s�m��ԿS㠿�;ž}���v�=��<笩=5'��4������F�y��t�=�	�>#�>私>sr�>dul>�X>F��+�*��Q����vh;�>j'�xu&��i���{�@{�������š��oݚ<��;H��5D�5��R<�`$��A��>oP?�E�>��5>��=v�>1
ʾpE��a��z�]� ��/��<+��Q(�K���d]���Ͻw�E<��2���>�IU>n���ŕ�>v+>"g�yt�>G��<i(>Y�z>*m>��q>|�A>Xj>��A>'I�>
H>)7�>�ĭ>�5���}��Eel�-~�>G,ؾ�JZ?�Z���#>���	�4�ӾO�e�a��>h�<��?��G�������>�R>�h�p�h��蔾/B>���>���>�+@��D�������½������F=Ā=�>*��p羖5���M���?�>��վ9O�=E��>%�?e�1?"�h?���>{�|>�_�<Lr?ڄ�=Už>�?"�>O��>��O?In?`��>N�=n��e�`�"���>h:��Js��V���c<�<g��1n��Α�cJ�nq!����=��>�)!<�z=�=̢�>z�6?3�1?$Q�>&���|T��y�+޽��="�>��?��=��M?�1�>-�!?g!*?{	>T���^-����>�>{~g��hs��7��4��>{/�>C?O|?,��ñ޽\0x���=׍?��?�j�>e?�:�>�Ͻ���߿XF����+���A���S�D�о�����+>�y̽���6g�=���>�l�>8B�>�4l>�V�>X}�>�Y ?ǁ>�v��q�z�$�d=�t�=o<ڽ7��>���=
%>ܿ^�_��=T�=�'�\K�|W��>�<	-�զ��˒?T�?U*��K��-̓�K�ܾS���O�>
��>�{�>6��>A�m=SM���wC��@5�{A�n�?݅k?���>E�?���=Q�켼:�9��>Mĥ>�*2>MQ� �ʽ������;<SV�>��?
i�>5��v`��n�V�	�pƱ>Y,#>Q�Tڔ?F�k?3gP�G��D�������m�
���ia������L�*�L�O��F{��̓��'>2�?�P�?ޞ
�9>�m�/�RL��ѵ��
�]����=/���C�>�>f��*�I��p޾(�Ǿ�����tؽS	B�(�&>��=`ܺ>=�$?�U?�
�>ٹ1?ݣ�<���>ȯL���?sJ�>me ?U�%?�~?-��>��?��>*�=�r�Z��o�=]����	�=�HD>�5>�@�<Me�����=K½�[o��_=H�=���;��ȽVР;e��=��7>ld?h<?�<!=�-�T����D���3>�'>5��>)��=��m�\��g��>��)? �%?��>�|5>g�m�+��d(��SU���t-?j�S?Ew?��ٽ�z->og��;�����>�+1>͞<�0���c��'������Yt=�~>䚲=:�>�*W?��\?��?��ԾWl��x����F� �>��ܾ8��>�j?'�c�,��7U�W�b�H�X�(&7�+^�W�������Q+�>O��>�=;7
>�,i>e�=������>�`>]�+�_F?��>�6+?SV?���>�Ը�����1�I?�ˠ�>�5���� Ѿ�����>s<>_����?(�Ӽ}�vɥ�q�<����>�j�?I��?�Td?D�]"�vQ]>	�U>)�>�t9<��<����f݄�+�5>���=�y�PZ��˪�;�X^>�w>Ƞ̽�tʾ@�㾣PB�yT���4J�*־��F�>V�`�i��X>�,���6>�$� }��Q��;���V������n64�}���]N���T�?�u�?J�>ԙB�<����S��6�ξS�=O]���h:�x�ƾ���=.�޽���辄�ܾ�.�Q�7��b�n�>[��<uR�����nk�"�=�2a>�V?H���!�� B�bve>x(� ?X�e��:ً�����(�����V?y^?n�ƾ��x�E��>Pݎ=`m0>IQ�>?�;�����k���
&?�{?�vI?=������E���+��U_�?(��?�C?A���թ5�C}	��N)�,��>�^?�R�>D>Ҿ��ӾR4�(�>?P?P(>��7�S�����;���>!ly?����p8>5?[��>/�V�E1Ǿ�ҽ��ݾ����&>��C>t����I�ؐf��`<)��>v�>26�����Q�>*ҾV)B���3��������1+�=�k�>����4<q=ںY>��>�H�K������?�b�ĺ'?3Z�?��_??�?���I�¾ �@<�A���>�ӟ>b�%=��w��>k��>1H��_�a�پ�d
?r��?{��??v6?�+q��Fӿ�
������������=�/�=?�>>b�޽^­=ƔK=���B=�݊>��>Zo>�8x>��T> �<>��.>ݤ����#��ʤ�ْ��[B�p �����vg��{	��y�ӡ�zȴ���효�E���9ؓ�i�G�x��zP>���߾�Ud�{M�>��h>p��>��>�%�{�
�'R�p��7ݭ�;$���	�p{ʾtݭ��G����)�.k|�&� ��=��K��>�d`=����r?�M	>�>�=l>J�K��|�=xA�>���>�W�>�@>Y��>�̦>l��=i��;�+�>o��=�|�Z����dǾ��>q��W1b?�z����y�Ja��d���꾟'�=��?�V�>jO)�M����u��?��`>z6��v�������c��>�{�>ڢ�>CUI�G������������<vO�=�e�=�����d�>�p��=2�>n۾/��=��n>��)?FDu?�4?܄�=a�>�.>su>���=8`>�n>l��>P�?�>?�Z3?Ҁ�>�H�=�
���8G="�F=J�9�u���h˽_fK�k������V���ђ=_�=�#��a��=U�<�ƕ�CY(�>��<���>�I?<�?&��>c��a@H��:=��.��p�.>Ȗ��mR?\�>z"?�7?���>�E�>�+	>����ʷ �deI>��*>�gI�|�^����Dǟ>�L�>5Ue?�� ?h�ӽ�󘾛h����=PDe>�R?�	?׊?L�>�?+�c�&���g��X��!��׻�;��/=Y`<�Vos�7��ދ��p�<>�|>&�>;�J>�Q>g�=���=�.�>�>�2�=��<�5B>cg?������$�=qH+�^�Q>�ԟ�3�p�&-սb���xF��T��?lN=�C����t��>d�?tR	���׼FФ�T�$�y���/{�>2�>�t�>8�?e̅��a���_�-�h�	�$�>�q?�7?/(Ѿ.��=�l��%�;�}>U|�>��i>?(ּd��·ɾ-	�=E2�>��?A��>I��=) �Y!��D��43T>u�>��K�u�?H}x?�6L����h��I:`���N�yb���4�����&��x�#��7��	1�qS��{X�Z�>���>Z��?kx��UՆ<��U��8���l���P-�oٛ>�#>�?���>t� ���罩����;P៾Q1Ƚ��'S�=�D?�R?�m8?�g?�A�>��*?>� ���8?Al>�&?�o�>�L�>��?��=?6�
?��2?���>�#~���d��e��2V�=��<� (>�� >^>9��=}�<b�=K�=낽=�.o�����N�=��=,�F����=���= �?#?y쬼���<�����@�+�=�,�=�">]�_��f=��ח>H�?��8?K�>]>GBƾRU��ro�r.�=4��>ɰ1?�g?F:�4�.>G���%.u�%��<y�%>D��:�t���5�=i�@���;��>��[>D�=�0�>��l?T�D?��?z��bH�wГ�L~�I[{>��4<�?p{�>够;. ����<���N��<��D��lN�xX���@}=ku
>�oS;�S!>*,>|�>�u=�t����'>�hv=0+e��y?��%?�K?z�[=YF�>�k�0�ݾ��I?�����h��ᠾ�}оE�g�>)�<>`���?����}����F=���>c��?���?�;d?��C����\>�rV>�>E�,<\�>��3�6Ʌ���3>q�=ňy����~��;z]>Dy>Pɽ��ʾ�<�s�H����@n�X&f�-�z�O>��m0�8I�<�쾱A�=���q־[�������M+�7a���]���ج�����?�F�?&��Q{�����,Ͼ�A���>��>9�K�=m[�io��*�����,/�5���^I��3�U���G?��нH۫�4섿'���፹>��3>�Dq?ٙ�������B�P&~>l�]>��P�0��������띿����o?Q�/?Z�!�K�����>T��>��>��>[ᄼ�Z3�����R%(>�q?}�M?C}��H�������96��E�?���?V�W?�k=�K�C���۽*\�>J�?��>pU������Y���I?G~=?Һ��̗>��5���WQ�y� ?��?�5�/>�zA?;9�>�D��!)$�
�/��e �?W>5�">#���D�������+�~��>�w�>� T��ݾ��>'ؾ0f?�!�>��u�tp�z�=:�?,�!�ܰ0>O>P�=��"�Ja��hڕ�vG��I�&?
q�?6gm?(�?����W&��ٔ@=���<vz�>s�u>��=�����R>9R?���Ka�l�о�?,��?��?��A?L�t�8�ٿ�����:�������4=�V���l^>�j�=+��=���O��Rܣ=asB>-�6>Fsc>2�> Q�>��U>M��>q��;���Y���ƕ��RC�W��T��Q{������퍾��Z����A��R�μ�"�K�>=ë��W$�$�&=-�[��&T>�c>���=g�>���>fv?=2wE��Ӿ�;�_�k��@���Ҧ�&)�%U¾�D����\��z��mz=v��(Ϥ>�70>n�T>|��>��X��,<�*�1>�
p>��:'��=�8>/�>0)(>Tf�>4[��f�>���=��>@�><�z��I����z<���>t����99?�Y5�ĩ�>���=80�_�yAH>a��>H�=wM.�܊��H����?� >f����R�0!k��9>a��>Nǋ>�"����+
ɽ�I><Ba��$J=d�b>6�=$��#	��U4�=5�>�ȾD��=�(�>���>�	#?a�D?#=>�f?&jz��	�>
=�P�<
ڄ=G�?�)?8�i?�ji?5�>���=j�����ؽR-��y�'�Iݵ�U�<]Ƚ�V=+�=[Z���i�'�>�o��@mf='	=��K=d����|=|��>8A:?g,?�?cr��;����I8��"x>N�5����>y`?���>�?�(?���>�w�|2��O|�W��>I4K>��F��[�D%4>��><$�>J�S?p?������j�<���=她=���>�}+?c�/?�/>�Qq�}>
��
Ύm4��+��A�,<o�4�`f�S�޽��.�x����o�_|��M�=��V=��>��>�^�>�ȑ>���>�>BI>��A>��=	p�=c�^=	H���W#=�&;+z�<�p���Y��n5����2=}ؑ����e�Ƚ�m �0%Q���>6x?�<���L~�s����3=���>�g�>�^�>���>�Y=4����M��I�<����>~�U?"�?��+�ԣ�<�p��m9X<g�F>^~�>?�5>.�s�x���2G��+�=!�>��?ꂰ>��2��G��co�ESԾh��>�>�.;��?��u?@���Ӿ���-oq��ྒ���
=u��������[�b�q����
�ƉԾI�U>��>:��?�<�?>;�W��B��բ��$I�\7>��u�l��>�0?d��XB����5Nƾ�z4��L�s���C>�32>�vC?"�:? l6?��>D0?�&޽pd/?T�>��?�Q�>%�	?�?e/%?��>��?�@�> +��b��b��̝'��.�T.>�q�=�3
>XJ�=ڐ�ϕ�7�ݳ��-0�� �� =Y �)$7�k�=�>|>�>k�?��%?�=��<Ȟ	�ϩq�J�<=Y=�<	#)>rf	�o�ǽόW=s��>`?+.3?��>� �̽׾�w��?��S�L=�[?5�.?�@�>�"�<29>�̾� E��!=7g>RG������yj�d�����vZc>��>#�>EE�>Ps?��G?��#?����l�g���~��N�*L��%/{���?�?�k�>�����GS�W�U�!sU�Nl1���л���S��=��8>�h�=#�>"n�>�ؠ>��x>-��=��
�C�P>1�B����>��?VMb?��>��\>R����3���I?h����	8��i�о���T>CW=>D��?j�
���}�����+=�Ƙ�>{�?��?�#d?�[D�P��]>uV>}�>�A-<>����G��s�4>�Y�=��x�!ٕ�Sx�;y~[>}�y>6-ǽ�`ʾ`_�}1C�2�����G��{��l��m����3RվxY�<�[4�W�K�b�"�徾��+�I�O��Ƈ��z�0������[-�?���?P�=#6վi���W�����x>��=�ҾZ����#����Y\����ۗ���\�$��OO?��)=㊞�͞��/>��o���Ơ>�4?H�R�Q�>�2W����=Aۧ����� g���K������_?|�?}
�ˆ׽�ñ>���;������>�k�����VJ�<Q�>NC�>��Q??�վ�8��a����{ε?e��?�.8?{m6��@���4�?EL�>���>c줾q�n��ZR��9�>��#?�>ͤ�`��	M$���>�?I?d��I�Q>2�>Ѩ>h	\�\���|����s�gP�;��=�ʹ���ɽ�?R�����2�=���>;Hw>4����׾�"�>�����TI�ƕ4�����V�D������?����a�P�`>�� >4�����q��ـ��k??漥?��?C_N?G��G�"��'�x�]����>�^�>��=E���N	>W(�>�"Ͼ�JX�S����>�g�?�@�?[�?�qn�� ٿH������f�̾�L=F��=V^_>F ��R	>���=��B�LԼ��?��	�>>YD>}�d>��=�@�=j���K#������▿�x3�������4u�MN�lJ�����>�Ҿhؾ0.��V@�&SνY���%L��w���u���*�-�r>���>��>#'���s>E�`>6�
��*�	B=��� ����c�������ǵ��!������=���!��>H1��D�=���>�����\H�E_�>��A�WI���;]>ռ='�>�>l�|>�>>ƋK>����	�>gr��s��m�����L>8�=_�@?��߾o�3�k���T;����x���>�%�>�������%⡿�@?��B�ٺ⾎��0>>V��>H+�>�#�=(ϻ��>
4Y���Ѿ�
=w�?��>p��!�ޛ��,Q_>l��>~J,���=>��9>�V?�74?k�6?���?l��>�_���=]�=Op7>�4�>�,?sjR?8�?y�>�zj=}Ƥ��P6=l�V>�߬��O���_�=��=�"������K�5�_:���=
<�4,J>��#>�M=؄������P�>U!T?a�?�ac>��#�6ἾEu�y�˾KQ>��=@�>��>��8?��>�(�>�Cf>k�=cv]�zB��1��>��>p@�켃�Yؾ�&z�>ǋؽ��Z?�?C>��=WO���o�=cd>�j=x:?Ĺ?>���<���	̿- �k|1����P���-�<���=ĝ�R0��._d�T\8��㽋/;>CRG>��=�@�=|n�=6;�=���>��>K >:1.>y쟼�o�e��G�=�.%��Z�<R��=����Q�=�+v�����]���	���=g�b<��?g!5?��$�卍�lܾ��˾~޾�,K>���>�I?�/?|�P>�m��s�(�0�u�W����>0we?��:?�&��1*�>z<Z��	0=��>���>��>��=ow=�������[b>���>�y�>r�x=�F��i�F��N)>���=���XG�?�L?�\7���i���
���O�C��Z��;">���YV��6������W��Q����J�۾f�5>��>Hɴ?奔�?\�>����?g���p�
�	�M9���I=z��>���=�8�#�7�����S���4��n�Fe�=S��>�-H?-�H?�?g?�=>�?���K1)?�a�>&/���?�>t�?+�?���>��>� J<�}�="��DxT��ʽъ+��>
b=���q���n>m6/=���I���F��ڰ^>y���\���M�]=F3>���=��>$ 1?$�<>61�>G��=�G=�����1/��`�>I��==�����=�t%?�g�>R|]?��>D�>=f���T�����Д��'?.� ?P�>�]��b��>�Y׾�Z�;�*>�\J>GS�>��0������&��9i�9v�=D�H>B�+>T�e>�M~?(?�*)?������_r���H�?�R��+0��iS>���=ܓU��/����_��O���h�-C�>::�SgZ>�@#>Ug��*�>�h?>�bi���.>e�,�d�E���-��3Ľ�S2?,��>\>!?�>�����dj����(�I?����X��VE��1�Ͼ�6 �W�>P::>�o��m?�s���|������=��4�> b�?��?]�c?��B�F)�D}Z>�U>q>�$<[�=���������1>�:�=c;y����s��;0b[>R�{>��Ž��ʾ(��~J�Q-��\�T��%���k��]���,D�[�b�Q�>�����w����c���7��t2��E6m�7�������Ұ��������?d�Q?̧0�%B�=�!&��W�+��o�[>u˾�:��������
�ۈ��Ntžn����b ��侷t
�Ge�>�Oݾ�̦���������A��>6y>�U?� ��k�}	���爼*NI>�ŝ>R��%�m�U?�����;FB?|2#?����1��[����d���>Ȃ�>S6>��=�u^���>�(�?��%?�A>C���F���^������?_P�?�BN?o�����T�0x�#پj�>ƽ?0#?Q�	����>%?vI?z
�>��&������eH���+?}�?*!��:��>��?Fg�>i�}�d��$�½�����נ�h��>�8�>����4��L��JPr�UyV>6��>��۾���Ӝ�>��2�H�3p&���0W2��u>�\?��`!��5��>q
>J1�k���N���8����5?Q1�?��?q/O?g��x��]RJ����=���>���>#���_�yQo>�ݱ>E�㾈r�A��f�?q+�?���?�.$?�Q~�����'�����Z���N>:�
>���>�����s�=��>�}���n@��_<���>Lӊ>�>61k>�_>r�.>XM���(�3"��4����9����A�k����og�4
��D�����舽5����*�������q����Ì�2�{>,��>�(	:��
>��>"�>����f��鑽����� ���ɾ�Ո�g����о��i�0������<��`D@?��Y��>r����>o2��i�=��>��M=���=�K�>�*+>^�O>��Y>r�>O`�=��>v��v�>����f���/On�XLB��q>��_>SU?H��1����*�F�'E	�PI�>{8 ?9>ND!�m׉��*��f�
?�2�����!¾��=���>KAi>��=b?�=L(�=%��iT
��H>��>�J�>y����p߾�q��w�<��>������=�9]>��?3�q?�|&?M0�=��>��>Ҏ^>�1>n�j>�a�=Ϊ�>��?�;?�4?x7�>o��=�t���=O&�=��6<��?G<����k����zO�٤<��ű�&}�=dЂ����=��>���*ZH<�;��0�?6�G?F �>*?���*�3����B�%�w>,��=8� ?�I>|?D�*>p�>��>Ϭ��o#ܾ(P�� l�>�7�<^-J��u9��O�=(�C>k��+Cd?�Kg?�Ÿ�zƦ�}Z>@�=L��=�>�	?`F??�*>=�{>����&ֿ���S�	�񨙽�%~�\.>��y�*=�L��>`����?�>���=�	g>��>�e=�>uR�>�xx>~ȴ=3�=�@A��Ea=�f���z=2\F����#�_9�-������X��=�н��H=���{��5�I�]�4?4�&?ٰ�����}���+S���ED�P�>vr)?��S?N�>1G�>w�� �S��E���`�o?-|^?G7?��D��>�=�=~<H�S>`�>_�?��)�񾞾���ܸk=A��>]�>�6>�>uiV�Ô@�1����>��=cd�Vw�?A�c?1�7��������4\���-�%�Zʥ�<	��Ѐ�y��;��0=ӾP�˾ �=X�>e	�?�����>������yi���ܾ��	<��T��>�ˇ=�پ�=��4���R
��	�'����+�=\�<�ײ>��/?c��>���?�LA�5h�>���O�)?�;�>�p2���4?�;ƻ�?r?���>���>��>u۱>cu˽��g���Լ	ؔ��	=d��=Nw�=��Z=�9��Q�=μ�=Z=��(��5�<ő=G���Ck�D�8�ޟ�=\�	?+7?��s��3e>}�=��P��k;��H=�x�>I�&������A�=	��>z�=N19?ǩ?Ci>B��=Yܾ���� �=[8#?�5%?�"?�=�")>���pS>��<�MԽIA���B����ž��=8�=���>9V=�(e>�4w?�~F?� �>�IԾ�t��<炿�?��ҽ �����_>ݢ鼊�*<
�'�����'�A�B�N�[�n�Y���l½�k	>`N>p˥<h'>;���y�	�=���{��=H�]>+�¼�9?<�>���>A��>����������kJ?����*\����G�о�)�~>)}=>�N���n?���={�)�`>���>� �?8��?�.d?��@����ҺZ>��T>�>�_<�W=����z��v3>lҺ=e�x�o�����;8�Y>�,>碌��|̾�@�БV����Y�X���5�A�[���ƾ�ھ�r˽��
>Kp��Z�B�|�콊ۼ��J��-��nu���*u���;�|[i�੧�T2�?�M?�j�=�j�=B�C����-��٥�>�B%�M������G��ʚ�.���b�¾>>��v�澾"��Q��wx?{k�n��d���2��ݴ>��c>k�?�4������!���O��R�>x�q=�����������Λƽb�@?��(?X_q�*p���>��o�<?y7>cD�>��>��T�����<"?:�?��b?�[��䏿���b�5�p��?ϔ�?@?�ch��m�ٯP�I�׾���>��?�`0?=y#�F\���1�>6
�>��?.�f��Xk��î� BF�M8M?�"q?Ծz8?�O�>�ǭ>s9�=x���#d�Њ�RE?=j�>F��<���7f��Vv���o=�8�>$ͧ>l
پu�����>0���^�
�Z� �ޗ,��->}�(?s�/�>"��>��=>R��◎�����}��0\?H]�?G�Y?��?Ċ���z¾DS�N��<�f\=��Z>�٥������?^(�>t��=�p�w�hg�>���?���?�*2?�r�Rӿ�������:���0�=&�=��?>��ݽ���=�_P=�ʻO�G�Q�>҃�>��o>x>�T>�\=>H->�V��T�#�$椿$5���A�y����� (g���	��v���������H���ަ��r���~����E��[�C�Ӛ��(�y>Ҟ�>�7>c+�>_�>c�>����菉����&����ؾ"��2��*>��X���͙�����oн&�影P/�Rs?$�>S�`�
?9��q>��J>��ڽy>>��=�P�=]�J>8��>S��>�i1>`�\>|�=,]g>;�/��F�m���<�Q���$�=�6?�WӾ����J�#�]�T�`>[��>�RF>��-����9ݚ��?�̽�o��=��Z�=�2�>���>d�P>�>uPͼ����G���i��=*�
?��>�� �F�ƾ:�(2>�߱>۱��2�%>.L>T ?��~?�+6?(�=O?�>�=>�>�_>	�>��D>�,|>�?��?��,?o��>u�=�~���f�=�)>����g=]���V �������Z!�z��P˸p4���2�<��=)��=$3;p����&�2`�>dN,?j�?B��>�8B�9� ���x��my=�Xk>��]?�>�> �?�#`>�H�>U��>vfӼ�%��Oξ��>��>�x��.l��CA=��&�kC��Xf*?jo?v����پ��B�>)���}H>@�P>�w?|v�>��>���=�s���ӿ���)�uN��bΑ�?��=��ֽ"y]�a>�=��J��#ҽ�Cj�&�>0��>�\b>��J>>m >@޼��?�f=`���X1>��<]Dg����7L�=����t�=��˺�h��v�I<%R����9=��`�	�|��<)��<�!%?v
?V����K��Fӡ�zL��3��/|>f��>�;?���>k�>�*ݾ�]�$v� Z��G?��9?��,?z6쾭��>����y�X��x�>bf�>e��>�����{=�|��e¾J/�>���>��>M�#>ǺW�H�j��;��YPy>�ʾ=w	6�R�}?�Ѓ?�T"�#��H=���h�^� �u��5��F!����!�E�ﾣ73��,$��;�4�̾4=��>���?o����m�>E��������k��4��i_<�f�=�`�>w�I=�,���0�-J���'�ef!<��P��k�=̗����>�|R?:�>)_?%>>MN�>y0Ͼ =?[�?��q�>B�>z��=��>`�.?x�>���>&��|�g>�6�䷗�@H>�ߠ�c���<>3<0>)|0;Hyg��U�=��W>|h� T���S���.���1��P���f�������>c�>?�$��N7�>B�>�a�>�<^K�;kI�>U�^�MR����>k|�>S��>��<?v9#?F½>+�[=z�\���/�V�=C��>E�?,�?�'���>�4��);[�#j�=��g�8ZG�^���NJ���S�(�G<�>K>|>�=�>��g?��Q?�+?>��.Yf��Ǌ�(rR���`�r��$Q?��L=Σm>�׾��־��r�C�5���H�8���F��諼O@}>�˫�,�\>��_>�FR�YS>΀���g��U��=�M��W�+?Rґ;�_�>(�?���Y�:�Ծv�J?�l��1��Ʃ�U�ھm��J�>R�T>+����?�}��0^{��롿�^B�I��>w��?���?�e?��2�����$z>�X>F�>��<p�U�1���B��f2>���=L!���ϟ��F���R>��o>�LȽ0�ξ)�㾣�[��	����o�-o9�<ͩ��������>�X�P;!	���%�;��������M�Md$����I�$����}Ħ�Tm��.�?T
O?�k�G���-���ھⳒ�,�=J}ɾڭ����C���}����#���[�\º����+���+��/?Gd �*7���v���)о.�}>�)�>�~?m�Ծ؏�N��(�"��ò>���>����0et�,�������10?|Q?*o�ps��*8;�%T-=�F�>�)�>c�>�qG������>_�?�S?t�ds�%͗��h�A��?W��?+NK?������T��W-����jj?�&-?b&?��ǾZ�뾐��=�&?��8?�>ho�EU��(���^*?a-j?r����X�>���>�X�>��|�Kӵ�~ߊ<�7����Q�&�>�b->�g|������������>��?��j�ˌ����>0���^�
�Z� �ޗ,��->}�(?s�/�>"��>��=>R��◎�����}��0\?H]�?G�Y?��?Ċ���z¾DS�N��<�f\=��Z>�٥������?^(�>t��=�p�w�hg�>���?���?�*2?�r�Rӿ�������:���0�=&�=��?>��ݽ���=�_P=�ʻO�G�Q�>҃�>��o>x>�T>�\=>H->�V��T�#�$椿$5���A�y����� (g���	��v���������H���ަ��r���~����E��[�C�Ӛ��(�y>Ҟ�>�7>c+�>_�>c�>����菉����&����ؾ"��2��*>��X���͙�����oн&�影P/�Rs?$�>S�`�
?9��q>��J>��ڽy>>��=�P�=]�J>8��>S��>�i1>`�\>|�=,]g>;�/��F�m���<�Q���$�=�6?�WӾ����J�#�]�T�`>[��>�RF>��-����9ݚ��?�̽�o��=��Z�=�2�>���>d�P>�>uPͼ����G���i��=*�
?��>�� �F�ƾ:�(2>�߱>۱��2�%>.L>T ?��~?�+6?(�=O?�>�=>�>�_>	�>��D>�,|>�?��?��,?o��>u�=�~���f�=�)>����g=]���V �������Z!�z��P˸p4���2�<��=)��=$3;p����&�2`�>dN,?j�?B��>�8B�9� ���x��my=�Xk>��]?�>�> �?�#`>�H�>U��>vfӼ�%��Oξ��>��>�x��.l��CA=��&�kC��Xf*?jo?v����پ��B�>)���}H>@�P>�w?|v�>��>���=�s���ӿ���)�uN��bΑ�?��=��ֽ"y]�a>�=��J��#ҽ�Cj�&�>0��>�\b>��J>>m >@޼��?�f=`���X1>��<]Dg����7L�=����t�=��˺�h��v�I<%R����9=��`�	�|��<)��<�!%?v
?V����K��Fӡ�zL��3��/|>f��>�;?���>k�>�*ݾ�]�$v� Z��G?��9?��,?z6쾭��>����y�X��x�>bf�>e��>�����{=�|��e¾J/�>���>��>M�#>ǺW�H�j��;��YPy>�ʾ=w	6�R�}?�Ѓ?�T"�#��H=���h�^� �u��5��F!����!�E�ﾣ73��,$��;�4�̾4=��>���?o����m�>E��������k��4��i_<�f�=�`�>w�I=�,���0�-J���'�ef!<��P��k�=̗����>�|R?:�>)_?%>>MN�>y0Ͼ =?[�?��q�>B�>z��=��>`�.?x�>���>&��|�g>�6�䷗�@H>�ߠ�c���<>3<0>)|0;Hyg��U�=��W>|h� T���S���.���1��P���f�������>c�>?�$��N7�>B�>�a�>�<^K�;kI�>U�^�MR����>k|�>S��>��<?v9#?F½>+�[=z�\���/�V�=C��>E�?,�?�'���>�4��);[�#j�=��g�8ZG�^���NJ���S�(�G<�>K>|>�=�>��g?��Q?�+?>��.Yf��Ǌ�(rR���`�r��$Q?��L=Σm>�׾��־��r�C�5���H�8���F��諼O@}>�˫�,�\>��_>�FR�YS>΀���g��U��=�M��W�+?Rґ;�_�>(�?���Y�:�Ծv�J?�l��1��Ʃ�U�ھm��J�>R�T>+����?�}��0^{��롿�^B�I��>w��?���?�e?��2�����$z>�X>F�>��<p�U�1���B��f2>���=L!���ϟ��F���R>��o>�LȽ0�ξ)�㾣�[��	����o�-o9�<ͩ��������>�X�P;!	���%�;��������M�Md$����I�$����}Ħ�Tm��.�?T
O?�k�G���-���ھⳒ�,�=J}ɾڭ����C���}����#���[�\º����+���+��/?Gd �*7���v���)о.�}>�)�>�~?m�Ծ؏�N��(�"��ò>���>����0et�,�������10?|Q?*o�ps��*8;�%T-=�F�>�)�>c�>�qG������>_�?�S?t�ds�%͗��h�A��?W��?+NK?������T��W-����jj?�&-?b&?��ǾZ�뾐��=�&?��8?�>ho�EU��(���^*?a-j?r����X�>���>�X�>��|�Kӵ�~ߊ<�7����Q�&�>�b->�g|������������>��?��j�ˌ�����>��	�n�d�cT����������Q>��?�(��l4>���>���=P>�`t���ꗿ� =��U?�O�?߫X?�-?����|ھ��� f�=�!>>�ǅ>	�цB�A��>�	�>s��+�x�9#(����>���?f��?�J?^�i��Mп�����Y���)����=p�r=�G>]j��Aw=�DH=e+����;��=�q�>���>1�y>��P>��8>/�9>c��@�"�.���eÑ���G�b�"�����l������w�����ù���Ͼ��ýG�m��?T���-��{�$�3�����f�v>v"�>�>���>�G�>zx>�9!=w���6s�&xݾ��(ా����/N�������E��������$��( P���C?ז9<���[!?Uy��1�>MF>c�|��:(=�#>F��>��>X=i>9/�>S8i>U�r>GN켢г>��ؾ皿|򑿑&��9R>)>4
6?52�~S�R����[�Ҿc��; ��>>��> a*�#�����d�?��M����s��ZO�>�~�>��>��>��0=�ek>�BO�R�������ba�>�?4e����Ӿ&=I�D�)>���>�ӛ���>!�>+�?=�p?a20?s�8��q�>`�s>J]=��=�Ո=��>x��>f?��$?��?[N�>Ӣ>+,o���=>�,J>����	�����Ov��!�R"b=����$�<��X0L<�N=�=5�<��>���oo�>�F5?o?.�>�˅�I`��7t��3>iU?>v�=;�*?l|8>�8>?f%H>\N�>��>���<+}��ta澅�>�>*wt��C���3�� ������F?��l?�^A>b����>R��$�E=]�>�[=?��5?�Sl>�I=���3¿���8龜k$�Wپr������1�A�,F�;��߽ HS��S3��b�=uW�>�V>Jo>���>��=���>��>f��Am>^��<O�Q��A7�F��=�,���(;��=�&e;ϥ*<E��Z�̽���� �ὐc%=L�ý�%!?��?6Z��Z���v.}��Ⱦ�+��kV>X�?}A?4�>��>G����E���I�'뗼�dV?R�V?�b?ゕ�5�=��#����=./�>�>٠�>�V�0Ͼ<�����Լjٔ>K��>n��> �H=��`��AO��);�A�>6��=L��{S}?E�Z?j����=,v׾�d��F��uN�0&-==����N=��~K����\��RҾ	I]=(��>���?	(;�\Y>Adƾ�ᮿ���}$ξeM5��G+>W?GGF>m;=&M�+&����Dj�4�k��,�>�*��%��>0�^?o�>�X?��E>�`?�-Ҿ��?
�>������>��^=�Y? ^?㒜>��>�@�yC>�.���ZD=���}=�g�=a��=S��=0I�]���S>�W	��ʼ�w^��Q���w�S����|���=,d�>��%?zI=uo�>��U>���WN;>	d�=��>�{d���r�� �=���>m�>?i�j?��?��F>��r��!���]#>L�,?m-�>˗?���<ך>�⤾锽��=G9ý}*��떾:�)���Q�T�c<�l;DZ�<�1�=�n/>��k?�//?��;?w°��
�_�s��m�ߙ���쑾��=�h�>k�_>&����������a�q�[�����L�)�ǽg<��4>���=i�G>��=�M�=(�l=�6�=M�۽���=�s��>���>t��>r�>SYG=����0��YH?�����/�o޹�)
�èŽ<�>�hg>�N��?C ��텿���G�R��#>���?��?UH�?� ��d��5��>\r>j�P>t�=`�s��+[���ɽ��>�t7=;����6����5��`�=�l�>�ʔ��'�3kᾟzI��}��F@j�\3K�n�_�B̾IY��Ad���ď=@*��0����Č�����5�ؐ�<^�y�%8;��Pm����*��?%?�n���������"��v埾��"=L�̾۱��1	��2,�r4U�4w �Vi
������ؒ��`C�a?���-U���"��������'>A��>�`?�W�e�����s��<�L>h�c>�_)��z�����"���G5?z?"���b֖��>��7.`�yM�>8�?�>\�� >�>Ԑ>��M?b�5?�@u=�>��>����">ڽ�?�t�?��M?>Ϻ��V�0�)�c��?"�)??��Ծ�Ծ�C'=a�?�-?s<�>���䴑��a���Q?�r?��>�t�>�]�>��g��.���e=q@���'N�"]�>�2�=�^V�M'��)٦��B����>{?�MJ��V��v��>����>z�N�X�6)�V�B��n>�
?�h���=}�c>�>�� ��b��H^��Zq��7C?,��?� \?e�=?�$�w���|�=�Z�=@�?��Q>�@��L����>?�S#��p����m/?Ӣ�?���?��e?�݁�7Sӿ_��@������*u�=��=�>>�߽D��=L?K=����5A�t>ѕ�>k$o>�*x>C�T>u<>��.>������#�Zä��Ғ�@VB�j�����pg��f	�8�x�h��״�⽾�̨�zݷ��ۓ�6�G�0��9�>��oh�RJ>�ޑ>��>��?P�L��I0>����4�1���+ᾝ�!�f���(���v�H�0=�5�=CP����fc���$�aA?�'�FW�=��>���;D�=���>K�=���>0>�S"=&�l>���>��>��>	�;>�L;[t�>l��<�͆�I�}��r1���0�ןr��:?�)l� ?��I5��H����
��>qb?B"U>��$�@�����t�*!�>����R�)ƽ.RS�D�~>�q�>��=&�=7y�b�����߽��>
0�>^>:�k��$����!��=��>Tپ���=��r>�(?�r?G�4?�}=�Ƹ>�^>�>���=�$K>ЙU>Oݒ>�_?�7?>00?E[�>v��=�6\�x&*=��"=\�K��.D��˽�	�x�ټ瓛<��h��+=��K=���;e9}=/�t=V{ȼ�X=< ��<vg�>�K?��>��>�.��$?��xF�<g���={z��q>"�>��>C	�>3)?�T�>��N�`�҃�=e�> ��>�Bi��w�h�f�M>]h�=f]S?�[?j�	;�?;������#���-k>Q��>h�4?Q3�>R>>�۽���.���_������Ᵹج3���l�����2�����Q<�<�g^���<a�>1�>#>ts�<�!=�/>\��>��>�e���'�A�u�~�n�L���8J=78g��J�=O��	��=�Ut����P6�� ����k��=߽2���>�<?=n��M|c>1(��W6��u@����>��Q?^�L�O�?��Q>{�<���t�e��WM�5 @?���?u�>�2��3>�Kr��-,<�=>��>y]���E�<"x�<E��7cF> �2?(z?/O�>W�/�f��H��LL
���(?�wK=�D��ď?�a]?A4�j������:�C�4���5=�'��x�g���M���.�M���l8���+n��`�=w`�>�?nj��nF�=��|�[��j��yF��RC=��=F�?�w_>�K���¾�� ���˾�c;���=�u�>�O��?ԃ?vRM?��N?(�>��*?V��qV�>���<-�<?���>wp? �>P	�>�Ml��'�<�ф�A��F�/����l >;NN��M>��>\2>Z���߉�j}?>�3�=������;ٙ=��k��|�=�SZ="R
>���=C�?[�?n���l'>o�|�b����>ES+>>!�݇���T��R��<��E>�A?W ?&��>�5 ��������oP�1�>F�>X�a?���>I{��4j.��b-��{���`^���>�8��׍�!�'��ɾ� ���>kE>z3�=��(>Wl�?��N?�N?T���J!��S-���(��	4=d������>>��>�>Xξ�N���b��=I���Z���������18�=��8>���=S޶>9�M����=~��<S�|��%H�	]�<�-=�ʗ>��h>���>�.>YӅ=S��Ͼ����C?<ٹ�k����
���Լ��=�Wz�,�>�M��?�[?�+���ㆿ,���j�A�S�>P��?u�?�-c?��>w��v�9>Vֻ<��=_�c�v��=�)x�p��=�y�>�e�>f�7���ʾ��]>��|>�!=ԥi�;H9�LA^�Ơ�����͚D���@2��g��iᾩl���NZ�G��=�孾"�Ľ����ؽ����}�9���;���|���]�?��q?���JMS��d��Q��tp���ٶ>���p�8��t־��ڼ6������桋��� �� 7�gvB����ۉ�>V���_!��<������
����=e�>?�|��ί�Z��X);>��>Dý=�I��"���H����(�dpO?ًi?�)���.�#1뽛j�>A<�>�\?:�8>B,�����rc	>�5?
:?��<�d��8Y��2��<4��?��?\=O?v�7���/� ������xu?�?�? g�Wq��.ľ��>��?��6?_*���(k���K���>ǎd?R�����>��?\Ad>���ՉϾ���>j������V>�L�������7���-�=��>�#�>T�A>⊹����/�>�	�6/*�!ϊ��C��]F�9��>V�>b��%�;`�>2@�>�0�~|���Y�� �"�(N:?�G�?�XY?�EZ?�Z�NL�b�=��>	�?�P>ԑ4�F3Ƚv��>?g?@���%���X��T?���?���?gqE?PV���ֿ�⓿�޽���0=>�O�=�>�=|~8��<�=�=�4ټ�E���L�=���>��0>�R>@'>E�='�5>�u��A`$�����m���!-��~�Ԗ$��I��t¾�p�h��&Ӳ���ž'#���r���s�ш=�#�4��,��S>���F>��v>���>��?O����{>�� �}��a@A=?�����>�uھ�+~�4�ɽ�q��ʺw�Atv��h��u���[[!���M?J1���=T>[_ü��.�Z�>���׵`����>xP>��>��>�j�>˱����e>do�:�O�> �Ƈ��{�sK� �=B���ϴ%?Xe:�ˤ�;m�=��p#�J����I�>��>?� �>F�&�*{��\�Y���>=
>{��s��%��⥭=��?D�T>.>��M�p����+�ݴ�>�.�>Gtݻ��Q��s).�ΐZ>���>�a־ď�=o^x>Ӳ(?_�u?(�5?���=
��>\#b>���>J�=eL>=DS>��>�%?/!9?11?U��>$v�=��a�/=b�:=|4B�W�8T��vPؼ��(�t<�"8�#GK==�p="<�f=�:P=�%м�d�;��<y��>��?��?dw�>j#��"�J��������߅=�,�����r>t��>�?Z�?(�>n�ֽ����T���Z�>I��>ɺP��&���ہ���Z>��>eɄ?�p?i���"=�y�������0>xi�>�=?8�>��X=��=��W������P��>��<n��Q�(��l:�ʜ'���ýRݫ=��X;�U<�1�>>���<\��<Ri>>�d>#��>A�>x���M�<@8!�����~ >�K�=�V��yh��S�<Xq�=58B;��
�w���l?��2�s^=��<��?�K?h��(ʽ�Qq�&��] ��f?�� ?f�=��?2i�=Hc�,܂��/V�(ꆾ��D?���?ğ�>4���s��=���Z<=��*>�D?=|=*�c��擾�Ͼ�=�=�7-?B�A?�I�>�c����{��D��R�Ҿmx�>>�9=��렘?Y_?�����~�&� ��G��O���#=��۽�aZ��ı���!�9�G �����%t����=�>(ݤ?��~���=eq��Ʋ���J��EU��JOl=x)i=}��>lD>�36�y"����J�Ѿ�tO�s�<yK�>'G��G?�n?mrZ?w�'?�;f>Y�?�o��U�>T��=��?���>+�;?��>T>�NL�8%�=saO�A�=����t��>p=����[>�>F/>�=��l=��=-�a<>
B���½������iw=~�y=u�>�V=�z?R�?�1O��>C~�woĽ2�Z>��x>�>�=�J=9���N�o�*>p�?a�?���>�J|����V��� ���r�>�F�>�J?��>s��ñ?<�,��6r��Y�>��?l�=f����<��0�����?���>T(=W8>>�h�?�O?i�E?�g����#�&HW���4�l�ν[�����>i��>2�>�����!���k��?���D�^���~Q����e=>g>Y��=ʉ>E��=�$�=Ӡ<���Լw# ���;G=�<�>�3�>g� ?�:�=_0�=R��|��[�P?0��f 9�,;��27>i�>$�ӽ��'�:'����;?PR#>�S��m���^�X?��?`t�?�;?L�m]���2=c�=VJ>��>��s��|�R�<��=��>hfƽ�	�x�>uc>���>rv��ھ��6G����R�$�,�I�Ҿ叓�)꾧Z~��Y�O�r����ڮʾ�/5�|�k�}�ҽA>t��KI�Ѣ��OG��sq����?"�?�D>�a��@0����=%��\ >��"�d��?��:V��;��?��W��Oc��F6���%������s�>r�����v��Q���L�u7ȼ�p >�7,?�ʾZ����+�eͫ<K]>\:�=����ҁ�$嘿����Ps?k&U?���������Vf�)�)h�>��?��>>����q�+�'>��G?ß:?#H�<�1��z0����ǽ�c�?��?eT?ȯ�=� '�L���Bܻ�Hf?:S�>�Y	?.�;ߥᾒ&��^C?��l?�F�>����m��Kah�.+`>�/h?*�.�Й~>p��>-��>Ѹ��5%=j'��Y�7��W�>��p�I�Z�Z�˾��(=�Fq>���>�,�=��	����<�>�=�5e8��g�֍���-b�W�W>�?a���h>�VL>F�_>�a���}�U���:�#�@?o�?=Mg?��W?ܹ�Y9!��Y��8E><9??�>,m<������>L��>�� ��^n�J
�p�*?8��?�� @�c]?�Iw�;.߿�럿jJ��������=��5=�]w>@���=��>�m��e��00>�ޑ>%ze>8t>>���=��->q\>����3,"�;���3!����(���1������Q_�����	�����(�[��{�fQýkn����9��8�|�Z��[>���>��>*��>ťo��ͷ=	0վk��]�m�g�ԾA��P⫾��ξ�l��` ���"�k�V>����s<�$��`?+�9�H�����>Ӗ3��#���^>�P��@>�Ď>�K�=F1�> Ӈ>(O�>� ^>o_=����đ�>AUx=�ʁ��{|�?�-���C���o�G�G?��=�����F�3�gᾑ���>��?�G�>�N$�O+���p��$�>���δR���	#㼹�>L��>
�=�  =J���v-��'����M�=Or>��>��H�%l��y��:�m=c��>a^ھț�=�Vz>��&?�s?U�1?�e�=���>$+\>0]�>xz�=��P>��_>M[�>�'?�`7?ʄ2?�Z�>�M�=Eg�V�%=Y[G=�F���^�@@���\���>����;TzB��>=�Ђ=�B�<��g=h�V=|���g:�,L�< ��>T��>���>���>E��PB��d<��b���:ͼ�!���hO=��֍�>P�O?�$?r�?��i;���W3R�L��>C��>�yr��;�,>�:f>�Ҁ>(}�?�8b?������Q������3 ���v>d� ?�9?�c>���ܻ����Ftǿ ���A,�S�<��;A�ۗ�������ƽl�=h�g��1�x�����_>/$�>;�">c�<=���=�QI=�L�>���>RR>x������K�ֽ�b����=1��=����Z�~<|�Ż���
^}��X|��V���[��R{=�
���1(�>ՏK?4"W��=����难��N�g�>8?*?��u�q��>�:>Ă0�ܾq��a`��A���(?A�s?��>�����>����u�ڽ[b�>8'?Q�}=n��=d*�<|z� (=��?�h5?�ه>Ƃ[�پW����FR��)�?�u=��	�m��?<!\?���ƞ���`��A��p&�6E,=��7��S`�+E��`�4�)�p���H�����a�$>Y/�>��?�#]���&>N�S�8����.��F���$p�=��>���>�|$=����0˾v���ʾ�I���=Xô>�A�sj�>i�?�q{?̨?�q>:l ?.f����=C�8>W�j?�>1�?�b<��=�HҼ�k�>���o���6�ʽ�2\����;|�L����=8z��$�>�rj=6gc=��=�����ٽ�'�f��E�����=�*=
\>�u�=�]?�.4?=��1�a��Q9���O��yL=��> �>#\�=�/�RM>��⽝t^>m�"?��?�%��~A�����(����>��6?�a?�{�>�}̽�C�b'�n��<��=��>c`佱�[�$$	����������>�
�><�>>݌R>X{�?ǘA?	�'?"�	��~!��i�)
,�Y3��,��;Ŕ�>�%�>��=�پ�q+��gl�TrL�y8��D��*�b�݋,=�*>�;'>Z��>���=�D>^2H�S5e�wዽG��;�1���>���> p?-]P>U(�=%&��a&���H?����I�����(墳7��=gJ�=J��>3��>	 '?��߽aч�J���9�4�M?g�?{h�?6�&?-�*��C�<�r�=
�(�tn�>\�ۺυ=�����h�j�=�;<��e��}վF�)>���>�ٝ>��r�K���j����j��Pÿ�M-�۞K����HG�e��2Wվ�JD��f�Ӧ*:k��AiN�!ߏ���Žc��-��ƾR���ù��?!�f?ND�=�ҽ������xgɾ�$�=F�]�J���$����I�t��۠��4�_��F�3��F3��v��o9�>���K�z��yo�0�꾞������s&?�ۇ�;\����ޮ=f�%>�S>����[�l�|��CQ�:O?�I?���0@��ѽ�>�j�>�\�>9V�>�_��\�v�=�I?d#O?��2>���90��N�h�0�?)�?��^?x���)����;�"�<��Z?��>ړ�>U��w1��Ծ��,?�Iu?�?����{���F�
��>�?��d��Ħ>�;s>[�>��־
�%�>�Mv��f���b>6�9�Nڮ�S�����q�Aǁ=5j>5M@>�̾~�8�?���es�OJ���U<pPӼ��=�+�>����y$[>Qu>���>�g���q�K��L���;?�%�?7�?@�/?�+���j�a>+� >+�>��=��i��=b��>���>��������7�0�?���?��@W�@?�F���!ֿp��$����7��`�]<��>���=׾����Ɩ=�]4=�)�3\N=$��>��R>�Q�=�G>
�5>�_>�߂��*��ѥ��_����*�K�꾂$��d�����;�ƾ�* ����O̾w�g�����a�q�w�+�ý�71���=�f��=�>��?j��>CЖ;�A>�Mᾱj?���н	8 ��:� �߾���CC�կ@����RT���� 
��>��zw=?${\���=���=�����|)�;��>�C>=r�;h�H>��=#�>e��=��>�>3J�>bP�=�>�i[>�t���~����K�=�n�=�u?��>����R.���i����e�>��?RB >��I��-��
�����>�Z�ڰ���k)��v�;��>+�>$�^>�O=>�q>���0�i�YQ�="}�>���>��>�4$�#� ���[��>)	־m��=9z>��(?�Cv?E�5?�}�=ʄ�>�a>]��>���=A�M>�P>=V�>�g?&P9?_#1?;�>/��=��a���=�P==O?��vU�<!������*���<D�4���D=�Km=��<Z�[=�L=�������;�=�c?'�L?�E�> �t>�f��}Q�$�[�a�.�(��>��оD��>���>9?�E�>��=���jQ���D���q�]�?c�>���0@���+X��+?D�?}��?jG1?8�1�pI=��S�;=*�>+�,?�(? )B?I~>�R����������Qk���S4�����Q[��i׽qH�F�{�[�]>�_<(�循3=9�>�#>x=�@j=�ܩ<�ԑ>N0�>�դ>�k�=9U=�༱�s����=�;>fƸ=�p�=Ӯ�=�{�=��Z=�>,<i�����*�<��;gj�������	?��1?3�<iЁ���Ծ�:V�����*?07�>�>˦?ir�=�5H��M��\�j�X�h��% ?���?1�>�_a�m�'>Re>�ZR>x�L>I��>�Ż��∾�M-��Ⓘ�R�=�7?�Q?���=O� �!������6��7�>C�;=��
�h�?"_?����� �0�G�ޘ��'=�2�`�[�c�����!���8�������!�r����==��>Z��?u~~��?�=K���%����U���k��cnp=v"l=��>��D>��7�&��>�s�о�vN��I�<Q��>���U��>?��?"=o?�yn?!��>�-:?��I��H�>��i���??��?-�F?���>��g>'���C�=�Ȩ��\!=טٽ<R��C�>Q��:��>.��=E�<����2���v>V�7=��X�1��/H[���ǽ�]�<�ӵ=�.C>d>G?��4?F����a(�Nx�>Po���(�>a�)>,:�<:Q��~[�>��>���>5&?�n>��d�q���{�o����=:�?�l?�?IC�3����D�&>���>pT1>�����#���޾�E���a�>�x>� �=�b>~m�?A�8?�1$?5\��6WL�ȷ�����ʛ=��P��^�>��>�f3�B�"���M��Ԉ��H_����w�0>�D�7>�==P�;ϧ[���u>�e)>���==K��Q��=H�W��t��os�<���>?M�>z�>}	>����e���;t��S�S?�޾���}��:���vm��g�A��<3��=D7?5��x���⫿KL�X?l��?芵?QV?@� ��� ����>�#<u+���[Q��ų;�m�>�'>/ϽL�]���Ӿ�X���uI>d��>�(��{�5U��Ȼ��ߴ���>��@�D�߾ >����ľ��m���Ͻ�咾1ɔ��H��ܸb��JG�D�D��5޽�}d����������G����?	��?� ��!X���#�?���̘�֟�>z��ˆ���ھ��7<BD�������˾����6A�F+���ܾ�>0�d�����܍�L��Kl�;���>iP?���m���
6��5">��V>�)>�W�����Ü��o
�C^t?5�w?^v�]�J�8�A��:�>#="?1�>�T'>�>��Pٽ3�#>�QJ?Z ,?��v�m���Wu�Y�\�Q��?`��?�W;?��]�=�?{ȾU/5��l?\��>Ar�>�e��uB���u}=�N%?c�E?�'�>�U��)��E�@��>�8N?>�����x>/0?�ʻ>��*�D���}�5>Mʓ�~��<'�Ļ��v:G�m�$%��!��1>�;>a!�>=�g�Wa��V��>7�
�D�+��W��o�{�\����>?O�?����V>�\�><ԟ>�N=��z�1㎿�3��7�f?"��? T?�iz?
�5��$3�>��<�1�>�s�>�>���;_�ܼVc?���>Oк�#�v��?���%?���? �?O�G?�ʂ�k^޿�x������N���r=j���$6>|ى�L��<1�F=�F���J�{�3>���>�J>�L_>��U>�_>��=a����E"��g��31����;�+h-�������ي��������t����ž�`>�������[�l�7���S�'R~�0�=�ɏ>���>/+�>�^�����;.�ؾ�ݾޭ�7����0	�Q�;N���8�����CM⽋��z�+�Ǵh<���bM5?V(���7����s>m�=|���1o>�ǻ�F�ٽǏ�=��>]L�>�B�>���>�=���>i�ܽCI�>�>R������Z�S�����<�\�.%?��S��zR��uT�����=���H?�??�L�>�x#�5���$����>.F>���;9�ý̵��$��>�>��[>���>����6����Z�|��>��>
f�=[I�"������� >h|�>	�׾�d�=��u>�C%?st?;*4?_��=��>	h>Lم>! �=4H>'�\>ȍ>b�?0�6?#1?�\�>"��=bY��/=	i=vgL�=	;�����jt��3 �}͵<Bi&��=~K=x�<�Fk=�]=]g���KU;²�<5f�>�q?���>��>����4���*�o�?��S>�
���>��&>�\�>?:��>��>��=��B�n��y�>��>W�N��ă�&�>�R�9>4��>i1{?��M?�k��[��<����Dl
���c>,��>�?<��>��>�hv�N��i�п����)�:��h���9/�GK��I����0ܼ�%��d޽�T=
|D> o'>�RQ>��B>:�=��=���>͋V>�|�=�t�=-��<)��N᩽�l�=�:3=I�	=�/J=�0�=̪�1���u�����k��`����H��=?�?��Q�kA���d��3��b����F ?��>����?U�u>�i���{�q�\�O�s��?N��?�|�>�=�W����!$��,�>*/?��>��>4��Ԍ�~`>�b?l--?�{l>Di޽}y��Ѐ���ʾ{�?/=���2��?~�_?y� ��e&��7F���#�'�j	��I�h������j!��(8�0�뾽���\�>~=���>�S�?����}=w���TF��)큿 G���/g=I��;���>�hA>Z12��>!�Wrھ��9�p=���>�B\�9?�Wn?�X[?B��>��'>�`>�6�ĺ�=�\={<9?(A?��H?>,��<��������!%��r�g���p�[�>�K����=��6=x%�=u��<��o�D
V=�،=���� X?�m ��Į;�p=י�<!�=�>��>�*'?�̻<���r�m�:f��;v��>��?{2>᭟��������u>��,?gk#?���=���b��ju
�[��>?L�>p�R?�>?�d�Ur��EN�#�;����>��=kϽ��(��="�����Q�>�̈́>G�Q��@�=C	z?AG?��O?\��R��Q��� ��_ֽpk�Z��>���>�e�>��ξP,�5io��F�u�0�X�q�)j�[�[<:,>j��=��<>/m��]�==�ӽ2u��`��e�=�L���Z�>��>���>���=+��=��7����0�P?*%�3<�����=�v=���=hl�<x܀=HCh���%?9HA�:�Z����f�G�?���?!��?Gj?2��;C;/�>�j�;�Uk>e3����<,�ʾ�0�<��V>l<T	�����|�=K�>��)?�z$��'�̎:��r:>�"¿�H�p����۾�	���������� �"�+��H ���ǾEg���n��p�U5��E��9��Ne��0��Ԙ?݃?�D�<����$�!��O	�����>ڤ��~�+��0��P\ҽYC��$p����龭s�lq)�Ue�bj;�>Z�f����������,�-\>��?�J۾�hþ��OG�<���=��=��3=��Uu���k��ol?�$T?7ƾ�t⾝����}�=�"?��?��>�sm����u>��H?v�?f\$:�����-��Za�<,1�?�n�?��X?�%��GH��߾J�=,�}?��?��#?Ff���S��(/5�?W
?$SC?'�?�����{��fZ���,>�H\?��y�ƨ�>,��>�>�G޾S�ž7%>�C�����[�c>�?A�$g���<��I
�=��u>QZr=�3Ѿ5𾗾�>����N�ҙH�:��Z��b�<E�?9��j>�ih>5�>��(��#��҉�%���L?4{�?DjS?�98?yr���w����@�=^ڦ>��>zH�=*��xڞ>j��>3���yr���Xi?�A�?m��?60Z?��m���۔�i���S�]��>�n�=���=Tײ���U��j�]�(=Gb�=O)F>dS>��$>M��>���>�0c>��>`���.$�J���E9����%�&�*u�[�:7�	�+;ξ�
�ߟ�&@��'�L�Q-/����u4!<4�����b��N�=�A�>���>�0�>��'>�y�>wK���ݾ@߾7���*Z�M��j8� �Ҫ��鮋���������Y.�Zh��q�>y�'>
~�=�\�>�"�=�m�=9t�>zF�>51Y>��&>��>/��>�E>M�>A\�>�A�>��7>_-y>�Ճ>o���Dr��/�V��y��am>R��?P=�b��x�p�g=�5��-��>��Z?_o�>�A�駿Sʟ�R�>ي">�;kd��.e�� =?��>�6>�Ci=]n���#��_���j(�h��=ۍ>)]�8����C[=��>�Z?�ҍ�h,�>]�>rM+?;��?��?URɽF�?�1?^�?2��=���>E�>9�>�(?��:?�1?�s=?[j�=�Z�2>n�㼙��b�f��r<���<�LT>��n=8�=�`�=�W���=��=��c=�E����={?_�6?b�>�Q�>�dg���4���7��'��c*>[�R>-�?�>	=?��>�b>�%
>;�=	���g��Z��>� �>p�0�\�e�	�S���=�.>Qz?�;?�3��U��BzQ>	��<�8x>d�?��7?at�>5��>6��=8����Ͽ�c��N0�Ւ�=}���I�<>�A8�?nǾ,O���5ȼ2;���L��P��=}	�>�Җ>12�>p��=,!�>�ȑ>Y�}>,�	>�6�Q�!=�s�IL˽x�=|�/=��������<ʼ'56��G�p�۽ոP�3���BH��T%?@k(?l��=r>3�#{��m���O\�es�>e:#?���>M�>���=�vʾn�0��&���k��S?4�?Z�1?��4��-e=G�l�!,�>_?�>�-A>E������)����;��%�>���>)�>dG ���Q���h���%����>�?�=��Ͻ�ǜ?�]?um*��ã�.,=�%�G�P��V���ǧ�����t�־��4�>[n�*j$��d�������Zy>�a�>R��?
ǽ���¾�꪿F���t˾��P'� �?Ga�<a0��.$���F�OCH�m�����H�>��{>�3�>x)?�e1?D(l?~�<?�<,?qfg���?���>O+?��k>��?q?��>נB>R�>�S>
>�j��⁃�Y��;�Բ=���>�A>Q�C>�I9�e�v��Ͻ=#��>sB>��!=efU=Qr�=5�>_r=�.W>��I>ƈ?`�$?���=��	>��<�ߕ��@��P2,�Of�>��ڻQ�n�@Qc�,ԓ>��)?&?jE�>���=�ؾ��X��/�2�>�9;?y�=?<w�>xF�>�>���
����H��W�>������X��R�{���>Ȧ�=d�=���>Ў?-3?���>���r�Pe����t�=�B��\���M�>쪥>��>Y����ml��My��G\���ľe�νNS3�M�l�'>��}>�*�=���=���#�<�uT= L�={��h�>ٜ?��(?S��>�;j>��U�4(���I?Š���������о�*#�b�>y�>>�� �g�?�
��u}�"����=�)p�>�v�?º�?�d?dVB�����#]>��V>0�>1z+<o%>��P�룃���5>�="�{�h앾��;F1\>�z>a�ǽF�ʾYr��=��:��s�X��b��ڼ�;w���=���ž��=ǿk��Ӧ�Q��X���p������#�������Z��Y������?�g?�=P�	���?��\!�;��*��>*��8x����+�]�Y�"��&?����i���پ.�.��VN����P�>V����ӓ��L���M�mxZ=Yn�>%`?"���u�LT=�]���=�G��Ey�-���A*��KJa��*2?K
?a�վ��"�ͧ>���=E�>�[>�~v=��������ł>?�?X�?�Zb�s2���x�������=�?���?3o7?mc��X;�AM	�U�b���>E�?,��>筘� ��HG���>�"?�nw>�
�5D���2���>SM?�����>��>N��>��*��⢾_��3ݾ�z��a'.>��=��9��1���T�|[@��0�>���>i�y�p=�����>|���qL�v�F��p���p)�<0��>�1�Q">��t>L�
>ap)�J׋�*�����KmL?�ʰ?�iT?��7?J1������I8�z=�Ǥ>���>�Q�=	��T��>�	�>j��,�o��M��?Q:�?,��?0+[?�k��Dӿ��������ѩ��!x=`RP=6�O>P�0��J,=Eɿ<
l���ۻ�eY$;qG�>6�[>>[�>q�\>$�J>��>?���k�)��-��I����U��$��)��Í�7u�	d�ײ��2��d���=������μ-Q��F��Q��
�T6�^{w>���>�.>bx>(7��g¾�wž*��4�-�|���H߾\���Sd�`����7���o�@Mh�%��#����>Wea>Kf =4��>���21��zø>ծ�>><�>�Y�>E�s>Wĸ>-К=�;�>���>I�?#T�>�����>e?���Ϳ�nY��B���|M�9D�?�uU>��B��� ��=2����B���;?KO�>��o�ĭ�)ÿ���>���=�g���
�aD���>�A?��S>�U���� �]f����}_F�PAC>~��=}E
�R���K���=�	?,����˽y'�>ĸ:?�S?A�@?c;���>�a?<?�� =�k�>ji�>,��>d�?��@?
�Q?��?�\>>��4�@�ӽa��=n��;E����0�=���=։��I`�<3N��d�> ��=�`;>a��=a��<����z��l�!��B�>�6K?Vp?�y�>�_��7�/���$�Pq3�C�>���=���>�d>	D�>��>�$�>B��>��>����ʖ�}m�>��=KT�{�������w;5�>*�b?�aB?΍;�����޿<���>g�?�1l?��?�q�>��7�T��e��2Y���6��Խ��K��n7����MA�e҂=ܫ����޾Ez̾}�>u��>��?>���;>}�=e�>k��>��;>��{>5<�=7x\=u��sɽ��2���߽�^[=��&G >ɸ������h����ѽ3+��H<���=�y?�?]�3=�O����ᾈh���h��a�>��>��><��>7s�[�����,�JC�V�<WJ?ׯk?{v�>+��pz=�#q����=��?�k�>��'<�5 >�2��p���]ν��>��>p�o>�����s�
Ԏ�m��][>3�����1���?�B?x(�c�+��+���Q�մ��t1�r�a�����s�,��K�{����Y�'�!���v�I��>��>Y�?�����F#�Z���'����������,�s8=��+?�>��'���$��l��c2��T����S�f��>'�>p�>|?+"?\f=?wT?z��>k�X�C�I>[�J>�2�>JKQ>!�U?)	?1��>�G>�5�>5>�{Ͻ1N�����=>�K��b5<�p>��;���wu�>إ >m]<j_
������0�2�%�T�:��=2.->��5>��:?��?O�=�VP>���=U� �
�+>u*>��0��HO>.N���RM>K�>%�'?:6 ?�]�>��A>F��� �辶���de�= X�>]'?�u�>^�/�Y6��m�˴c�\�<X`q>C����(�Ҿ�s�������>5��>�폽�� =�{�?j�A?2j�>�y��Ra��2闿R$p�0��J��r�>Mb�>��Z<�t0�D房�촿ԓ�U�F�]�G=�;-�
�|)�=�a�>��>���>�d.>&ý��q�2�����;�="?�?��I?�^�>+�>�"����2��??0e��� ������$��a�>�-6>#@¼�d?:;Ƚ
|�����5�Һ�>���?9�?�3d?X�.���y�;>V�4>�z�=��&�s*?�Zi)��H�W>b��=EG}��A���7#=�%u>?��>{t���Ѿ��ǾJ� �G�ÿK4����;�����W�f��������<-;�S���, A�0m�=@X
��6���?����F����h�p�D��?�9c?���=� *�ng��}׾�����>��˽����wAA��\���Y���K��+$Ž�t��˻��D�Ή&��S>i�ݽ���|�˿=�umy��;�>�s0?�����FH�V�(�i7�:5����оw~���x��<]��f�%?x��>� �R�����	>70�>�� ?�z>��i�ȡ�{e`��X�>'��>GL?�܇�R����	���3>yq�?��?ąC?��J�)=���������?��?R^�>��������փ����?~�7?+��>5���4Yz�t&��o�>p>R?�Ja�z�O>P��>���>�y��x�v�΃�x(��.���+�=��d������*�d$,�Q�=Ri�>��n>"P��n�¾��>`羣DN��tH��+��"��<�`?rg��>��h>�n>��(��\��������J%K?��?diS?p�6?�k���5�k蔽H��=��> ��>`�=fK���>���>��쾥*r��g���?E��?��?��X?<�m�(�����Q���N����X�>n��=:B�=����%2>��=��=%_c��>'�>L �>��>V2o>� i>��%>�S��,. �A���|������b뾸�.��d��F���Da�۰ݾ0j���T�3�B�C��O\#:��!�l�-�l�����n�x>s9�>$ز>�q4>*U>'��>��/��W��k�۾X�~��*�c��M�!����$�/�̼ܽ��P�J��:���q����>�^>d6@>���>c\����:=ϭP>KT>�m>�Z8>��>ݗ>��>�6�>q�>{/>$n�=�9I>fS>;��[^��a�ξ2l��4>��n?�L�k��`È�{ן=�����r>��?(*>�L�_2��}长�?�>��پ=_�=��?��?ˆ�>�E�̕�k���ѽ��=}�?>��J>&��M�����?t�<�z�>X��r�*>�>�?���?�/)?D*���p>���>�>]t$>r�?���93oh>�j-?��;?�3?�w?��H>����x�H>�@�<����|�=�=�:M���Iљ>��C���>=0�f=��@>���:d�A>w�?���\>+j>K?)?���>i�?ʸ���3��I����� �>K��>$�>���>-�*?P_�>S�>�?�>5��>`�U�~Y���>��>���|x�-~㾃g=��(>��c?"q?\#M=ĝ+��)�"+H���>nS-?>�/?���>��>a3w�o����ʿ�����}1�=�͒������>��齶�4=�3��p�	$�
��>�Yw>��w>��i>�v�=�r>���>9t">����C�<�O�<P���>�c�=^���=�-��K�9>F������o�����=�8k<���9�^�?��?���C/����o�
N���Z���G�>���>ׂ�>(��>��=r�7�T�9	<���9����>h?*9�>Y�;��H�=��F�C<��>݄�>� >=災���l�����a<���>�?z�>���IY���l��A
��^�>��=Fl� ��?� Q?7�7�����}̾�#3���5�0��<����Q����Y���.���n�/
�u����i6�Ex�>�C�>V�?ݽ|�~�<pu�����O͒�����=���7d?��>��ž����bX��0�V��O&��U�>�=�h�>�v?֎?�@k?9?)� ?a�G��8�>�jv=���>���>h�?��?h��>���>�R�>ݳ�=ۀ��ML뽘b��#�˼��^���=�`L>�G>
Y�=#�(=C��=��q;z.��ًļ_��9<0n=���=�#>��O>o?��!?��=�7>�f��㠾��X��Ҙ=Z?<ό>nT�=��8��Ñ>���>�M?�? ?�j�>� `�\� �پ���� ?�(?X?�%K>�^>l ��n˾5f�=B�_>x�ٺPR�I���������K�L>�E_>D��=���>���?�EF?š?<B��$I��z|��eZ��	6=�'ͽ���>� �=�2��G��V�_���[�eIK��-`���<����̻�<�>�>څ�>��}=�$=�	�<(\=��^�����4j��>���>U�1?��>�S >��u� [���I?�*��p��8B��A�Ҿ��6��'>b/=>����?�D�/.}�������;�'L�>���?���?�Fd?�
G�}��x�\>�WY>:>s�h<,c=�]�'G��f�1>3g�=cx��앾�6;;�%Z>w>a�ʽ�!ʾ����v@�=f��o�Q�ln���@���
&���	}�FN?�wU������ƾEfn�6��x҂>9�����[���c�;�C!��^��?( T?m��<�q޽�2�@��S����6D>�;T���}����,��=�*��?Yؽ���:�ZN3���L��*�2�>ޭ��3������Ҿ�+�><"�>j�v?�	�� �!�F���>����c�=]�{��{���Q��T3���?��?�-ɾ�B��f�;pf=��>wB->^O8>=x��U		�o}?�a.?&�=?(�;�u���������<J�?�?/c,?sBջ\<�D�)�(�����>Z?��?�b׾i�/5޽R+?HI?�7>+������5�_�?�Wc?1P��6R->�?�w?�����澈㛽�]���>�j>K�>垳�Ю��1q��j'���>d�>R�����y����>����N�ҙH�:��Z��b�<E�?9��j>�ih>5�>��(��#��҉�%���L?4{�?DjS?�98?yr���w����@�=^ڦ>��>zH�=*��xڞ>j��>3���yr���Xi?�A�?m��?60Z?��m���۔�i���S�]��>�n�=���=Tײ���U��j�]�(=Gb�=O)F>dS>��$>M��>���>�0c>��>`���.$�J���E9����%�&�*u�[�:7�	�+;ξ�
�ߟ�&@��'�L�Q-/����u4!<4�����b��N�=�A�>���>�0�>��'>�y�>wK���ݾ@߾7���*Z�M��j8� �Ҫ��鮋���������Y.�Zh��q�>y�'>
~�=�\�>�"�=�m�=9t�>zF�>51Y>��&>��>/��>�E>M�>A\�>�A�>��7>_-y>�Ճ>o���Dr��/�V��y��am>R��?P=�b��x�p�g=�5��-��>��Z?_o�>�A�駿Sʟ�R�>ي">�;kd��.e�� =?��>�6>�Ci=]n���#��_���j(�h��=ۍ>)]�8����C[=��>�Z?�ҍ�h,�>]�>rM+?;��?��?URɽF�?�1?^�?2��=���>E�>9�>�(?��:?�1?�s=?[j�=�Z�2>n�㼙��b�f��r<���<�LT>��n=8�=�`�=�W���=��=��c=�E����={?_�6?b�>�Q�>�dg���4���7��'��c*>[�R>-�?�>	=?��>�b>�%
>;�=	���g��Z��>� �>p�0�\�e�	�S���=�.>Qz?�;?�3��U��BzQ>	��<�8x>d�?��7?at�>5��>6��=8����Ͽ�c��N0�Ւ�=}���I�<>�A8�?nǾ,O���5ȼ2;���L��P��=}	�>�Җ>12�>p��=,!�>�ȑ>Y�}>,�	>�6�Q�!=�s�IL˽x�=|�/=��������<ʼ'56��G�p�۽ոP�3���BH��T%?@k(?l��=r>3�#{��m���O\�es�>e:#?���>M�>���=�vʾn�0��&���k��S?4�?Z�1?��4��-e=G�l�!,�>_?�>�-A>E������)����;��%�>���>)�>dG ���Q���h���%����>�?�=��Ͻ�ǜ?�]?um*��ã�.,=�%�G�P��V���ǧ�����t�־��4�>[n�*j$��d�������Zy>�a�>R��?
ǽ���¾�꪿F���t˾��P'� �?Ga�<a0��.$���F�OCH�m�����H�>��{>�3�>x)?�e1?D(l?~�<?�<,?qfg���?���>O+?��k>��?q?��>נB>R�>�S>
>�j��⁃�Y��;�Բ=���>�A>Q�C>�I9�e�v��Ͻ=#��>sB>��!=efU=Qr�=5�>_r=�.W>��I>ƈ?`�$?���=��	>��<�ߕ��@��P2,�Of�>��ڻQ�n�@Qc�,ԓ>��)?&?jE�>���=�ؾ��X��/�2�>�9;?y�=?<w�>xF�>�>���
����H��W�>������X��R�{���>Ȧ�=d�=���>Ў?-3?���>���r�Pe����t�=�B��\���M�>쪥>��>Y����ml��My��G\���ľe�νNS3�M�l�'>��}>�*�=���=���#�<�uT= L�={��h�>ٜ?��(?S��>�;j>��U�4(���I?Š���������о�*#�b�>y�>>�� �g�?�
��u}�"����=�)p�>�v�?º�?�d?dVB�����#]>��V>0�>1z+<o%>��P�룃���5>�="�{�h앾��;F1\>�z>a�ǽF�ʾYr��=��:��s�X��b��ڼ�;w���=���ž��=ǿk��Ӧ�Q��X���p������#�������Z��Y������?�g?�=P�	���?��\!�;��*��>*��8x����+�]�Y�"��&?����i���پ.�.��VN����P�>V����ӓ��L���M�mxZ=Yn�>%`?"���u�LT=�]���=�G��Ey�-���A*��KJa��*2?K
?a�վ��"�ͧ>���=E�>�[>�~v=��������ł>?�?X�?�Zb�s2���x�������=�?���?3o7?mc��X;�AM	�U�b���>E�?,��>筘� ��HG���>�"?�nw>�
�5D���2���>SM?�����>��>N��>��*��⢾_��3ݾ�z��a'.>��=��9��1���T�|[@��0�>���>i�y�p=�����>|���qL�v�F��p���p)�<0��>�1�Q">��t>L�
>ap)�J׋�*�����KmL?�ʰ?�iT?��7?J1������I8�z=�Ǥ>���>�Q�=	��T��>�	�>j��,�o��M��?Q:�?,��?0+[?�k��Dӿ��������ѩ��!x=`RP=6�O>P�0��J,=Eɿ<
l���ۻ�eY$;qG�>6�[>>[�>q�\>$�J>��>?���k�)��-��I����U��$��)��Í�7u�	d�ײ��2��d���=������μ-Q��F��Q��
�T6�^{w>���>�.>bx>(7��g¾�wž*��4�-�|���H߾\���Sd�`����7���o�@Mh�%��#����>Wea>Kf =4��>���21��zø>ծ�>><�>�Y�>E�s>Wĸ>-К=�;�>���>I�?#T�>�����>e?���Ϳ�nY��B���|M�9D�?�uU>��B��� ��=2����B���;?KO�>��o�ĭ�)ÿ���>���=�g���
�aD���>�A?��S>�U���� �]f����}_F�PAC>~��=}E
�R���K���=�	?,����˽y'�>ĸ:?�S?A�@?c;���>�a?<?�� =�k�>ji�>,��>d�?��@?
�Q?��?�\>>��4�@�ӽa��=n��;E����0�=���=։��I`�<3N��d�> ��=�`;>a��=a��<����z��l�!��B�>�6K?Vp?�y�>�_��7�/���$�Pq3�C�>���=���>�d>	D�>��>�$�>B��>��>����ʖ�}m�>��=KT�{�������w;5�>*�b?�aB?΍;�����޿<���>g�?�1l?��?�q�>��7�T��e��2Y���6��Խ��K��n7����MA�e҂=ܫ����޾Ez̾}�>u��>��?>���;>}�=e�>k��>��;>��{>5<�=7x\=u��sɽ��2���߽�^[=��&G >ɸ������h����ѽ3+��H<���=�y?�?]�3=�O����ᾈh���h��a�>��>��><��>7s�[�����,�JC�V�<WJ?ׯk?{v�>+��pz=�#q����=��?�k�>��'<�5 >�2��p���]ν��>��>p�o>�����s�
Ԏ�m��][>3�����1���?�B?x(�c�+��+���Q�մ��t1�r�a�����s�,��K�{����Y�'�!���v�I��>��>Y�?�����F#�Z���'����������,�s8=��+?�>��'���$��l��c2��T����S�f��>'�>p�>|?+"?\f=?wT?z��>k�X�C�I>[�J>�2�>JKQ>!�U?)	?1��>�G>�5�>5>�{Ͻ1N�����=>�K��b5<�p>��;���wu�>إ >m]<j_
������0�2�%�T�:��=2.->��5>��:?��?O�=�VP>���=U� �
�+>u*>��0��HO>.N���RM>K�>%�'?:6 ?�]�>��A>F��� �辶���de�= X�>]'?�u�>^�/�Y6��m�˴c�\�<X`q>C����(�Ҿ�s�������>5��>�폽�� =�{�?j�A?2j�>�y��Ra��2闿R$p�0��J��r�>Mb�>��Z<�t0�D房�촿ԓ�U�F�]�G=�;-�
�|)�=�a�>��>���>�d.>&ý��q�2�����;�="?�?��I?�^�>+�>�"����2��??0e��� ������$��a�>�-6>#@¼�d?:;Ƚ
|�����5�Һ�>���?9�?�3d?X�.���y�;>V�4>�z�=��&�s*?�Zi)��H�W>b��=EG}��A���7#=�%u>?��>{t���Ѿ��ǾJ� �G�ÿK4����;�����W�f��������<-;�S���, A�0m�=@X
��6���?����F����h�p�D��?�9c?���=� *�ng��}׾�����>��˽����wAA��\���Y���K��+$Ž�t��˻��D�Ή&��S>i�ݽ���|�˿=�umy��;�>�s0?�����FH�V�(�i7�:5����оw~���x��<]��f�%?x��>� �R�����	>70�>�� ?�z>��i�ȡ�{e`��X�>'��>GL?�܇�R����	���3>yq�?��?ąC?��J�)=���������?��?R^�>��������փ����?~�7?+��>5���4Yz�t&��o�>p>R?�Ja�z�O>P��>���>�y��x�v�΃�x(��.���+�=��d������*�d$,�Q�=Ri�>��n>"P��n�¾�?�����v�;��S��C��z��>�z>�1F��{�>V�>>��>�7R"�)�c�|Σ�g�X�j?���?�{?�G?x��0���N�>ݒ=���>0֞>��=2�i�M3�>���>��{_�~>���>���?�1@�~y?�����ԿV������O�˾��=���=���=�	��o�%>kf���'>6�M>�>:�>mQ>��8> ��=VTL>?O>,����n)�E3��p����mI�c���7���[��,��7���?�w��F���z����O�Ž��W�;� ��	�ds:����=Ӗ}>W1�=���>�v;��>�z���s���ֽ���~Os�P��Ix����q��N��98w�Z���������)�,?����k79>�p�=�a�=W��=�3�>���>Y!�=�L��ռa�>�\�=q�+>�m&>F��>�p>�03>
e)=����k���A�I���1~>�^K?����󦽱�6��G�좾��>R`�>m0=͑#�����$a^����>r>i�ݽ�C��$�t;>J��>0(/��,�����
���M���0:��>4��<Z��~���&	Q�P�<b_�>��׾��T>�%�=�0?�h?��%?gk�=���>�w>��0>���=ݷ=a��=�>�0?�?@?}�9?ّ�>��=�x���c�=�E >�g���̽��}�;�:Խ�'>�B���9>ѹV=�=���=x�<��z��;�8]��U?��D?k��>��'?l4��`�1N#���U>��=��ҽ�"?�w>>��S?��/?�?�d�=B��߂'�-k��m�>%�>%4��ɱT�87t�S�=���>N�?�w?�a�;N^���R�������>��#?�,?���>�*�>�y\�=����ܿ0��ּL��6=<�&.>,)Ҽ:����->Y4�����<�o�>)�>!hp>^��>Q�U>��!=)�=�C>���>�2>F =7,S=�6=��=5ׇ<J0�=�߽~�f��r׽:�˽GID��9�I�z�Ԓ���Z=�y�M>.��|?�(?,^�=Hӄ=��5�tEվ����p>V$�>y�B>9�>�ל;��-�k9n�7�?�c�_�FW�>F�j?3�>���Hj>G ��r+~�|f?�چ>��e=��> ~=ok��>H[�>#?9�M>�+W�p�Q�+�r�~����:>���=�������?x�K?���_��G�q�-��L�����>T�->7�k;ܾ��2�}8��p˾���Y
ӽ�(Ͻ�h�>�$�?�~���@�>�m�fӊ��ˇ��h���y8�(�VN2?v���=�.Bl���H�v:�S��~A�+PR>L[>^j�>�#?un�>A�w?9�e?%��>��f�`eH?�<��?�:?ʓ??H9(?�O?(a�>^I���	���Z��OF��v樽<h��ОL>ß�>nA	>�l
>o�t=�9�<�,�;�=�*��]�a�;F��S~<�u�=��m>�y�>E�?��=?�o�<:
�=�X��w�8�>m��><j><���8F�=�_u<`"�>�D?�k?ED�>���ep�����ݾ�d<�6�(?��>�?LLy>��%��<�~G3<�2��vl=�>m��З�C���j=y3>?2K>�ę=�Ռ>�.o?�h?�F?�t&�78����5��mK?>rD�P��>{��>���վK^*��@��6�c�,	��>��b:A�;��=�g>ON�=���<�:�>nL����N!:�X���c=h�?��?#�?yJ>�%%�,�	�ZД�дh?�ԋ�|DA�7�B>d��|��>6m�>��ﾑ*��i�E?I�6�2��Ҭ�����o"�=6�?�v�?�Z�?ԣ^>e3���/�>I��>���=��,�I���P%�q�>�'�Mg	��?<u|����TO�>�H��{�@󾄄��z&��3r[��y��E1�p����~�9�*4�=����'Ȃ�~ ߾�N@���
�V��a��0P����������=�QK�?`��?b3A��]�֋L���+������K>~�7��� >�ӛ��e���A��U�?���ƾVF��U2��g��rپX��>)5������n��Y��a-�y��>.��>l��x��%�.�0�ӽޝa=1�b=CJ"�T����J��KHj����?+A?�ω�/j��+��H]7=�e?!Il>��2��0q��ؽ�]�>�R?iA/?�e߽J���*튿q�(��d�?���?'�??��N��A���w{���?6�?�>�슾N�̾(�p�
?��9?>��>���MN��m�?v�>�?[?l_N�s�a>�!�>U�>�����'�(l���"��^9>�]
��.���g��[>���=�
�>Rxx>�\�L̮��٫>�+��Y���$Nm�����a���=Cs[>��2�bS�>DV$<�\���5�)������X�g���m?[��?�5>?�H?�׾ۈ��[s>c\;>	��>��>��>;Q$�)��>Q*?��o��av��
���>�Y�?�	@�x\?���-�ѿ�󤿧5ξ(���>�5>&�&>[u��`�=rǽ(�=y�2>��b>��>$qR>�ҋ>�yp>�k>V��>�U��TQ-����������)�W�u�cK�����v��\@�Ys��ځ���5� M�o`=����(P��b=���s�=�X�>
47>(�K?^g�>6��=H�)������?��͌�����ƾA��5��C�+�D�����z,�<�?������D?
簽��)>���>%�=���2>)�5>I���{>��?h�.>�J?�!>y����}���5>�X�<���=5��;��T&��]�=��rI�TrF>�&*?%γ�P�a����%�m���>{�>xg�=�d7�G痿oV����>�򵽍�b�^���l�<���>�3�>�>=��,����"s����h���B��-m>]�_>dYI=�5[�6� ��:�h�>�{ʾ5]�=ήa>�W)?�x?5?��~=3��>�O>��>��=6�e>�d>D��>�?�e5?Dg0?���>=��=4�K�=�&<P1�<�HK�YÑ�G���~@��8�o�=�r!�f�=��=N��:�3=��S=��9B<���<͎?��O?�K�>C^>>@�ξ���D���a���0>��7�=��>%H
?��?�B,?�?��N<�G�� l�U�ӾGǳ>��>�a�	o�0Z�<-#"��A]=�:Y?Z$??���V�T�R�=�/>hV�>a��>�0?�(�>B4�=�.U���������a�H��>�{�=�)�<O:��ܽỀ�g��'|P=��>��>�D�>۾�>D�	>���=�d>�(�>�>p�~=�L�=dÎ���黦�D=��M��0��5Z=�SM��7S�+ۼ�l�l��L��W;��S|��gQ��
?��?�_�=h� �y֌��C8��g�@��>)�>Z6?�i?��<�;���P�&=�!������>��K?��>�I���=N���Dc����>�d�>-B>h�~�d�Iv�8Z�=Vv�>��%?�n�>��O�EQ��!g�7�߾�Ĉ>$��=������?Ts)?�A��ם�4�;����w �:$;�,a�=�Ѽ����4���E5��c������{�6�=?��>y��?�؆�rw>�y-��î��I��JB�	U9=Y<1>�:C?lL��ھ�η��@�ٸ߾\�}y=���>	�>���>�&?/��>#Z?�C!?���>�> pA?�;�/�>�"?]<?��$?t!H?vD,>��<B�H����x���(���s<lS��^�=�S�=�i�=�+���.>�U>Y���@M=e{0����� ��ɱ=��=�Ʌ=\�j>f�$? �@?�5!=^��w"���X��5=���>v?��۽)wS=�k�>�_�>�7?�CO?�m�>�\j�ǎҾg�������q�?	.+?S< ?�>'�>�z��E�@�fr>f��>I�I�����ꪪ��Ń�ޘ��}�>�;>Ƌ��/ۆ>ܖL?��]?�R?Z!����d������cْ>�}><�?=@>�⨾�_���� �z�f�uK�]
�\|P=�Z�����j=�ы>i�>t�>ƨc>��������}�ϯ�/pW=<R?Ep�>��?��F>Ih��cƷ���Ӿ90?5�_��y�{��=$���Gb0>_�?���O�%�/�_?�'��Ր�I���Cw��ڜ~��U�?}v�?�ܖ?��=��Y��*_>>�>(�>�ڦ=L�����c.6��Ƞ>]���N�����hA=���< ��>˯ʽ,@�$��̍�=!A���fW�^EZ��ƾ�õ�7ƹ��m]����@���F� �qǪ�5N��5(��a ��(S�QI���b���6Ͼ/J�����?o�?�r�<��AM=�����*\���=rX����=�g�H��]-�;����������Y�F��B���;��>qm��u��e�n��5��=���>�	�>֣�u�!��*��}��� >�������5쉿������1����?q�R?A��@)�y���MO�<���>�� >N���9�`�p��<���<�n0?��?��%.��������=���?���?��E?P2	�4�9��w�;%��N?'*?֏�>B>����¾ގ��9)
?�m@?7��>�k�~����$�>��\?�c4��Sw>Ai�>E1�> �<�K��̶����=!�s>�Vt<�U�]�G�Jw-��ZJ=W]�>jue>0�c��?��|��>�{���Pn�#�I���ؾqC�:�=��^>�'�A�>4>�=P��D��Fx������j��b2v?��?NyM?�&?y���[�վZ>&��<V3>4x�>�m�=�잾K%>�?��˾�熿)��u~>��?�U@��^?V���e�Կ~��������$�c��<-E�=���=n����<\���<�<3�;��}=%˫>�[�>���>�*>G�=�D>�����^'�錄����wI��v4�L,��������վ����ɾj[����K=��j={���`���h�z���{����-=���>sTY>�p	?�Q^>͙>t<��m�ͅ���uM>�μ�����S��g�����ux������M�;��!���?��ql0>�>_5�����=ڨE>(�>�]�<��?xc�=��>����}�=ϯ�>�\P>���4jh>o{�=[}|�^Bk��+T�s���� >S!??Cjc���A�������%>����>���>C�J>"U/��ۍ��Ex�ʜ�>�{��?R� �����=뀀>���>��	�?b�<�����O��.PB���z�hx>��:S�?=��K��'���7=���>*�׾�%>�4S>:\.?Kt?�i2?��=��>B�b>'%�>^�=��A>CR>�+v>]�?\+9??�0?iF�>/�=Oe���K=�(�=��K��蠽����p�>����O=��v�d=�M�=�=�>=
={96�H��E)$=�]?�L?t �>Y�>�3��!�q�����>:�o>�m�=R�>���>���>n�#?
.?>�|�
���
�ϡ�>���>���#����͇�^6!=�t�>ui�?	�-?Q���𢾧ܯ���x��s�>ZS5?�(D?<i�>?�>B��tL���ۿS:��NX�lu���\���?�����$����a��v�Ľ#9�>���>
��>��D>�@=��d�Ko=V_ ?">�=�]R��y>�_:�5��<�;�<�C2=�仼/�|>�ī��W�?�=��ݽw�2�����`(�]��=���<�?��?lW���%��s׽�����é�@ј>���>�8�>��>q�����U�t�A��"�_S?��U?��?^����M=yr5=}0!���?j!�>�o>�U=>lZ��7���2>�k�>��?Ԑ�>O� �35���~��Q�s!>$�=��ɽy;�?�'+?u�龰���U�;���*����\��=��==�;����k�*��W�s?"��h���a��[C�>4��?�竾�m)>����ߘ��֠��,վ<�>��<.4?
H=4�þ�	�������o[��"�=(7�>]�>�>�%?0?���?���?~�>�5�=�C?�#m��^?��=?�%W?>t9?�M?@�J>��=�м���.�x�d��q�=�w��P�=9�=*k�=c��De<[kL=�z�թ�ң����z��3L���%��~�<s6�=���=a�;?��R?o�J��9�Rd�+-N�q�>�!?M��>u���Ω�=[L�>um�>�+?� K?��>~�,=ڮF���o�˞н�?V�9?B?� �>�]�����{���m�Qá>��>��j=閊�8O�n�6]>�q�=R��=��>�{a?�|?�T?�w�mc&�O�����#��κ>�>��A?:S?�`��E������{��q����J>{���l4�<���=�V�>�(=���=�i�>5(>����{���尽$w$=b�>��?C	,?��=>�Ă<�Ш��ŕ��>?+UȽ�0���;��bς��l?�ƾp�-�e�K?bM��K��Ο��������+���?�?�?#S�?{�l>�H���N>�s	?e��=W2��fT��O"N��ν���>�v=�y�^�*�Y��̖���x�>����E�R�)���*>�I����N�ܝ���ؾ��Ͼ�2����g�1^���ț���=����щ��9h�0؅��h���"m�$���Gn���y��H��?>9�?U2>���1�J�?)���F�(躆yȾf �<De:�I������VԾ�M�Y
����:�V<�`����>W�4�k����a����v>��)|>g�>]���!8���7����9'>O��<����d������J�ڽ�rn?��??���/q��ʜ�E��=,�2?Er�>!�=����5�<�K�>��4?Q?�-��Dx�������u=K�?��?8B>?>�>�w�B�F������?��?(.�>���[/þ���j?a0:?F�>�����������s�>#+[?q�H�8�b>���>�H�>�ҽ,���+�x��GW�S�;>�]|;]�$��=_�G�9�j3�=9��>v�z>�N�;@��t�>�Ḿ�|����|�쮽ڬ׾�03>ȯ>TJ�^�F>��O�" ���]�p�x�� ���:�m�}?���?I9�?h�??�g�<i�0�zľ*��<�F�=��w>�<�>��F�]>���>߬��aI��m�G����<�*�?�@�2s?�=e���׿!ѣ�����Ӿ7V�=��2<�I>�5��a9�=p��=�15��@�OH�=� �>h�M>�<�>Ǧ>->xz>���1�2�����ܞ���4�������)aj�ݺ4�IT�����]��e���6�G���@���t��)�H�}�����U�=�{�>g]�>���>�%�=*!�<I^�����Q����q��/1��/�"���r혾޽�H��GxE��g�oQ���s?�T�=�o�=q�?�߽���=��>c40>�M]=o=�oC>{��=�&!>�q>=��=�^�>��=2�f>��<=I��<I����4�i�`����<NH?�Cv��L��M�1�#\߾�r�����>��?22>G'��쐿�ol��9�>0�]� ,`��ǈ���ݼ��t>���>>��=o�μ�8��/Y�������=�-�>���=㽼*������=���>��ľ�k�>te�>2C?�}�?�x?7�
6�>?B�<��^>��>0��>�U>hΞ>�t�>%�?c�?�$?�f�=�$'�B0�<�!=B�;�LI޽R]��7��N2O��[>�Լ8��<7?=�G�=n��*[�<KF���9�;:�F�?�4M?2�>4	?J�%�6"��5V��T��%|�>߀�=6�>�I�>�??��>��%���VT.�1�;���>ɼ�>��G�LP�ܭ-���=?��>��V?,��>��`�����>w�2�d��>�/?�?Bi�>N��>�.H�~�q�߿���Lۀ�p_�U<j�;п���9��[ּ�r����;r�⽊>��>�a>���<K;��޷����>���>�J;��1�<���<M�9=�
�
�=|Ѥ��Ɇ<�̽��;=��=�A��f�8���ٽ���<������-��y�>?��>�w�;��:��b��[���r�W��>5J�>�!X>��W�b�27����M$L�FF���>|�_?��>T=���1��=̫>�N�>�R�>���(mG��7>Ձн}M�=��><�:?��k>[�\�\�t� ���x���n;>A>=h���FI�?�LX?	���^���B���K��ѣ�Z`�>�	���<¾65|�KT��(U�xJ�� ��e��A!>�T?��?�6p��8V>�/��	���*� d��b�k���9>t�*?���>�q>Ӻٻ����ؤ�-��C���a��>4�~>�V�=�Y??a6[?�Zp?B>�쾽)� ?+߇��%�>@�&?�s1?��>4k?���=hg#�s�E��St<�eM�o�f�c���~���h�<r��=��!>D$�=A�;�n�=��<t��d =���=�}e=��=���=��>b�>�?�MZ?��:��=��D��o��>�Y�>���=���=�@j>ʙ">)+�>��?	�?��R>�Ȣ�y������4�Ծ�۹�GK�>��?A?L%7>�끼٢���K�uL�=��>>u&�)�A�����þ�@���R>JK@>��\>c�?C�z?0��>�EC?v���m���F�
\Q����>B�s���?��0?�B>g����R��E��	j��Wb��긾���+(�<��\>%5=��>{WL=�]���=����_;/ڄ��
彔l=�@�>v��>�+�>�i�=X_���dﾘ��_f ?R�μS$~����nJϾ��/��D#?wj>��K�@{?�sE��V��kcſ�y��x�m�?+�?�͟?�V>vLD��=�$?{�o>5! ��,w=w�]�լ7�s��>L{߽�~���%��[� =��W<;e�>�l+�.'�����TY�Se����Y�Gn�+:��Ͳv��񵾀0��ms;a����H�޾�Ic���c�>zw�lܽ",T��H�O6��~��'S�?)�?�jĽ��r���1�/��r���6>���`o���������Z��X�o�?ž%�	�r02�9u���y��=�T��-h���on�y����(�a��>��E?�
�[e&����2�V�*#>�@> ��s
���-�����+�j?ΰ:?Gr��%�ܾ��y=a"X>��>��>��;��þ<	���>��>�n�>��~W���t�����e��?�G�?8�7?�t��?����(����>�	&?�k�>쟾�@��4�.����>�,0?���>�w�d��������>s�R?E�E�J;>C7�>�/�>�]���A�P;����<Վ���$>"r���^�ږj�!%-��>{�"��>���>u�X�I1���}�>�޾��z���F��{��Ia�M�=R��>��;��:�>0~>M���m�+��[w������5S�|.m?��?_?#%<?���C�����>�僽NTt>ҕ�>�1p�M;��>�!�>վ Jh��NZ���> f�?�� @�<?}Ɂ��ο������p���4�$>9��>s�<>�C8�vyF>�
)=�!L=ܾY�ZCG>y�>�ϒ>�x�>�t;>B�6>��>���CM%�v�������,��8	���	�=LI�������]�a���J����aۮ��{����U�U�/��B�����yc�(i�=���>�i�>� 2?P�>jZ�==���E��/s�T��N���P
����n2'�U�;�4ƽ�����3��Gg���&?��[����>�2�>��&���^>x��=c��=�>�D�>�~n=j1�>�"㼯3�=�Z�=��>�#���=�_=�o��-������Lu�\h�>�>�п����m{<�M���%��,��>��>J
�=x�H���������R�>�g<�����	�]|Ǽ�Y)>ؚ�>x{�=9��:͹�=�"���K��:��x�><�9|���H��3Z�0ߤ=A��>��J}#>b�W>�ZE?r_�?�#?�Z�=*]�>	C>v8$>�2&>J�>�:>��U>P�?�\/?�5)?ԭ�>���=�^���\ >�&�<!������U��0��<##�չ�='p =A�ݼ{��;K��+{�<KK��kQ��ͫ�e=
;?̧I?�%�>/�?H����]��E$�Y�I>Ԫ>/����?ڌ?�y?�H-?�� ?WC=�ࢾ[�	��
��c�>T|�>T��%ڈ�g��;���>1��>��V?�B%?Fk �Zs�o�M>7�6�X�>y}?��!? �>CG�>�h�S��:޿ju���T�\�콫m=>ҡA=\������=f��r�K�n��;Ƈ�>��l>��>�{Q>��>��=]�G>-��>��>��ļ/޻�����|�R�<���<X��^�����������,>�������;�O<P)Ľ��ǽ�����`�>5,?�5A>�ⅽ����u����}��>U�>�z�>j�?�,��uK?����M9�`���=m�>�0S?���>]p0�K��=C�v����Z��>�{>�w�<($">/�	>�aȾ�S]>�J?-6?�vm>�����d��=��� �Gu�>�A]=�%���?3+?�-����'<�M�{�0�����><b;5M�����2�
5��y������iZ�P�����>n(�?V<��T�=�w������7n��̾�.�<�l�=T�3?x��u��r�ɾYN
�\ؾ�k<
��=�K>��+>�W�>�#?�N?E�Z?vw?��>m�_�+?�-��h?�3:?7+=?\�(?s�.?�cF>� >�j�������Jr����<��	�v3�=iep>t>5�[<�&�=��<��G�ǿؼC��=�ʋ=,z!���~;k>	�='��=ǥ?֑1?0U��P8;>�(,��־�`q>�J�>��>l���=>�n�>�E�>�\D?��;?�_�>'>�K3�@�����ھCz缕�?W'1??�>T��=��M?� �r�4�=�Wg>d����G<7���|k�4��!=>��=j�=��B>:�b?R#j?(0?���G���ـ��;���68>������>�Қ>Y��=���+�!��F���6g��J���=v7�u�;<�=�I�>X�=�P�Ѣ>Zh<��n�<A���A�b�L=c?��?v��>({8>0ޜ�J����񾆞X?�&���_��e�=�GE���r=LI?��ھ�5��b?4m�YD��������l�m�>@��?���?T�n?x*�>��}�W�>QQ�>,��>3Z�.�w�BN��?ULA���S�f�P�=mZa>q�?��L����Q�9ߙ<���O�A�Z�>��t�y/���~��\�����e��0e�:I��LҾ��p�Qr��,��@����'���;�۾����׎?��|?p��=�	$��9� (׾�Fm�3�X<u ���t�;��׾�����ž��־�����پ��7�5�>�(���>�D,�̐��׏�d��<:1�<+X>���>��վ�R��E��\�&��U=��=�� �����|G��#�.���d?6<?�̾o�V��{r>���>�i�=���>�վ3�Q=_�>�?x*?V>3����V}��>�?|��?�@?�-B��i@��`� g�Rb?�?��>���˾�8�_m?��:?O��>.������$��P�>��Y?okN�:Y>�-�>�4�>��M%��Ә� ��������@>�|��j �<�\��3�$F�=�>93|>�S��G��N�>���l�b��b1�:�!���P�Q�E>�"?��2��>QE�>k>������dJ�������?�Ͻ?.�b?��`?9����%� ����%���� ?���=:��<P͋�qQ�>��?�(+�) ����<?�M�?f�@�	Y?iW9�"u���������w����w�<W�=t�#>���-�A>�Q�=�$�=�8�<�E!>H��>�[V>pR>��>�>��\>�ӄ�����̣��}��}����X8����Ne�����/�� �{�߾��Ѿ(G�Fn"�x�:=���j/�?I�W���O���!?"��=34�>�����>�}"��e��1�}=t@������)��*s�ſ��E�Mӭ������!���Z�>���:��>��>���ȗ�m��>;*"�$D8>Ӽ>g�6�2%	>�ۄ=N�ټG�r����>H�w>�L��~0<��n�>�o�.�Q������a�;ԋ.?Eɸ�t��`�#��˾3�x=讣>pK�>{0�>��&� �����,��>-�T;ސ"��.G=��>�0>�̔>��}>�����<�<7�=��;K�>��K>��j=�b�=��(�.���S3=��>�ɾ���>Mu�=L�H?��r?�W;?nR�=˙�>�d�=i�>�(��GB>t#�>���>�?�>�'�>�?�G�>�ˬ=�Ľ��>��;>���tJڽ�8ʽX��k�z7$=�rf=%.:@�>Qn�=c��<]�ּ����=bz��?ӐO?)ާ>gO�>+�Ǘھ��w�d։�Z��>7��yߐ>��>>h?類>!)�>�^�X�_��־����Q?���=Nڎ����oA;��O�>��˽l�?I�>?'�q�,%F����=6��>G�>tI?��??�[z>�E�NR�W��K���-Ə��9���Շ<��� �P>S�"��E��O>>�������%��>[>~��;���=E��=7D�= ��<m��>#[m=]7�<]��<z=�� ;�����5	��Խn���'�<Q䷼�Ȁ��۝��g輁@�=��=�*	?%�U?��|=�,Ͻ�־˵
��ƾ!����?�c�>��H?q"�>�2��~�"W���þ�|�>"E�?��5?���l\>R��)�����>���>U"��2��php>�Kn���R=q=5?1S?��>�B}�>�0�<G[����e?��=qݽ|ʛ?�J$?��ξ�ꎾ���m@�nkӾE�x=�2=�|ʾJ���]�N������^2S�C?>���>UF�?�~��6��>��G��D��v�y�V�о��|=��=f5?�O�>>�!�D���Oz1�Jx�f-�=�R�>�ƿ>[K\>���>M,?�sg?��?Ɗ?�@�>!����?ɠ<=��?��?#F?B��>6?��ѽ?�=�׋>f�T�#�����>�<���=�A&>d�=.<�,0��fi=��@>4�>��=��[=���=��g=
�^=�̬= ��=O+J=�'?J*?H����ƽx�P>]�+>�+����>�@>1���b�N��= �>�$�>]?Ѥ�>�"�=`����־У��04ؽ&�?��/?s~?���=��>�;�����j"�=e>NT�=0�����꾶"}�~,�>��>+�k�g�>�8�?��-?�?�)��V����&z�_��>���ϲ?~I-?҇�=�y7�GK��>��/9[�##��U�>FL=�H t���">��>ip>1�v>��=��ּk��X��"E�[���>Ao�>���>-g�=�l��ض��3/���\?��&I���ʾ{)�����=a��<į�>z� �i�	?�G������`[5=x�p?���?T{�?�2?>�4>dT�D�=>B�>7�^�Q>���^E�=)\;>v��>��p��$����刑�Z��>��>�	� J��p'�e1N��ƿ�d���E�M��������
��=�<����=>�<�\䁾|����ԽAH�����Qx˾����?+Ӿ��m?�V?�&�=�%ɽE'!��9� o0�@f =�
��n=��[t�у��K��qm��5���:�
�@%��a0���>��t�����Br�(n#�в��Dl>|2&?�Ծ&���GJ�!��=ZH>C������2����ב���7�U?7�<?pX��|9��_ �&�X=n�?Y[�>�t>Ħ�(��ɚ�>��.?!?������%����p=~�?W��?3J?ۄ��]\�љ�_-�=��>?F?�"�>(hQ��A�����"�?��P?="y>Ry���p���ؾ�d�>s/?�~�4�>��?h�>��r¸���>�ɻ�<e>��>��ս���b&��=j%�JV�=M�>m{>s�S�J���ζ>4���#�՟F��!�:����֨;5/?�O��!�>�>�k�=�A���e�y�h��X�9@:R?cs�?�F?N�X?q}��5���P�q+>�?1�>}�>�'
����>Q �>	e ���n�n�^�?^�?���?��A?6�b�U)߿;󟿞�������={.��f�=�����h->�'0>fS��*���dvk>�ѡ>���>� �>�f�=ȶ�=qS>�����)�����m0��:04��� ��q��K�A�c��Hl�f4��Ĝ�ZЊ���{�̜�#�����
��$���~v��+���28?���>&�=�����7>5^��Z���Y�J�+x+�"���8�X|��z����վ�����q>�Ծn�>���=t�=�4�>�e��^���b�={��=�+�=�u>��<�y�>]�7>"!R>yy�>�y�>:Q�>P^>�-<Y傿��{�o+� �p���}:L�>?�Os��eV�N1�. �N;��Z��>�?EҎ>�$'�5��I�v�Г�>J4ǽ�����*��h�<�|�>`��>�)z=F��=�+ǽD���k|%�e	>��>3�>\���Z���,��m>$��>�ξ1,H=�}>�?6 ~?l)?
�=jg�>u�>�_�>I>C#$>��>9>>Ub?�??�4B?J�>���=�+^��]T<�c=oG��]����ܽĈ��D�K��R<���]=Zy�=�FȻ�@�;��C=CA�<�v����2=���>V�?�y>�t"?Y��;�b7��N������ X����M=6�%>|4>�?q�I?=?��>mΤ�FI8;���>*�>�y_�2Ai�o^�����> o>�%O?>�Z?�N��T�>�k>٥��x>K?$�P?!
f>(x>c4����,�տ�k
�p���S���_ý*=.=�#Aҽ�"U=ё��q⽼��=Yh>\�W>IW>��$>��>�{�=O^�>��i>ۯ�= �=X��Qv'���>)��=�;P�$q��߬�ݸ�<3'q�����T���5ʽ7G�;�U��"u��7?��>�8��J䝾�ƾ�8�������$?�M�>
F�>�O?d/?���\҂��>}��c&���0?�h�?A;�>�gB�
 �>^A�=�L>D��=��H=
'>�C��r��C��`Q�p(�>�D	?�f>E�c��5{�*�w�r!O��?�L=����M�?`J;?���z��S���b�����/N=�Qp�� ��qt��i��8���ھ��ھ75�[�W>�2�>^F�?�ȥ�tI|>�5�!Ĝ�Oⁿ�~���F:�5,*���>�>7�����ꛫ�ݲ=��8�=��ͻ�?�>r_޽�%?��Z?|w�>��?��?a&�G����g?ji�BU ?�֎>��>���=&N�=sM��\�=�E>�J�q��o���Q,=�O��F���R=��0>�j�=��=J�=����u��fF����=j>��>���=`B�=G�m>j��>�|?�+����>x#>�Sf����A��=��>=f�¾>ȯ�>�:�8��2��>~�_?V^;?,�>�J	�.2����ɾH��=�?D\?>-v>��[�>p㽂������>~FS�(E����~��hL�J� ��۾���>}Nk>�f�?!>�P�?�G(?W.?L�=�v��}��~�M(g=g�a�:M�>�<�>�=ShP�8f�fӇ���F��Q*����|f����=�J�>&av=��>)�/>������fG�=g�����#=sĽw��>���>��>�T>:�.=��+�#��W?S6����9�J��kBؾ0=�>' ~>��%?���=1R?�;>~$�]�����$���r>�h�?9��?S΃?�Ǚ��`�=S�����ySa��G�>D�]>�ލ�M�ʽ���>aB�=
�#=����
i>>��|<��O=pVԾ�Li��[q�HGʿ�G��={��A��dJ��:U�.��=�w �ћb>��DT����-��8�<�?o�+�ͽS��������.t�?;�?K��=)!��j�>���
޾`��=0��
ɼ�̾ٓ+��1˾�M���\I�������>�V������>��x����B�BҾg��=^�
? M1?b��,���e��ʾ�r�>�י>H�½s<E�#���n��|�q?Z0?V��np��X�=ǹ$�� 2?@v�>��l�P����߾��[<RV?�|�?s~�= ��kv������:#�?��?8A?m/���LC�����ҿ�pI?��@?�⼽ �ɾ�����l�.?���?$�?\ 6��mw��}+����>�!x?q޾�b?G�?U=7�6>��ɾW�*��t����J��X$>�������ξ[��d�ݽn��<l��=�!i���˾� �>�q侅�5�ի:���'�Z#n�۝̼�?����G>cu>�wB=��+�ۻ���v�ݻ�HL?�H�?��H?DK?R���<�Lr���q����>�Y�>i�_>Y�˽���>���>s��f�v����"�!?��?��?��K?��e��ڿ!ޘ�|��@��z�=W�=+�>�(���,=�=���ļk�>ʒ�>I�d>��>�">>�>��%>�Z���L ��Ơ�����@K�F�.�j��)�L�l�}~R�I�j檾2<ƾ�ڲ��2��vռ�L��WA������;˾�!���� ?�z?Ր>��i��q�>xʾ�O����7�J�wI��4���׬�x�%���.��]��Ӿ � >��쾀�(?�┽a���xR>h��=�=t�>R(>pB>���=>ۼ"/>��>T&s>��>���>� ^>LƐ>
|j��΅���v��E�lWe�A�;�sK?�/t�!��yD7�}.��8��$k�>ɳ.?^��>�6:��"�e�2��>|��_qվ�߻����=ԉ�>�>q}s=��>!_A��dc��m��q�>��>�`>,n��C�Ⱦh���NQH>��>���p��=�~>�_#?_Nk?�(?�"�<�)�>��F>*��>��=�$>v�C>�9�>��?�j9??X1?���>_��=��X���@=�2�=\=�����&ɽ����h�>?=����>E=���<ݍY�	�d=kW=kG� �r;��<�t�>��&?�_�>{��>�ᗾd�0�Mi!�;����2��&���Ј>�S>�L�><��>V?�L�>���>8$/�� }��d�>�!�=jW|���W��;���x>8ԃ>��P?��6?�4l<��<.e�=#63�D�Q>Q�>;uB?0'�>��>��~�$���mӿF
$���!��$��������;V�<��N�F9К-������e�<1�\>�>�p>��D>�>e;3>)[�>�YG>=Ǆ=���=1��;f�;��E��?M=~��OTF<ήP�}S����ż����������I�%�>������ؼ��3?��?H����H��~���L*>|�y��R+?���>±g?:af?*��>�
�?�T�&O���&��"?u��?Y}6?H���=1���L4���W�>��>�G�=�|G����Η��=Й�>�*?���>��s�'p�O[R���#�2П>/������P�?�G?}���&Oľ�o����M�"���ؚ<pM�����wy��ǾU�#�-䜾O�þ�ս	[�=��>��?�`�̚Y=�>��^莿�&��@͘���?�͵�'_�>���=�<?�<ż��b���_�#��=�U�=&V�>p4�>&?U�J?�G�>|�?p�>��>�D�~x?w�ƽ�
?�>0>^�>�m��K�>� �<W(|�wG]=�k��W�s������<�t����h�>�ҏ>��9H�<e��=�4v<Q��Ǣb��AA>�a=x�|=��>$�H>�)�6��>� �>@׻�CZ>$�A�u"0�j炾�W��0^J������"���O=J�=N��>"B>?]��>#(Y>1��o�ξ���5�>�A�>��?Hr�>h)���=�X��ѽBt��;���r��<Ŵ����÷���ܔ���W=^�_>�=8��=�D�?��??�? ��>�{ʾ����w���K�>3�����>:5>j�4;H�=�}�����dׄ���h��p$>��Ӿ0�>D��>���>?�>���M�=G�'��2>xw�ܺ=ʜ��+��>�4Y>�?���>/G6>L���%} ��0?b9���������.�ZA��>ۯ=�E�>ek�����>c��Po�;����|�?�?�E�?�T`?�8�r��=����eq��j��6>���=�鋽iz>>9O�>/f>H�?�,�~���*��>��v>^(�=��޾��e�o;���$ҿFrZ�t��>Mf������O��ܽ/����ݾh�$>F���Ф�����ē=$����fN=�u��k.(�;��<�~?��?�b=���=�� ���ؾ�Ns�6Lg>��X�Q�M=�㱾p�b��_�qdU�>h����t�*EӾ�����׮�>�'ᾍ����`V���,����<vʧ>z�9?q�Y��H
��7.��8�ٹ>^`�>��'/O��d���~B�3uW?�m1?����Q��Ө��t>7$?`]�>�	�=�f7�J1��K��>��~?ko�?F�->[Y���K��5.\���?F��?;�Z?�E��o?`�J�K�yS��F?���>g��>.���7��/��>��?Eg~?t)�>7� �� ��%��w�=��>�����J�>W�>���=�'ؽX� �˔�D����W�*��>�;���>d��W� ��w�$>�f�J#�H��Y��>�,�S�N��H�.g�jm��:�<�?QX���>�Bh>�>KY(�}،�t����� ���L?n|�?BTS?�f8?����S��0��EЍ=���>���>��=���Q�>x1�>%辈�q�Iu�e�?�/�?!��?7Z?lm��ۿB���YS��>�Ӿ��M=��=�'>*� ���=S��=w�:#��=�>�>~�I>ŹZ>3G;>��/>0�>��_&��𛿮���0W��)��9��g�з��� ��@�-"ϾȾ�퉽�z	��ˤ�>�Y�-#-���H����Z+>�!?�<?�2�>u='�#J�>O-���}D�h5�T����2�TL����(4 � ]�}���ި�������=^+�0��>��߽I��=��>��!����Y�<>V��=��>��7>:��=\�G>��=��>E�i>5By>��S>"�>�"�<��y�<�{��<����TKH=�Y?�Uf��A���!�D����ξQum>]�%?��>����Ή���c�6�>!�(�R����i��<@:�>Ht�>Zs>="">�=��+���%����=�DI>�1�= ��<�ǭ��}�O��F�?�j�����m���KH?R��??�bf=�?�ʓ>���>�4=z"��1/=�'`>�1?|!G?.
?a�>BY�<Yt��z�=�Z0�Tf����6�`�5>��K_��(nʽRX�<�h3>6u�=����$$�Oㇽ)��=7�>S�>&��>�F�>��>y�>"���	>���}�'���xɚ��uT�����M�>�t�>l9#?B�D?:�?�\z>:ͽ�Mz�>��>�׽�F�y�B�J������>~��>T��?=*?Y{��������� �S�\��>�x?|$?��;�(J��p�����iӿ��#���!��u��ӈ��;��<��;N���9Z�-�AZ��l��<?�\>c�>8�p>�E>%�>\3>
b�>�SG>B��=���=�;�K;��F�[�N=ʎ��ZJ<Q������ż"x��@���LI�j>��.��׼��?��1?��T�Fb=lXp�J���"���:�?C��>��?(�.?xQ�=�M���m�x�@��{��;?�?�O?Ɓ�,1
?�ɂ�IZ{>���>���	d�&�Ͻ���{{G��y��K�>���>��>�[+��>��P/d���-��@G>k��i�!�?�9_?6[�Ԉ��p_�a�O�@���3�=�����*ʒ�`p���3�)Lþ�9̾p-��V>,V ?�?:�c��$F=Ǡɾ�������y���m�V�M}>N%�>�W> ���z�R��*վQ욾��	��<ix�>+-^�2z,?v?��>>�?��>XL�>���&�9?|�=�p?���=��=ћ=��>a}������ǰ=qҽ)���ӆ�ź�>��@=��<9G�=
�z>���<���<b[켼b��#n�<G:=��=��;��֔=�[�=s9<�^=e��>�(�>�0�(�;���<B�0��޾�������齭�`���־�Q>+��>Q~?.O2?>$?��,>��f��;�=�
�����>3��>�?=�>/?��"��<d�����T��ɘ,�_�H��c���+�0%⽪q^�^�>���>���;��>��?�	?/i$?\\�=z����(d���ʾ�#>�6���>�5>�w��_��W'�^���;�D�y�%�L5Խg2��Z�<��>>*>�=�vs>Λ=~	>���<�/�;H���� �D��2F]>�D�>���>| 8>��̻[�������a?����uH���⾘s�����>�f�=I��>3I�>��/?��>�=b��[��"�#�6?�.�?��?�G.?'`j�kR�̇&>+7�=��[>xb�<s|��NA=&5H��pL=j��=��';Wn�600>��>��<��k��]�Ś���<�ԿA
]�P�>�$v��)��)!�x��l ��辦�>�-�0���J�*? �}؉�^��yc �e!���̡��ߐ?x�,?d���B>�%��x�臾�X_>B��w=�Xk �i���`��Gѕ��kZ���**:��0�\�׾�7�>͡����#x���\�٧:����>g�V?X�Ǿ�e�0�T�j�����>��	?��}���g����E>`�R?E7N?����	r���#��>_T9?��>�<k<o�h=���3��>9�R?l�?�#>/Γ����� _�T�?ɰ�?�[?lX��?s���-?=��?�j[?���>�#��۹���1>�v�?���?�?�$���S��� ��>�q���i�@�?���>s���DW�g�r��@u��ؾ����� ?��a>��c>]����1]����>��H>���XC-�n��>���I���-���u���l��?�?���a�>(rw>��#=b`H�yB��*�m�!��v?#��?�4#?B]?������|%��%v�O&�>�a?K��>ju�=(��>�#?dK��:�N�?<?!&�?��?rRd?��H�Ҿ�U����*��]�0�V=�:�=w��=Π�ǡP=��=X�Z=y� ��7>���>f{Q>��_>:|G>��=��^=!S�����蘿,|��qf�@	)�n��Dd���3�j&����y�Ӿ���|���� ����������F��n*1���
��ȼ��%?&c�>�>�4���v������ �����v���!�h��}�8�ݾ����Z�eش�k���6h>a���!J�>T+b�<] >	~�>j�ý��~>�D><�=
OT>`Lr>]����>d�>wt>��>%0�>�)^>J�>2�/�nя���y��|$�v%N��a="??�3H��/1��:%�q=�����1o�>Y?,?^��>�8 ��]��cv��A�>�w��_�*�^��-�ռ;Ç>=[�>���;�nA=.7���,��,�ɽ�>�x�>���=�}��9��z!��7>3��>�B����|>��>��>�R?��?^����A�>�@�>`|P=����*�=̑W>��`>k=?]�D?l??9 ?!��=hAڽX�=j�,�������;��ȼ�	��C��D��=\��=�H�<��=7�	���L����=��>�)���
�=_�><�?Վ�>�D�>�:���9�ЌO�Qܾʔ������]>��>��?�F2?_�?� �>����߁��E��Q��>-��=�D���a!-���4>j��=�G?��?�r �k䎾�ż�
���ܠ>�?=?'?���>i�G>�ٽ���u	ӿp$#�"S!�.q����"ٸ:�\=�rY��x;�/�!��N�<`d[> Y�>�q>{E>n�>�43>���>�(G>m�=gŞ=n��;�n�;�G�q-_=��5�Z<��H��۬���̼�藽'����F�"�2�&���ݼs�?�*?<Y�=��:�*�Q�(�F��v����>1?�>��>�1?kF�=�U��T��O�l8Z�n�*?;��?�m�>�k�-#�,Gͽ���s�>g�?6��=i��%T������^>L?y 0?P4�>w97�nz���7d���쾏�}>���<}i����?��\?W�k톾�4 �9G���'k)={���e�QX������7�/y���� ��.h�.G�=}�>n��?�
t�q/�=V��񼘿bƄ�߮���H=�gH=���>�-K>�2��u�����Շ̾|hH���<zC�>*b��;O?���>���>�W�?�R?��>�u�=�=?�����R�>4��>Xɖ>���=I�>�d���&�c�m���ɽBS˾Q&�=��=��=�i�=�*$>)Fj=�WU=�9s�����5n���<�=�N�=Q?�=uf>���=,T>���>���>-i뽌�T��Q�<�i�5�E��W���/Y�M�䌖�5��<���>�m*?��"?a��>ai�<Ƿ��v�`���쾌U/>�d�>E�??���>�gؼT|ѽ����XE=V\�M���5����g�7�&}t���=��e>�$�>!�`=��=��?�4?��?�/�=�������D�����>�Fj����>xp�>� <�� �`/�%�m�-N_���I�"<r�Z0k��3>�,>��M=�nJ>�A=��>]�o���=�ܽ�>�Zd>���>pѦ>� �>��d>=�qi����4?0U��U	���.�}U�ʝ��<�>z�k>�jt��EW?� $��-��Wʠ�Ih�j[?Q��?P�?��B?�+s��=�	z;r5t���7�l�>�W���4=5�F�"5>�>����ƾ��"M=r�> �>�j��!R����i#�>ٿ��X���=p��=�P"�wQ%�����������=z��XԾfoe�k�*��L����>�nR��!�ƫ#���8?�b�>�l��	I�<���"T��@�����=Α��ٟ��xվ�J�W;�L���N������Y���������g>�>L�辒뛿�?S�M���!=��>E�?��b�	�0��_�y֤���>A�>��q��X�I����o��V?X�%?�����G5�̏��%ý3�$?���>X�ٽɈ3�ߏ����;�o`?�z?��=%[������O�޽?bǺ?��g??}F��vk��"��P�9�k?*7�>Lh?��>���_�i>��{?�ba?�>������c�S>}ER?K�w�� ?���>8J.>}��=�o��Yc�� ��߿�#�>��[�/�����%�JcM���;ec�>��~������辄�>״Ӿ��`���5�Ѳ�����<�W=S��>�龵^�>���=-�b>Sh�����l/���ye��D?�_�?d�?�)%? ^߾y���ؽ���\�>�1>%�;e���nϓ>���>��վ$������~� ?Cm�?ߟ�?��_?֪h��ο{���J���ަʾj�h=ٯf=ބ=V���N��<4l{���;�ȩ�!>2�>tt>���>���>H�r>�B:>��5T"�����
���M��'��
�/�i���g���I9�og���_žo=k��<H�h�:�M�a�m�ԁ��w��G�ۼ���>d��>_�> T��+>С��f�L�N�@5���5�1{�1�kg���ƾ��6�F#
>�����!(���,?pN�І>i�/>�i	��K�>v��>�e�>�C�>_d>���=6�>��>�ի>�ǌ>��j>^��
�$���X��]Μ��w��ޮ�s�=W7?�񂾙��րR�h��J>�� �>}�?s[K>��4�L��`Pm���>@�G��󒽔�%>�d�=�Wm>8>X>_���'
��������ّ"�ߛ<��(>���<��ټ��\��	x�8��=��>~����>�d�>V�9?�Q?��?ՒT>���>�>�ְ>K�`>,$$>���>�ɷ>��?�k7?k/?�^�>��=�R���=�	=cq��	%�N��n*D;)�н��K�,�0L�=�r�=��=�4�=�u�=���1�q=�.0=�?m�8?ؘ�>#,�>�柽�O��F��n�=#ۑ>M)I��?=��>�ֲ>$?�Q
?���>���=eVy��{޾�س>x�>��@��N��ŽHQ�=_o<>�K?��>?�I��@E�J��<{�=���=Ha?��/?�x�>b��=p{ >k���ؿ���!�j�'�|<����i=���>{���� �v�Z���6�����>>	��>vZB>�!�=" >c>�>�>">>⚭=���=β'>�����ѽ���>���U�A;�K��Q��Q?����(�7����=�=}�?0�:?���^�Y<��^�9����1�$y�>M��>$l�>��>1>p>
tӾ�Mb����dB�f�>�`l?b�?�t���=L�V>������>�>"��>�x.=��-��_¾\0�=̾�>�}?a�@>7!x��b�2���1��	>�t=g^��j�?xzG?������F�^&\�I^�n�=��
�s�ڽ��̾�l"��y3��H�&`��u��M�k��_�>��?�����q�>2u����ߋ��͌뾳Z�=I�
>W�?��>Z���	��I����̾��u�����w�>z�>uR ?�@?�P/?Rm?�>?�L�>�D�>�N@?rv��6�#?�K?2�"?�� ?!?���>T?r>�=g}���
��䤾c��=��<&��=��/>�ج�T��<	A\=)m�=<Լ��&���ʽ�T>�dM<�Hs=��>P>�>��r�?�(?��U��K>&�; bC���'�F�'=d��>�k�<gM	����=D��>'r7?�)�>2�L��.����þ�<�"�>�D#?-k?�I>��`>� ��������=D�Y>Nnٽ������ξ�V��ʕ���$�>\��>I��=:��>��b?<@??eW?h4ϾkM'�)���q27���?��>aT?�ѻ>K��=au̾X��TH�����)x-��Wn��p�� q�=S.ѽ,u�=�2>��=���>m �>�����b��~=H1��`�>|3�>�"?��>��9�!��Rǳ�RF?;���������^C¾�{���
>� B>�׽�	?�[�ssz�Y�����:�W�>^��?R�?��e?��9�J���N>w1f>~9�=M �<w6��}(��ߝ�&�%>��=>Ʉ�%���a�:�R>�Bx>�*Ľ��ʾQi�* i��C������M"i��U�Mˀ��̾�����錭�� �����uV���;���	v��.нn񌾤���B$��aj?%�?bi��
����]�����F� >s���;̾�/�Z���j�-� �R����I>�7d}�Nz�^/�R�6>�Ӊ��`��l%m�����
>2�0?i�>|4�^V����U���&��+�>�kL�t�=�Xp��L���W����j?�K?�㮾����=�=;ͣ>'�?P��>	��k�����=��#>�Fk?=��?N�׼d���h��J��=���?�x�?j=1?$>�QAv���E&\��4?�?�a
>�wϾ�P�-����!?�N?p	e<�=��ꍿ=����?|?�?i�<�
jP>�k�>iӈ>�B`���Ծ�u���->�J>��=����y����	�1>�>Ԓ�>�@+�;�Ǿ���>�U��VN�*H��E�Yj��<(z?�����>\�d>:>r9'�>���鉿2x���J?�A�?T?��6?+���/��/���\�=p��>�i�>�2�=i	�:p�>l��>o��oms�#	�M?�q�?)(�?hZ?\qn��ӿ+-��[�̾�����ֽ�����Q>��d��	><�v>"�<�
���:>�ɘ>���>�`�>��>Hu>��=���*_#�3���U�����d�lM@�����t�8'����<�o�� �?pܾ�}�ص�V*���3 �{s&�s[9=� Ͼ-�G>��>��E>��|>��L>�B>}##�����ɾ2'\���0P���s���ޏ�P�����=��<��	�s@��^�?����?>-4�>�x@<n�>ge�>�pP>k�>w3�>��=� �>E�>D�>5F�>��]>����K�=�~;�k���Z���;����H�O>V]5?����K��T�E�j�"�oN��k6g>3?�>�rc>��.����� b����>99�=*)b�e"x�F���U��>/6�>3����-нǢn�3�c� �:��K>���=*t59���{u;�#R�=;>��?�g߾�I�><�>m�p?:ws?W{?��c>�T?�/�>�>�o>(�w>gz�>'��>�)?�d?��R?�t>��=��ʾ�j>��=#�=��[�ZF��F<��>�޻���;�!=��&=X4>R��=�T>��>֌?>W6*�X
?�#$?���>���>�*��#�234��6>�t�>|��'�>�'�>x��>~WD?��?%J�>�O]�X�վ>��n��>q��>�eh��܂�`�W�WY�k^�=���?��L?�b�&��s@���ÿ<#�>�q&?^
/?��>�w2=����-
�0Fܿ��'�D��aS���½Kwq=4 �ҨX���=��-��p8���<i�A>���>�S�>P�u>�)>�3>��>�L>T;=*L=0B�=ެV=|�=�R=�[��)ȉ����y��o|Ƚ�����ν�J)��I��E:�e�<�?;�?��'��2��� f�M����G��R��>���>�h�>r��>x�=2�
hU�)A��GF�<��>�[h?��>�8�ٽ=[D,��z�:��>'o�>"E>�^d�F��t��F��<c?�>�?�0�>H��@[��|o�M�
�i.�>����"<�`I�?��K?�����׾.;.���`�R�ھ�P/=�2=��/=Oq׾�� ���=���߾���D��m�i�N�>���?X��@�>�8!��܅��Z��^�Ѿ/tf����>�?G��>����-��P.���Cs����N��#�>B�+>�Yl>��?JX9?9r?��$?��>�H3���?�b*>N��>���>��>���>���>Qp>�r�>"G�=������)�x�e�C=�=�{J>
xS>s�>NC=�ɻ�7ؽ&��=
ɽE'<m�� �E�S�Ҽ�9�=��N>`�=��)?ǞO?/F��R7����=�F�l5���>`?� ���������=�nU>&?NK?��$?g,�>�����?�$^þL�s<�>�-?H�?5P�>�>������D[}�A֣>_z�=;f���b;ߦ�wh��}�>Gљ>S�Y>��f>��V?�j?�@A?ٙ���@k�2����`P���ս(�>��?y�?tϾ�?&����B�q�R��S�B-B����T��jŽ�s�=;3>���=�">}Ӓ=�O��n�b<_����|���e>)��>�?���>^�<B�ݾ@Ծ��I?J>��jK�3���D�Ͼ5o�>��=>4����?_��]�}�� ��, =���>b��?���?o(d?$D�]��4\>�U>v�>�]:<�=��~�DK��)d4>˧�=�Qy��啾1��;O�\>fy>sDȽ�Qʾ��㾼bE��`<���.6��,پ��m��䱾�I�o����B_�}��)�n�ܾ$���j�<�>�C��7N|G��j��%�����?�8�?���=<,
��P�_9������$��R�о���ූ����m�� Ӿ����k���d�qe��L�=���;Ȯ��gI��A��|�>��>q��>�2�<�;�^���.�kV�>�bi��m0��ǌ��M��'���_v?5?�����
�2�����&>cB�>��>��I9W|Y�����}>W�V?y
Q?�*��ʐ���T��y<ý���?���?]H?!����#b�T/�l!����>�M?a\>#��D�ܾ����?�||?E9�E\O��W����F�d	�>���?I�}0^>R�>?���>$����ƾH�*������<p��=���=�?p������Î��>�>�Q>���L�cM�>l�z�2Ff�i�\���Q:̽�Z�T�>s��|v<�ٽ�Z=>P!��_��ڇ��u����C?_��?���?�&?��Ӿ����z�V=�|_�d
E>�֫=�H7<u®���>��>��Ծ慿!3(��n/?��?�5�?�1C?� ��,1οl(��Yl̾�&��'�.>��=�>�0��=(�=���= m]=ܑ=�>oM�>=�_>�8�>��i>`lA>�a>�l���s'�Od��A����6�q*���<U�S��fۑ������W���[�������u��+�a�u�i�kg���������	�����>�8�>���><N>Fma>	jP��q��Vޝ��⽑�2��� ��꾑侅�Y���=W�u<�1�� ����3�+�?�G���>F�I>[8�=X@!>r��>I> G�>#�=>�i>��>ǌf>(�>�:�>��b>���:�K >20=�t���}� 47���b���=�R*?~��7[���N4��!��/�Ӏk>�O�>�S3>(-C��5��\�}�r��>���=Vq?��=V�b+�}�>��>��x=K:޼����r־h�e.�=�`L>>�8�A�ҽ�2ƾ�#��L>��>.�ؤ>�f�>�#G?��z?�eG?��=8q?��">T">#�\;�0�>��>e��>8�(?��K?�}0?ck�>8b�=�W��=LL>F�d=K�=��2<^�-��x�R���>9m=ٿ3<]��=)E9=F�n<�a=�wA=}�׼Y>�����;]�
?E�0?(Q�>��>�޶���+�.m"��!>��>������>	�?l]/?�9?._�>��>��d={`�}j����>�:>JT��Kv�.�:��a�;{��>��?OW?˵��U�-���M>FQ/>X�>�?�g,?��?N��>(/`<�����п�]?�%��lF=���2o�.����þ��=���>�ҽl����>� �>@ �>�0*>W���l=N�>'N6>�=�X>)��=�د=���<o��<�\#���U=� f���齏-���2��. =�=V�u(�Ph��A��%?��?:��c�4�/V�����ɾ�Ԫ>���>P��>���>�o�=_M��f��+F�i�r����>*Hl?�??[_�A2�=On=�]=�>�v�>�>��������#���]�=�8�>�?�^�>���	J�kDm������>}ؑ=�rB�¨?��d?d�Ⱦ���@�A�R�T��e��>V�>�~U��pýk���l,O�Ø1�i��ъ��~~'��{�<�Z�>
��?��:�>�D�/R��vM���&F�[䵽��>}��>�=w>�5}�\W����L�-�d���Ѧ��޼H>�)�>�>kw�>I/?:;R? �J?Z�?}>ɳ4?�Ɯ=��S>cM�>�)?�)?k�?�Z�>�>:�=�V½����������`���Y>H{>�8>-�s�!Y�(�L����=���L�/l�=�H�<4Q�X�m=��>��">�j)?�y7?�c���<6�p=�<��.> ?RE�>�ky���C��>r�?_Y ?v�5?0e?h�[>�PB���Bk����)�? 7?���>�h>7Z
>O'������!G>�#7>%�u���p�����9��1����=�у=Zc�=�{�>5Av?]?D�?����[�����(�ż��Q�>�JB>>8�='�0�A��'2�������n�����U�9�5�/�\= �Ͻ߄ ��{>�`[>I�>�+���-G<C�ž&h��?�w���F>�P?\�?'�>�7�Fα��p޾�yI?�L���>;��о�$�B�>�;>ӷ�"?�W�V}�Zʥ���=�I�>t�?���?2�d?¦A�f8��'\>MZ>��>a�;<O�@��=�.ֈ���4>�Z�=-@x�R=���zV;�J]>1�y>��ȽD;˾S��ydQ������e�ᑾ����r#�%���pmn�i�~��6��zȽ����Ҿ���� gὫ$�=����Π����2<Ͼu��?E
�?��T>N`��w0�K��tF��?�>��:�Z�^���eѾ;���ཾ���UE �XN�&�A�A���e>'�<j���E�����%�DdP=�c�>��>kO�Eg����]�e���X8�=9,㼹s:���������>[��I�?S�>?�J����.��i>T(�>��>T'>�*���f�4>ʽj?�j�?soE��������2_>���?Jw�?y�6?ٽe$M�o�p�����>��?lz�>e����޾� s�9X?��<?���> �b����f��'?^Gz?�B�>�7>3�>�ȡ>~�����:�n씾�$P;�'>�e�<��v┾D���~>*��>�2�>J2�G:��">Vh�����_� ����-��X=���>hy������=K����E��~����q��
�½��9?t��?c�?�s$?'�ľo����m>�0�:�V���6>���=O�j�;��>)�?�5[�d���������>'�?�)@�nl?f^��$g��,�����A��P���Z�=�8�=lT>����-�=�ϛ=xwF=T}���J=��a>��B>��j>�>>��.>��\=�m���M&��������P�
�=�d��>5�����MӾc/�v��������@�B�����»���S�B����������>^�J>	j���>��>��>}:���c:�k�pg.�Ū$� �ɾ�ξ�VZ��x�<2is�Hմ��r�����t?8܎�2�>�<q>Xu�=�B�>�?3? x�;$�j����>���=1��>f?h�>(n+=�D�=�g�4x]>�U=@���+|��I:���V�ݹ�<�wL?�:3��0���05�cᾁ����(�>��?bvT>�@�b퐿��v����>�ڇ��:�C���a׼�wf>f��>~?�=��=}`�f�n��$��%��=s�>��+>1sK<X�����ʖk=/?9�����>���>�?v��?�3?�̰��e4=��>z�$?t>�>�>�>\>��?�O?2?.X�>?�>t.L>��
��!M<�p=U��9
��xv�[+n�N����އ���4�l�&��Y=��z�_s=J1�=nO�f�?��)t= �>�T:?��O>|�>�a�i�$�a�9������r=�B�=�t�>P�>���>��'?��
?Q�>|�%�ե��V�3�>@�f>��;��ad���n����=�h�>(8e?�?x���h,���ǖ>o��="�z>y@?�l]?*!?�D)>*�����lӿJ$���!�w����N�2	�;��<��M�*՞��-��������<��\>��>M�p>+E>�>+;3>�R�>�FG>�҄=q�= -�;o�;��E�_�M=��wYG<��P��]��� Ƽ�9��:�I�j�>�>1��Cټ)��>YF?n��A���ʾ���z�����>�v>
.�>��>��<:��>�\��V��I���? �q?
��>��j�=w�=��5>�+�U��>]x�><>r�<ɡ��.\ξ|�\�`-�>q\!?�8�>Ƚsh�*���� 1���f>a>�'�ٽ�y�?�H"?��-��)|���.�\�H���Vu,>"E��*Q�mꌾ5�<��?B���������ý�z=���>b��?�;��䱜>ښ�*�v�qҙ������}=B�L>�H�>L=�Q��/���"�w�1������S%��K�>|S�>��>xV�>TZ?��`?h�,?���>�s,��t�>���>���>�
?�[?�0?�?s�>���>�����b�E����o��.>�=����?>�3?>5_���<-<�71>��<��!��Q��?�=�<׽�*�Fp��O=7˟=^�?]�5?9O^��c˽9,�=̹���g�>f�?>��x�\�=�Xv>�؊>���>$�a?��?z�=�Mþ"�쾚¾�0[=K��>�>7?�w?)�>��7>[��-�b�4w��G9>�T1>-�H� �󾄨پ4A�N	~>���>�E>I�`>)u�?9�?'O?�X����o��촿i�8�7%o>띱>f�6>��@=�r����پ�d4�I���/҄��.��ƴ��֌���j=��½��!>���>L�@<~�'>�>E����A�|�n=��P���>�X?�\?d�b>K��=����о�(?������'��N���q�3,<��X&>2��=d����+�>����7y���/fV���N>���?<��? j�?��7�,��pc>�v�>���=b���2��\=����V;)> >�"V�ɐ���I=S��>�l4>�
7��	ؾ�������輿�I��*Y3=�'��\��kZ�����(� >n�<�U�� a(��Ed�ޑž�䏽\X������䥾�����qȾ��l?��y? W'�'U��E�;z��˾f*�R�X/�@Ѥ�2	A�Ls�<7��)���2�T8�a��r����;c�/JL�pU��r���ǚ�uצ=�ؾ>���>�ﾪ�s�A�Q����D>M7��*�����7����L�GX�?x??f�G���Pn&���>�F?6!<>"��=�x@�n<�=J�a>��$?FP?hV��ӏ��Y���&=q��?N<�?�:?��@��:@�qc�����%?�D�>#��>P�f�{O���Ž�~�>'�1?6�>�����ㄿL!����>rMQ?�FA��P>Y��>p>j>n�C�+��[V*<6쉾�cƽ6�,>z��=Sޅ�[=^��~-����=���>�lq>ꢈ��FžcM�>l�z�2Ff�i�\���Q:̽�Z�T�>s��|v<�ٽ�Z=>P!��_��ڇ��u����C?_��?���?�&?��Ӿ����z�V=�|_�d
E>�֫=�H7<u®���>��>��Ծ慿!3(��n/?��?�5�?�1C?� ��,1οl(��Yl̾�&��'�.>��=�>�0��=(�=���= m]=ܑ=�>oM�>=�_>�8�>��i>`lA>�a>�l���s'�Od��A����6�q*���<U�S��fۑ������W���[�������u��+�a�u�i�kg���������	�����>�8�>���><N>Fma>	jP��q��Vޝ��⽑�2��� ��꾑侅�Y���=W�u<�1�� ����3�+�?�G���>F�I>[8�=X@!>r��>I> G�>#�=>�i>��>ǌf>(�>�:�>��b>���:�K >20=�t���}� 47���b���=�R*?~��7[���N4��!��/�Ӏk>�O�>�S3>(-C��5��\�}�r��>���=Vq?��=V�b+�}�>��>��x=K:޼����r־h�e.�=�`L>>�8�A�ҽ�2ƾ�#��L>��>.�ؤ>�f�>�#G?��z?�eG?��=8q?��">T">#�\;�0�>��>e��>8�(?��K?�}0?ck�>8b�=�W��=LL>F�d=K�=��2<^�-��x�R���>9m=ٿ3<]��=)E9=F�n<�a=�wA=}�׼Y>�����;]�
?E�0?(Q�>��>�޶���+�.m"��!>��>������>	�?l]/?�9?._�>��>��d={`�}j����>�:>JT��Kv�.�:��a�;{��>��?OW?˵��U�-���M>FQ/>X�>�?�g,?��?N��>(/`<�����п�]?�%��lF=���2o�.����þ��=���>�ҽl����>� �>@ �>�0*>W���l=N�>'N6>�=�X>)��=�د=���<o��<�\#���U=� f���齏-���2��. =�=V�u(�Ph��A��%?��?:��c�4�/V�����ɾ�Ԫ>���>P��>���>�o�=_M��f��+F�i�r����>*Hl?�??[_�A2�=On=�]=�>�v�>�>��������#���]�=�8�>�?�^�>���	J�kDm������>}ؑ=�rB�¨?��d?d�Ⱦ���@�A�R�T��e��>V�>�~U��pýk���l,O�Ø1�i��ъ��~~'��{�<�Z�>
��?��:�>�D�/R��vM���&F�[䵽��>}��>�=w>�5}�\W����L�-�d���Ѧ��޼H>�)�>�>kw�>I/?:;R? �J?Z�?}>ɳ4?�Ɯ=��S>cM�>�)?�)?k�?�Z�>�>:�=�V½����������`���Y>H{>�8>-�s�!Y�(�L����=���L�/l�=�H�<4Q�X�m=��>��">�j)?�y7?�c���<6�p=�<��.> ?RE�>�ky���C��>r�?_Y ?v�5?0e?h�[>�PB���Bk����)�? 7?���>�h>7Z
>O'������!G>�#7>%�u���p�����9��1����=�у=Zc�=�{�>5Av?]?D�?����[�����(�ż��Q�>�JB>>8�='�0�A��'2�������n�����U�9�5�/�\= �Ͻ߄ ��{>�`[>I�>�+���-G<C�ž&h��?�w���F>�P?\�?'�>�7�Fα��p޾�yI?�L���>;��о�$�B�>�;>ӷ�"?�W�V}�Zʥ���=�I�>t�?���?2�d?¦A�f8��'\>MZ>��>a�;<O�@��=�.ֈ���4>�Z�=-@x�R=���zV;�J]>1�y>��ȽD;˾S��ydQ������e�ᑾ����r#�%���pmn�i�~��6��zȽ����Ҿ���� gὫ$�=����Π����2<Ͼu��?E
�?��T>N`��w0�K��tF��?�>��:�Z�^���eѾ;���ཾ���UE �XN�&�A�A���e>'�<j���E�����%�DdP=�c�>��>kO�Eg����]�e���X8�=9,㼹s:���������>[��I�?S�>?�J����.��i>T(�>��>T'>�*���f�4>ʽj?�j�?soE��������2_>���?Jw�?y�6?ٽe$M�o�p�����>��?lz�>e����޾� s�9X?��<?���> �b����f��'?^Gz?�B�>�7>3�>�ȡ>~�����:�n씾�$P;�'>�e�<��v┾D���~>*��>�2�>J2�G:����>G��>�O�!�H�(�W���@[<�R?��|>�b>NR>��&�����M��Y���XM?EI�?gZR?C8?������1��[��=Qo�>�e�>���=�J��ՠ>t�>G�O�q�U��s�?�H�?wE�?�dZ?V�m�!�Ϳ����&�
���־�a�=�ݖ>��]>������=�f��t�\=��=�>��>in�>ky�>�Ǒ>��T>�7B>�L��CA��3ÿ�2��>�U�W*�j ���F�Pܾ1KF�'�"�	窾|������2���Lq=�����(��I��y�� >|��>k�>gg5>{���[7(>J䈾��ʾ�bԾf�����^	���^+�:Y��$�S��I�FG�M���_پ��>���=�NL>��?{�>Rޱ�$�>D+v=��d>r�b>Pe�>�`>e�>p�>�dd>8�>�U�=�K>��E>b3��jI���9��
�<��<��\?�R���:������� �qs;�M>;v?Z�">�z/�W,��i
���?�;�|����+�=9�5���>F��>�S�>h��w���ʽ2�^�!t��#�'>���=����>�� �����>���>��۾�
X>�w�>sQ?~tc?9fO?>��t�>�#�>�C~>褝=)��>.�>@�>�?T
<?o�.?�!?�T">C�;��=7>�����-=e��=!��;��o��\�=,㱽�q�=j�=TR��T]�=2���X߽���=�?nEj?��?��>l�E�i1���o�D�r��'�>n/��%�?<7?�+?��?2�?ގ>�W�=/���]�`ȫ>d��>UU�� ���{%=�?e/�<-�?%�O?ȋ�=�$w�=�->T��=@��>�g�>�H?L$8?���>%p��MԿ��k���E���=�O�H�\�(�
>*�>哢>�SվĲ<	]N>=�<VU�>$�?)*�>�f�>�5�>�"�>�?�=PY>���=��>��W����I�>���<�|�>�Ι���=׵�=7-�6:��9��^;�������rN?�9?�4n��#@���Y������+ة>*I�>!
�>���>�o�=�T���X��
K��ky����>`Cg?AM�>�!�b��=Siq�Mc_�^%�>�|�>C�$>���w4�gP��\e�<uB�>>�?Xƣ>� ��QR�@�k�����>zG >��ҽ,�?��h?]�j�[�d������a�eB7�T�>V:#<9���f����nW��:�I�.�x�	��,��B>|J�>�R�?̠�}=����Go�� �� ����=P|���?:�>�U�$��^��Z�3c��MM>�0=T�o>�;�>uk/?��'?+�Z?[�?���>�B���G�>�o�C�?J��>� �>z1?��?rE�>�>�+:>7<�$���}>�P-���=h��=�3=$jV>���<��1��=�OH>j�g[�<�-�<ZƤ�u��=���<"�H>'�?38?])S�_��W�1� a~��Fl�8/>=���>�M���U��'>ߐ>H�?�\'?,U�>H�I>p������
yZ==�	?LR.?�*�>���=�,>��	�+�X��>�\>��K?]�u���8n��T۽���>�Q�>�Zb>u�?�I?��2?]$%?�m}�b=��ng�I_3��zӼ��8���?Ok�>�����~���g��?f�~㴾S|>�f½j����=���=WƯ=��:�'�=�Va>��=Q/V�4���$m�=���>�|�>��?���>���=����i���I?8���Lj�m�qо=G��>��<>����?8��M�}��
��kG=����>"��?r��?�?d?��C��)��\>NV>?�>�8/<f�>�'������3>o�=|y����T�;�]>SHy>�ɽ��ʾ2侒xH��	��P�L���������wռ > �>�����	>�g5�ȣ�>Q����
�!��:]�8��������I����_�?Eݚ?���=.l��VdY���鎾�C=�l��n�&���ྊ2ľ)����D�a���kB��`�� !����>8N���Y���~�QtP�Q �=���>��p?���������u�9�B���)=�����݅�*����,���gJ?�%?�߾K�E�ƽ�=�����)>!T�>�'�=k�ھ�F�����>?��)?�Y�=IY��Ք��*=�K�?���?��8?��'�D3�.�=%��%ǟ>�� ?X�?����þr�;�(��>"?7o�>����$���� �Ax�>oe?�{t��	>?�R�>1ޛ�ȷ�O@M����[��<���>/)ػ3�c��v����>��[C>)��>@��7٤�F*S>��;4�<G�a7L������e:��
?ƭ1�l�w�	c=���0��o���Tj��%ྺ&?�x�?@�t?���>�|��]���)�=gZ.>��>���>?�L�ǂ_>+�2=9�>�ؾ��z�(lh�:�L?��?kR�?�)?�b���ȿ*���(��[�ܣm>�*C=�l��Ž�	<���>$�J���='��>�b�=�Ї>�>L��>���=�F>�ن��(�ۖ��Ľ��4ξ����g+�Y�$|�g�̻	,e��.�C-b�C�G�Ar�������������@<���h�;�V?^��>(ve��%����=v�k��Q�t9�,��Ƨ?����)��(�ž&?վ��;���]��g
���6�yv?��F>.9�>D?n��>%x�>��>o2�>�>�%�>4��>���=���>5)?��=��M>��>0�x>�[�=�������>;�BVS�ix�;�t@?�`�h����(4�W�������>,?iL>�3&��C��� t�H�>� �_c^��j���}�4�>���>��=Y�<:v
M���r�^�ս��=祊>��>9Ϲ�,k�������n=G�>
j9������>�R�>�^E?f�?��=�?��Ͻ>�P�>z��=k��>1��>�{?��G?1K?o�?	>>�Z�Py5����=�p�<�G�̨v����<��<�=YeW���	>�4Q=�SB���;q�F=�V�=C�V=���=�[�>y� ?��>��z>_!��nf��A�	���5��=���j~�>y~!?Ϸ�>�~#?�.�>���>D3�=�����[[�>u��>�s���D�(�=�V��[ ��&?�+?B`[�u����>�<M=�>*A�>-�?�
?��>������|'ӿ,�$��n!�JM��ӏ�d�;%W<�"�A��i��̋+�9G���Y�<�B\>���>�wq>��E>�!><4>G"�>��F>�!�=��=d��;�KM;c3F���E=�n� �O<��Q��Q��5tʼ	���2���eI�eHA�Z���ԼP7:?��`?ڒ���/+����H8־",����>�Z�>��?_L?u>�۾U �����HʽU��>*1_?�:?GýF��=vC�<�>H*�>�J�>7ɷ=���N*#��t6� �>n�>�~(?�>��,�F�u��_���߾6ܴ=*=���ㅾ���?/uA?�G�p������h}�'~$��H�=0��1�B��}Z�^9c��~�<��X~0�wX�yI\=��>��?�h�1�?��7�9ߴ��#ä�����rU>eu���>��9> ��ʋ���U(��
%�J��r��������{�>ď�>em�>�K?��;?0w?�o�>l�=�?1��={��>n��>��?Q�.?���>�>�>��>�&�=}���bJ���� ,>	(���b�=��>��>%�3;Š��!��:Cj�������n���	���*<.GM�u��O�<���=�i?1�?�B���<�+j<��*����<�:�=+φ>����Ͻ^?>�$6>��?�0?,?�z>>��K�OṾ��꾲o�=LA?a /?C��>�;�=-UM>з�xZ8��c:��bj>m�6�7s\�W����Ň���;�e�$>u�>��=yν:tq?8S?7��>m�|�wPl�v���@1��g��ڼx�%>M�>����
�h��q���k��X��/�Ӄ�=�Y���ϴ>��4=	1>��>�ڶ>ґ����ͼRB�4�z<��>�M ?�K?lL�>�KQ>�Xx�R?��I?���9~�IZ���Ͼ�SD�� >n;>���"�?@4����z�y���x9�+��>I_�?6H�?��c?N�6���彉�k>Q�J>� >V�O<��;�p7�Ww�S@=>���=͕t�~���W-<��Y>�Hp>$6ͽ�˾]�߾nPS��Nȿ߸���"��t���#Ⱦ�Ο����=�ϥ�+�J>�-b�rԽ �0����Z{1=_4�Pcr�mZ��{���?+��?c�>�˾G��#��e̾��>���Ӟv�6� �5̴����^���(��
��D�c�����p3������O��!=ʿY�s�v��7Í����?���Zt���ͅ��`x����;�g���c�j���%(ſ5ͼ���]?c99?*���y�I-B>'�C�p�>���>*䋽ʋ$�=���@�?�>/?�l�%�������V�Lk�?Xn�?U`4?��8��AE�~[�P݂�(j?��?p��> ���;b;ѽz��>�@?���>A��Hy����Q��>�an?n�@�S->;2�>�%�>R
�!,������C�K%=�d>�V�;6sĻ�7M�_�l�j#�=���>�4�>_W��>�߾1��>FﾀGU�{�M�m��V$���Q<�?��!4>+J>��>Ʋ"�� ��������uqM?<�?��T?;m6?������ni�����=�!�>�>�5>ƽ�"�>��>�Uܾ�d�:>��?�8�?�m�?�Y?��q�;Hؿ5���_�վ߾G-�=�~>��*>Ԫ�֖�=;�<=Ǧ�<떽5��:k)L>�1;>BW�>V�%>N�x>��u>������b�����?2�U�	�xQ�e��L����(��*羾p�&1?��j�;C���G���	����<i�����c>�{�>C>�%?;�q>qV{>�9K���f���儽���þ��"��;n������l�e�#in��:]kS�����X�><�>�$�=���>&����i3=!��>S��>�)�>� >=�<�-��:N�>#.�>�j�=�Me>�Ƚo�|>L)�>�:���휿�?"�2f(>��<�'m?�㳾���<�G}���"���ݽ��I=��?@�->P�0��t���M���L?��<����?I<�f0���>�{�>��>�)���O��þ���K�>��=��ͻ�M����B�iѮ�Y����W ?ߺǾڽ���>v|*?��A?Ϙy?�L>�f?��Z<i�>�T?�����b�>y}�>��Z?uz?�]t?�h#?T�="���������$��E����<i<��=Ct`<��=D<G��x4=R��=;
�xU<��b=�����༷:F<�!?s6�>2}?��!?����O�>�n�5����m�=�'*�'*?�q-?Y�?��1?���>�>�M^�|���5,���>��"=M #�dUV�@�ٽ_�>x��<�`4?��-?�m9�<zs��x�m�=kg�>.�>O?D��>��q>&.�a���wO��˧Y�(rW�m��}�eE���<���>J�3>T.ľɥ徸�w�&=��l>�i�<�g�>t� >�1�>U��>��>UD>��;3>ς�����:V�,>�ݑ��>��N(Ӽ��<4� �m2�=� N���<�����ɖ<�?�??w#����{Qg�n��LϪ����>G`�>���>���>ع�=6���U��<A���E��S�>]�g?˧�>��7��A�=)#)��?�j#�>���>r7>0 j�t)����_��<���>>�?@��>]f�B�Z� �o���
�NQ�>�{�=�5K����?�{?�����I�g��Y�c���6��	>e�����}�o�O^��D��+���+���q�%�\>��>���?�g��>��1���������ܾܣ�<�E9�_s�>]�>�@d�-����V�p���Z���r����:<5�>�'0>0��>J�!?ǟL?bq3?[��>La�:Ma�>24��?�v�>!?%�0?��?�G?�
?n��>c�n���7���7�7[ӽ� �dE>�3>�I�>P<*B]=�)������(�� �H��u��1��RK=���=�S>�{>�="?���>��=��=��d���ǽ,�_��~=��_>.����0=���=��>]�4?�L$?�$�>Ys�=�G�����5� �]f�=r�>:?�
?�E>�8>����#���x�=���>��V�SB߽�QҾԩ��[X�*��>q��>�Ml>���>��?�1j?��?Dƾq8x�l�|��`��Yx�z7���ɡ>k#�o�����3t�4x���i���i��������)��-Y=��1>��%>�fU>�E>�3�;'���LJ���_>��=��R>��)?�W!?���>_>>Y���b�þ��I?��k��ߠ�gо 1�c�>��<>���l�?�����}�����8=�)��>���?��?�Ed?��C��� �\>�MV>��>,�-<t�>�J��~��h�3>�@�=~y�E���8�;�]>�By>j�ɽ�ʾ{D侜�H��"��v�2�u|�������2�̛o�^�r���>Y��@C~>Y��ꃾc�{��K�p��=	W���(��@��M۠���?���?$4�����PT�'{�S:Ҿ2�>g��D��j��y$��t��	���3z1������^�.��g)�,��>�pD<���	����F��O>�A/>|ӄ?�5��(��l_��������>��¾|�K����D��T�W�])?!
?#��xn�=E>�����9�<B{�>��z;��Ҿ&��r ?��\?m�(? k���ͭ�ո��I�=��?r��?��;?Q>��,����~��Mo�>��	?�m�>��ҾK���U&.��t?T�D?q�O>!�1�o⑿|&�T>�>�Mn?�ꂾ��z>�?^F�>F˽f¾�d=a ����j�>{$j=��W�������F�=�,�>V��>-=����u��a�>��$jN�^H�>x�ζ�3��<��?������>�i>R>��(�("���Љ�I��gK?��?o�S?k7?R��zZ�L��߰�=�>�)�>�4�=�՟>r��>���1�q���D?t��?�z�?�WY?�6m��ֿ.ћ��ᵾmB��ō7>{�>>��=6z���;2m�=	��p
F��	G�H��>�>�-M>~��>'�R>�@>�����"��������� - �*��cq�٭M��i�Pb���,����5�������a�{(����ҽ �0=�ߚ���<R�>( �>֠�=)�#>�Ŏ>��I�7��,þm󩽤;��.�Rv����!�J Ծ.�¾�Q���ڻ�W�E��:��>̤E>,>>ű�=�-N=���>	�>~��=�"�<��>{��=f�>dX�>�h�>\h8>���=��e>�T�<�}�~e��#eY�Dݵ;�����o?�y+���Ͼ�
[������G%ؽQ� ?Q8q>�>�Mߧ��A��|�?3�>�]�/~~��🼘�>�= ?��>V�������1%����G��>�B>(��/��M���+> ]?�ճ���P��w�>�;A?TU�?��u?��>�J�>]<�I�?ݯ?�½h>C�>E�D?�C?�u?��>*u�=`&\�W�t�_�+=�jH�N��3�_<㐪<{����=����\=�*;�8�b��=�E�=��F�
ā�ҳg=>�?W I?^�?
q!?R�e%Y��Q���[=�N�>���>���>�n2?��>�8?�̺>AW�=���9�
��2�>�B>�8�N��$��=�q?rH�W�P?��Y?����X[���>1W<�wg>�1�>\�'?���>�Y�>�\>�	��Կ�P�Ē8�f�>�D�=a$���-��)C�>�;.>I� ��"���\>|�>�ö>�v�>���>�M�>�)�>^U?�\>�Rb�2%(��k�>RG=i����=8J>.1>�jپ..=�s�>-�s�ĉ��>U���Ƹs����<
N?�?�$�������d�%���{骾�s�>��>�m�>�`�>���=�L��AU��r@�j�D����>7�h?O��>�=9�?w�=� -�A�:���>�ǡ>�H>g�g�?���z��f�<Ѽ�>9!?�Σ>�,�q�Z�r�n���	�%�>���<y1�AD�?ddo?<��Ѿ ��"�Z�V�%����=*�彄PW�`!�jN�H����^=���:����>��>�y�?s,�;o�� |_��d���������ZD<��o��G�>��>�־���P4E��Z��X�|�ڈE�u9>��>(K?D<	?0MC?�N)?݆�>Z3n�5+?����?���>��>�;?���>��>��>�>C2>��@F��W��;�@�<=�u= �(>UP>ŽA��;ɖ�����u�1��<i9N=���<��<H�n=��^>�p>�s?119?w�r=��=�L�<[Q��6Լ�@>��U>ʵM=Q�ͽ\���L�>��>�D?%��>#�>{aɾY�a�۾4u�{$?g�M?T��>/.���}�>mݳ�q�쾵
>�3o>=V�W����v������`���j�>fv�>^�> �o>�F�?�k?/�>��s�X�a�%ᒿo�F7�UJ>�}�>���=��G>���pQ8�����M@��'�wÚ������k�=���<��>67/>�X>��4>��=�)�=g�->�@<�{�.�>�V�>�V�>ݢ�>\g>%�����?J?�9�����sF��q�;0���>�s=>kw��?y���w{��E��A�<�^,�>N�?SK�?Ke?3�A���R�[>OW>�>�Q�;8�C�����j"4>~��=M
z���_'�;�vb>�1{>5�ɽ��̾�⾋7���Pm�F�����&�k)���2#��Zž֦�=�̻=�,��<��Ш�@�=w��GW��ˢ�)�ϽK�˾bFӾEć?LPw?�u�>��1�����3��4��ul>Q����"���ڽ~��������ܾ㏉�a�!�r66�w�j���Y�q��>��p��<���$K�MP��6�>Z�r?b�� ����h(��<��L~;��Cu���������7,F�809?h?A�׾^X��i>Ƞ< �9>ے�>(_���4��������>AV-?�?|���Ф������5=�ʾ?���?́6?1B�G�5�T	��B��v�>;Y?��>��߾�"�ƽ��?b�?*�6>S(�Y^��S�7��]�>5�l?�!���>g�?�/�>·a���t�������rά;��g>�s>#��Ɵ��(G�z��=^a�>S�>�|z�ݓ����>��J�M���F����dY(���Z<L�?C���b>n`>�>�"(��莿ՠ��c���EF?[Z�?�W?�A3?����R��f����=��>���>1�e=���ş�>���>�?���u� ���Z�?���?���?�U?�o���Ϳ����̉��zQ�����=�:�=>
E>��Q����=2W�<��}=;B��=�v�>O��>Mx>r�>�q>߬8>����'�U���+�����3��%��#���D�@�������_��"����BѾn�����!���[l�������z�oCI���=hC�>Ί�>��b=�D>� >�n��� ��h{*�0�ؾ־	��������L�������+�L�?��jP�4�A�I��5��>gz=�DL>�0�>�:S<�4�=E�?�F>�O=am�=p��>F�,>5o->D� ?6��>�D>T��Е�=±:>�Ђ�"虿9���c�u�<��D?ۣ?��,�<��0��*�����g0>��?��=������g����>��= �������>�?��>�9q>SA��*��������2�o>!Y�=o��='�H<?��?�ݾ��@=��>X��J\>�
�>��>�tc?�s?<��=N��=^��z�"?�'�=#6w����>}�?��E?"�C?eX?�>�I�;�4�h��܃������Ee><_�;OZ�<Q��=LK=�ؽ�bp��=4����=5j=�˺=x>�,=$��>�BH?�M1?��?¹��a�=�j�4�t�O��C�>��=���>��?��M?u�??7�> �>�\�=�ʾ�K�.�>,�	>���z�w�c���W �>��?)K3?�0�>Y6��K��^H�Y�����>9~?( 3?Br�>kX>4�c>lJ���ݿO?R��::�u�=	�Y���S=���=ڸ����]=����me� +����>��?H�~>��>�v�>���>���>/+H>)$>H��m�c=ڔL���W��F�=�&�<���>I����4�=���=�]���B�"��=�N=��2��Ľ1�?h�?cQ'�ɕ�� r�+� ��i��o�>���>��>V1�>�>�=�����R��6>��W����>l	c?_�>��9�*��=��0�g<׶�>g��>��->2lb����蠾x!�;�>d?��>{�����U��l�]�	���>�G>���?�:w?��
�ɸ��;� lI�v�\�d>jO��o����r�=r^�OFZ�;�2�ѾQx���Sa>M��>��?�:~;�">�{~��뀿J5����� �"�">��0>�:�=�Z�Պ�u����� ľB����=��[>�m>�
 ?�7?�7?A"?��0?���h�><ӽ�E?���>1C>�1?p�>���>�k�>�"�> W��+J��f���NϽٸK��A)=f<�=Mj>��.�w9��ف<_�d=)�=	R��Շ�o8�=}L���-��=v�=:�=Iv?��.?�=���=x��=�e���Ѽ���=�?�>m���Խ�M��@o>r�?��?;%�>Y��=����S򾫱�����>ǻ??�u?�]f;�~�=D�P�k���+��q��>\c:��ԾNA������$�8���>o)�>;��=�~>T��?�YO?��?��>�2@�sM��)�S��>'g��w��״�=@��>T���Mo���f��B'��1w����	m3���>[��=�X=��=n��:-�>��=�K�=nb(���>?̧=�F{>I�?�k�>ẵ>՘�=�+���Ǿ	�I?�󡾳������Ҿ]��p>�=>�����?�z�fC{�����H�;�lO�>�d�?-��?��e?�k?��B���Y>,�Y>{>T\<8�,���o���7>5��='d���疾���;e�W>��w>j�˽B�Ǿ���[�7�l�����,�ƌ���-�>��x�9��N �=�j����>����@��Վ����󟼽�����˽t�a��ꩾ�B�?]��?)�� P��}�:�%�¾����˽��G�(h��D�2��Ҁ����Dо&a�x���(��t�s��>j 	=�
��t}���)<��e�>w&�=�Fh?����P���F��G�����>@��F�ک��>Ϳ
"˾�_[?"]/?=F�a��?�>�'=8�:>(uN>`'�>�ݾ%ێ�a�>�>�?�� ?�l�?��������/����?��?�C?ˑA�7S9�=�j��
��>���>n ?�&�������M�V�2?��?���9������G�wD�>��?���4h�;{+?v�?�q%�0x辭�f�:0�?�=s�u��+g="��q%��=�WP>X�>3�>��w�OH���>״Ӿ��`���5�Ѳ�����<�W=S��>�龵^�>���=-�b>Sh�����l/���ye��D?�_�?d�?�)%? ^߾y���ؽ���\�>�1>%�;e���nϓ>���>��վ$������~� ?Cm�?ߟ�?��_?֪h��ο{���J���ަʾj�h=ٯf=ބ=V���N��<4l{���;�ȩ�!>2�>tt>���>���>H�r>�B:>��5T"�����
���M��'��
�/�i���g���I9�og���_žo=k��<H�h�:�M�a�m�ԁ��w��G�ۼ���>d��>_�> T��+>С��f�L�N�@5���5�1{�1�kg���ƾ��6�F#
>�����!(���,?pN�І>i�/>�i	��K�>v��>�e�>�C�>_d>���=6�>��>�ի>�ǌ>��j>^��
�$���X��]Μ��w��ޮ�s�=W7?�񂾙��րR�h��J>�� �>}�?s[K>��4�L��`Pm���>@�G��󒽔�%>�d�=�Wm>8>X>_���'
��������ّ"�ߛ<��(>���<��ټ��\��	x�8��=��>~����>�d�>V�9?�Q?��?ՒT>���>�>�ְ>K�`>,$$>���>�ɷ>��?�k7?k/?�^�>��=�R���=�	=cq��	%�N��n*D;)�н��K�,�0L�=�r�=��=�4�=�u�=���1�q=�.0=�?m�8?ؘ�>#,�>�柽�O��F��n�=#ۑ>M)I��?=��>�ֲ>$?�Q
?���>���=eVy��{޾�س>x�>��@��N��ŽHQ�=_o<>�K?��>?�I��@E�J��<{�=���=Ha?��/?�x�>b��=p{ >k���ؿ���!�j�'�|<����i=���>{���� �v�Z���6�����>>	��>vZB>�!�=" >c>�>�>">>⚭=���=β'>�����ѽ���>���U�A;�K��Q��Q?����(�7����=�=}�?0�:?���^�Y<��^�9����1�$y�>M��>$l�>��>1>p>
tӾ�Mb����dB�f�>�`l?b�?�t���=L�V>������>�>"��>�x.=��-��_¾\0�=̾�>�}?a�@>7!x��b�2���1��	>�t=g^��j�?xzG?������F�^&\�I^�n�=��
�s�ڽ��̾�l"��y3��H�&`��u��M�k��_�>��?�����q�>2u����ߋ��͌뾳Z�=I�
>W�?��>Z���	��I����̾��u�����w�>z�>uR ?�@?�P/?Rm?�>?�L�>�D�>�N@?rv��6�#?�K?2�"?�� ?!?���>T?r>�=g}���
��䤾c��=��<&��=��/>�ج�T��<	A\=)m�=<Լ��&���ʽ�T>�dM<�Hs=��>P>�>��r�?�(?��U��K>&�; bC���'�F�'=d��>�k�<gM	����=D��>'r7?�)�>2�L��.����þ�<�"�>�D#?-k?�I>��`>� ��������=D�Y>Nnٽ������ξ�V��ʕ���$�>\��>I��=:��>��b?<@??eW?h4ϾkM'�)���q27���?��>aT?�ѻ>K��=au̾X��TH�����)x-��Wn��p�� q�=S.ѽ,u�=�2>��=���>m �>�����b��~=H1��`�>|3�>�"?��>��9�!��Rǳ�RF?;���������^C¾�{���
>� B>�׽�	?�[�ssz�Y�����:�W�>^��?R�?��e?��9�J���N>w1f>~9�=M �<w6��}(��ߝ�&�%>��=>Ʉ�%���a�:�R>�Bx>�*Ľ��ʾQi�* i��C������M"i��U�Mˀ��̾�����錭�� �����uV���;���	v��.нn񌾤���B$��aj?%�?bi��
����]�����F� >s���;̾�/�Z���j�-� �R����I>�7d}�Nz�^/�R�6>�Ӊ��`��l%m�����
>2�0?i�>|4�^V����U���&��+�>�kL�t�=�Xp��L���W����j?�K?�㮾����=�=;ͣ>'�?P��>	��k�����=��#>�Fk?=��?N�׼d���h��J��=���?�x�?j=1?$>�QAv���E&\��4?�?�a
>�wϾ�P�-����!?�N?p	e<�=��ꍿ=����?|?�?i�<�
jP>�k�>iӈ>�B`���Ծ�u���->�J>��=����y����	�1>�>Ԓ�>�@+�;�Ǿ��>״Ӿ��`���5�Ѳ�����<�W=S��>�龵^�>���=-�b>Sh�����l/���ye��D?�_�?d�?�)%? ^߾y���ؽ���\�>�1>%�;e���nϓ>���>��վ$������~� ?Cm�?ߟ�?��_?֪h��ο{���J���ަʾj�h=ٯf=ބ=V���N��<4l{���;�ȩ�!>2�>tt>���>���>H�r>�B:>��5T"�����
���M��'��
�/�i���g���I9�og���_žo=k��<H�h�:�M�a�m�ԁ��w��G�ۼ���>d��>_�> T��+>С��f�L�N�@5���5�1{�1�kg���ƾ��6�F#
>�����!(���,?pN�І>i�/>�i	��K�>v��>�e�>�C�>_d>���=6�>��>�ի>�ǌ>��j>^��
�$���X��]Μ��w��ޮ�s�=W7?�񂾙��րR�h��J>�� �>}�?s[K>��4�L��`Pm���>@�G��󒽔�%>�d�=�Wm>8>X>_���'
��������ّ"�ߛ<��(>���<��ټ��\��	x�8��=��>~����>�d�>V�9?�Q?��?ՒT>���>�>�ְ>K�`>,$$>���>�ɷ>��?�k7?k/?�^�>��=�R���=�	=cq��	%�N��n*D;)�н��K�,�0L�=�r�=��=�4�=�u�=���1�q=�.0=�?m�8?ؘ�>#,�>�柽�O��F��n�=#ۑ>M)I��?=��>�ֲ>$?�Q
?���>���=eVy��{޾�س>x�>��@��N��ŽHQ�=_o<>�K?��>?�I��@E�J��<{�=���=Ha?��/?�x�>b��=p{ >k���ؿ���!�j�'�|<����i=���>{���� �v�Z���6�����>>	��>vZB>�!�=" >c>�>�>">>⚭=���=β'>�����ѽ���>���U�A;�K��Q��Q?����(�7����=�=}�?0�:?���^�Y<��^�9����1�$y�>M��>$l�>��>1>p>
tӾ�Mb����dB�f�>�`l?b�?�t���=L�V>������>�>"��>�x.=��-��_¾\0�=̾�>�}?a�@>7!x��b�2���1��	>�t=g^��j�?xzG?������F�^&\�I^�n�=��
�s�ڽ��̾�l"��y3��H�&`��u��M�k��_�>��?�����q�>2u����ߋ��͌뾳Z�=I�
>W�?��>Z���	��I����̾��u�����w�>z�>uR ?�@?�P/?Rm?�>?�L�>�D�>�N@?rv��6�#?�K?2�"?�� ?!?���>T?r>�=g}���
��䤾c��=��<&��=��/>�ج�T��<	A\=)m�=<Լ��&���ʽ�T>�dM<�Hs=��>P>�>��r�?�(?��U��K>&�; bC���'�F�'=d��>�k�<gM	����=D��>'r7?�)�>2�L��.����þ�<�"�>�D#?-k?�I>��`>� ��������=D�Y>Nnٽ������ξ�V��ʕ���$�>\��>I��=:��>��b?<@??eW?h4ϾkM'�)���q27���?��>aT?�ѻ>K��=au̾X��TH�����)x-��Wn��p�� q�=S.ѽ,u�=�2>��=���>m �>�����b��~=H1��`�>|3�>�"?��>��9�!��Rǳ�RF?;���������^C¾�{���
>� B>�׽�	?�[�ssz�Y�����:�W�>^��?R�?��e?��9�J���N>w1f>~9�=M �<w6��}(��ߝ�&�%>��=>Ʉ�%���a�:�R>�Bx>�*Ľ��ʾQi�* i��C������M"i��U�Mˀ��̾�����錭�� �����uV���;���	v��.нn񌾤���B$��aj?%�?bi��
����]�����F� >s���;̾�/�Z���j�-� �R����I>�7d}�Nz�^/�R�6>�Ӊ��`��l%m�����
>2�0?i�>|4�^V����U���&��+�>�kL�t�=�Xp��L���W����j?�K?�㮾����=�=;ͣ>'�?P��>	��k�����=��#>�Fk?=��?N�׼d���h��J��=���?�x�?j=1?$>�QAv���E&\��4?�?�a
>�wϾ�P�-����!?�N?p	e<�=��ꍿ=����?|?�?i�<�
jP>�k�>iӈ>�B`���Ծ�u���->�J>��=����y����	�1>�>Ԓ�>�@+�;�Ǿ���>�U��VN�*H��E�Yj��<(z?�����>\�d>:>r9'�>���鉿2x���J?�A�?T?��6?+���/��/���\�=p��>�i�>�2�=i	�:p�>l��>o��oms�#	�M?�q�?)(�?hZ?\qn��ӿ+-��[�̾�����ֽ�����Q>��d��	><�v>"�<�
���:>�ɘ>���>�`�>��>Hu>��=���*_#�3���U�����d�lM@�����t�8'����<�o�� �?pܾ�}�ص�V*���3 �{s&�s[9=� Ͼ-�G>��>��E>��|>��L>�B>}##�����ɾ2'\���0P���s���ޏ�P�����=��<��	�s@��^�?����?>-4�>�x@<n�>ge�>�pP>k�>w3�>��=� �>E�>D�>5F�>��]>����K�=�~;�k���Z���;����H�O>V]5?����K��T�E�j�"�oN��k6g>3?�>�rc>��.����� b����>99�=*)b�e"x�F���U��>/6�>3����-нǢn�3�c� �:��K>���=*t59���{u;�#R�=;>��?�g߾�I�><�>m�p?:ws?W{?��c>�T?�/�>�>�o>(�w>gz�>'��>�)?�d?��R?�t>��=��ʾ�j>��=#�=��[�ZF��F<��>�޻���;�!=��&=X4>R��=�T>��>֌?>W6*�X
?�#$?���>���>�*��#�234��6>�t�>|��'�>�'�>x��>~WD?��?%J�>�O]�X�վ>��n��>q��>�eh��܂�`�W�WY�k^�=���?��L?�b�&��s@���ÿ<#�>�q&?^
/?��>�w2=����-
�0Fܿ��'�D��aS���½Kwq=4 �ҨX���=��-��p8���<i�A>���>�S�>P�u>�)>�3>��>�L>T;=*L=0B�=ެV=|�=�R=�[��)ȉ����y��o|Ƚ�����ν�J)��I��E:�e�<�?;�?��'��2��� f�M����G��R��>���>�h�>r��>x�=2�
hU�)A��GF�<��>�[h?��>�8�ٽ=[D,��z�:��>'o�>"E>�^d�F��t��F��<c?�>�?�0�>H��@[��|o�M�
�i.�>����"<�`I�?��K?�����׾.;.���`�R�ھ�P/=�2=��/=Oq׾�� ���=���߾���D��m�i�N�>���?X��@�>�8!��܅��Z��^�Ѿ/tf����>�?G��>����-��P.���Cs����N��#�>B�+>�Yl>��?JX9?9r?��$?��>�H3���?�b*>N��>���>��>���>���>Qp>�r�>"G�=������)�x�e�C=�=�{J>
xS>s�>NC=�ɻ�7ؽ&��=
ɽE'<m�� �E�S�Ҽ�9�=��N>`�=��)?ǞO?/F��R7����=�F�l5���>`?� ���������=�nU>&?NK?��$?g,�>�����?�$^þL�s<�>�-?H�?5P�>�>������D[}�A֣>_z�=;f���b;ߦ�wh��}�>Gљ>S�Y>��f>��V?�j?�@A?ٙ���@k�2����`P���ս(�>��?y�?tϾ�?&����B�q�R��S�B-B����T��jŽ�s�=;3>���=�">}Ӓ=�O��n�b<_����|���e>)��>�?���>^�<B�ݾ@Ծ��I?J>��jK�3���D�Ͼ5o�>��=>4����?_��]�}�� ��, =���>b��?���?o(d?$D�]��4\>�U>v�>�]:<�=��~�DK��)d4>˧�=�Qy��啾1��;O�\>fy>sDȽ�Qʾ��㾼bE��`<���.6��,پ��m��䱾�I�o����B_�}��)�n�ܾ$���j�<�>�C��7N|G��j��%�����?�8�?���=<,
��P�_9������$��R�о���ූ����m�� Ӿ����k���d�qe��L�=���;Ȯ��gI��A��|�>��>q��>�2�<�;�^���.�kV�>�bi��m0��ǌ��M��'���_v?5?�����
�2�����&>cB�>��>��I9W|Y�����}>W�V?y
Q?�*��ʐ���T��y<ý���?���?]H?!����#b�T/�l!����>�M?a\>#��D�ܾ����?�||?E9�E\O��W����F�d	�>���?I�}0^>R�>?���>$����ƾH�*������<p��=���=�?p������Î��>�>�Q>���L�cM�>l�z�2Ff�i�\���Q:̽�Z�T�>s��|v<�ٽ�Z=>P!��_��ڇ��u����C?_��?���?�&?��Ӿ����z�V=�|_�d
E>�֫=�H7<u®���>��>��Ծ慿!3(��n/?��?�5�?�1C?� ��,1οl(��Yl̾�&��'�.>��=�>�0��=(�=���= m]=ܑ=�>oM�>=�_>�8�>��i>`lA>�a>�l���s'�Od��A����6�q*���<U�S��fۑ������W���[�������u��+�a�u�i�kg���������	�����>�8�>���><N>Fma>	jP��q��Vޝ��⽑�2��� ��꾑侅�Y���=W�u<�1�� ����3�+�?�G���>F�I>[8�=X@!>r��>I> G�>#�=>�i>��>ǌf>(�>�:�>��b>���:�K >20=�t���}� 47���b���=�R*?~��7[���N4��!��/�Ӏk>�O�>�S3>(-C��5��\�}�r��>���=Vq?��=V�b+�}�>��>��x=K:޼����r־h�e.�=�`L>>�8�A�ҽ�2ƾ�#��L>��>.�ؤ>�f�>�#G?��z?�eG?��=8q?��">T">#�\;�0�>��>e��>8�(?��K?�}0?ck�>8b�=�W��=LL>F�d=K�=��2<^�-��x�R���>9m=ٿ3<]��=)E9=F�n<�a=�wA=}�׼Y>�����;]�
?E�0?(Q�>��>�޶���+�.m"��!>��>������>	�?l]/?�9?._�>��>��d={`�}j����>�:>JT��Kv�.�:��a�;{��>��?OW?˵��U�-���M>FQ/>X�>�?�g,?��?N��>(/`<�����п�]?�%��lF=���2o�.����þ��=���>�ҽl����>� �>@ �>�0*>W���l=N�>'N6>�=�X>)��=�د=���<o��<�\#���U=� f���齏-���2��. =�=V�u(�Ph��A��%?��?:��c�4�/V�����ɾ�Ԫ>���>P��>���>�o�=_M��f��+F�i�r����>*Hl?�??[_�A2�=On=�]=�>�v�>�>��������#���]�=�8�>�?�^�>���	J�kDm������>}ؑ=�rB�¨?��d?d�Ⱦ���@�A�R�T��e��>V�>�~U��pýk���l,O�Ø1�i��ъ��~~'��{�<�Z�>
��?��:�>�D�/R��vM���&F�[䵽��>}��>�=w>�5}�\W����L�-�d���Ѧ��޼H>�)�>�>kw�>I/?:;R? �J?Z�?}>ɳ4?�Ɯ=��S>cM�>�)?�)?k�?�Z�>�>:�=�V½����������`���Y>H{>�8>-�s�!Y�(�L����=���L�/l�=�H�<4Q�X�m=��>��">�j)?�y7?�c���<6�p=�<��.> ?RE�>�ky���C��>r�?_Y ?v�5?0e?h�[>�PB���Bk����)�? 7?���>�h>7Z
>O'������!G>�#7>%�u���p�����9��1����=�у=Zc�=�{�>5Av?]?D�?����[�����(�ż��Q�>�JB>>8�='�0�A��'2�������n�����U�9�5�/�\= �Ͻ߄ ��{>�`[>I�>�+���-G<C�ž&h��?�w���F>�P?\�?'�>�7�Fα��p޾�yI?�L���>;��о�$�B�>�;>ӷ�"?�W�V}�Zʥ���=�I�>t�?���?2�d?¦A�f8��'\>MZ>��>a�;<O�@��=�.ֈ���4>�Z�=-@x�R=���zV;�J]>1�y>��ȽD;˾S��ydQ������e�ᑾ����r#�%���pmn�i�~��6��zȽ����Ҿ���� gὫ$�=����Π����2<Ͼu��?E
�?��T>N`��w0�K��tF��?�>��:�Z�^���eѾ;���ཾ���UE �XN�&�A�A���e>'�<j���E�����%�DdP=�c�>��>kO�Eg����]�e���X8�=9,㼹s:���������>[��I�?S�>?�J����.��i>T(�>��>T'>�*���f�4>ʽj?�j�?soE��������2_>���?Jw�?y�6?ٽe$M�o�p�����>��?lz�>e����޾� s�9X?��<?���> �b����f��'?^Gz?�B�>�7>3�>�ȡ>~�����:�n씾�$P;�'>�e�<��v┾D���~>*��>�2�>J2�G:�����>�U��VN�*H��E�Yj��<(z?�����>\�d>:>r9'�>���鉿2x���J?�A�?T?��6?+���/��/���\�=p��>�i�>�2�=i	�:p�>l��>o��oms�#	�M?�q�?)(�?hZ?\qn��ӿ+-��[�̾�����ֽ�����Q>��d��	><�v>"�<�
���:>�ɘ>���>�`�>��>Hu>��=���*_#�3���U�����d�lM@�����t�8'����<�o�� �?pܾ�}�ص�V*���3 �{s&�s[9=� Ͼ-�G>��>��E>��|>��L>�B>}##�����ɾ2'\���0P���s���ޏ�P�����=��<��	�s@��^�?����?>-4�>�x@<n�>ge�>�pP>k�>w3�>��=� �>E�>D�>5F�>��]>����K�=�~;�k���Z���;����H�O>V]5?����K��T�E�j�"�oN��k6g>3?�>�rc>��.����� b����>99�=*)b�e"x�F���U��>/6�>3����-нǢn�3�c� �:��K>���=*t59���{u;�#R�=;>��?�g߾�I�><�>m�p?:ws?W{?��c>�T?�/�>�>�o>(�w>gz�>'��>�)?�d?��R?�t>��=��ʾ�j>��=#�=��[�ZF��F<��>�޻���;�!=��&=X4>R��=�T>��>֌?>W6*�X
?�#$?���>���>�*��#�234��6>�t�>|��'�>�'�>x��>~WD?��?%J�>�O]�X�վ>��n��>q��>�eh��܂�`�W�WY�k^�=���?��L?�b�&��s@���ÿ<#�>�q&?^
/?��>�w2=����-
�0Fܿ��'�D��aS���½Kwq=4 �ҨX���=��-��p8���<i�A>���>�S�>P�u>�)>�3>��>�L>T;=*L=0B�=ެV=|�=�R=�[��)ȉ����y��o|Ƚ�����ν�J)��I��E:�e�<�?;�?��'��2��� f�M����G��R��>���>�h�>r��>x�=2�
hU�)A��GF�<��>�[h?��>�8�ٽ=[D,��z�:��>'o�>"E>�^d�F��t��F��<c?�>�?�0�>H��@[��|o�M�
�i.�>����"<�`I�?��K?�����׾.;.���`�R�ھ�P/=�2=��/=Oq׾�� ���=���߾���D��m�i�N�>���?X��@�>�8!��܅��Z��^�Ѿ/tf����>�?G��>����-��P.���Cs����N��#�>B�+>�Yl>��?JX9?9r?��$?��>�H3���?�b*>N��>���>��>���>���>Qp>�r�>"G�=������)�x�e�C=�=�{J>
xS>s�>NC=�ɻ�7ؽ&��=
ɽE'<m�� �E�S�Ҽ�9�=��N>`�=��)?ǞO?/F��R7����=�F�l5���>`?� ���������=�nU>&?NK?��$?g,�>�����?�$^þL�s<�>�-?H�?5P�>�>������D[}�A֣>_z�=;f���b;ߦ�wh��}�>Gљ>S�Y>��f>��V?�j?�@A?ٙ���@k�2����`P���ս(�>��?y�?tϾ�?&����B�q�R��S�B-B����T��jŽ�s�=;3>���=�">}Ӓ=�O��n�b<_����|���e>)��>�?���>^�<B�ݾ@Ծ��I?J>��jK�3���D�Ͼ5o�>��=>4����?_��]�}�� ��, =���>b��?���?o(d?$D�]��4\>�U>v�>�]:<�=��~�DK��)d4>˧�=�Qy��啾1��;O�\>fy>sDȽ�Qʾ��㾼bE��`<���.6��,پ��m��䱾�I�o����B_�}��)�n�ܾ$���j�<�>�C��7N|G��j��%�����?�8�?���=<,
��P�_9������$��R�о���ූ����m�� Ӿ����k���d�qe��L�=���;Ȯ��gI��A��|�>��>q��>�2�<�;�^���.�kV�>�bi��m0��ǌ��M��'���_v?5?�����
�2�����&>cB�>��>��I9W|Y�����}>W�V?y
Q?�*��ʐ���T��y<ý���?���?]H?!����#b�T/�l!����>�M?a\>#��D�ܾ����?�||?E9�E\O��W����F�d	�>���?I�}0^>R�>?���>$����ƾH�*������<p��=���=�?p������Î��>�>�Q>���L�x�H?�l�z�������[��X>��Q�"?����T�:�@>~�[����^�h�"Ğ��MK?��?O��?� ?蛽�	����>@�C�$�>I��>�7���2Ǿ�^�=� ?oR�ԣZ�N�F�k?Y��?R��?t?�����Fӿ�
�����������=$�=�>>�޽�ȭ=�K=���}V=���>ڏ�>�o>a;x>��T>�<>j�.>9���3�#�gʤ�Nْ�?\B�� �����ug��{	��y�_���ȴ��� �������Γ�_�G����hT>�h����5~�&�=DO�>?~4R>_`�>�{	��"ʾ�E��'½�����U4ھQ��s�=���>L�9���v���"�I�:���&?�<9� �@��S�>���=%m>��>G�v��3�=�{�>/�=�C>��>�Z�>Ϫy��0%>/6J>o�t�8�:��{�o7������[ȾQ(k��_5?[z�>"精�Ԅ�;:T���+�>9��>�^F>$�2�o�j��,��z5�>�R��a�e>>�� >���>��>�?~�h�/>�C�=*a��@ɼ�2>@K�=T�>r2���FX�OE�=ٲ�;Z�>*c��S>�G*>q�>5c?J?m9,>�7=>_ڛ�Zc�>݇�=�L>Ri>>�х>�X?��)?n�?]g?ď�=��+��!>&�齲�����#�Aq�9ڃ��=�;��a�;����#��]<�<�>���=M�>�����<�x?|�d?���>�5>:-��M|�@�K��0#>><g�	��>'\4?z1Y?��?��%?��>Ŕ��J�p2����>%�a>����2��N���{�=�<>�}?�{m?��������>� ?���>z�W?+�m?���>���=�������տ����<4����;��<�!��W��b�P� �I�P����'ؼ��Q>ꏒ>HZ�>�3>^>��)>
@�>�13>R��=�Rb=��:=���=B��� V��F���r#=G!/�f���B���:������@���~�5 ���D�=�a?�?{-�X����.����ƾ�ꍾ�;�>�Q>��?�h�>�/������b�O�c��DW�7W?HJ`?	�>�=˾*�<�9ʼ٘=�l?��>�{Z>@²<_6x��A����3>��>+?��?N�Q���t�Nԍ��&�"��>f�����μW��?�6?I�Ծׇ�f ���1�F1��*�����=�d���ݾ��8�:�b&������}��K =y&�>�?�i���=�(�����������A��=ª�>��=�\>PS<��f��$*�Y�5����e�N����=ۇ�<�ā�0?*F?��"?�^?�o]?�@��V>��>헒>
�n>�P?��3?�K?kկ>l�'>�yt����>��,�\���֑�4eY�I��<�E�=�>%=�n�:Ƒ�9Be3=R��<<~�<��k=q�X�Kc^���<�'=Y/>%�/>�?��e?� �G�e�~�Ǿe��r=��(??h:2=�I-��<�=��?�D&?N�x?0�!?4w�;���*��������B�Q?6�[?��?ڢv>Ɖ>��,��i�Z���Bz$>������ �.�?
�"Y˾�ux>)��>d��='�=΅?�j?^P?U����x?���S�<~w�����iN_>X��>�o>�&�����a�������m��c]��}ǽw �����$�7=*>�2.>�m��Y**>��>!�>�?+��[��L��a�>���>/�?�h�>d��=�5���7ƾ�!a?�j���>�jM�<��C=㪆=E�=�׈�A��>�ٗ�{8��Xw���6���'>I�?+>�?a��?�r�zҾ���>{�>�q={CK>�����Vd>r��L}�=#��>ĳE�����p&>A_�>�"P�֜��7o���:�łܽ-�ɿ�"g�̳���\8�>4Ǽ{�������� =l�[�'l<��!��~������<�g���菉����ǽ�6 �?o �?��A�<���%�Ǻ�B��(Փ>M��Մ�0���+��LѾ^bþ4!�����9���8�9����>�g�����㍿�q	�H��=����K)(?4�u�j���N��t*>�>u;��H,����-ל�3�d?c�|?m㣾&�S�Z����=>7?b��= ��>#ι��&�%'?cW?V�?��%���4&��.�=���?��?F�??�R���@�������&6?5�?��>�)���Oξ���u�
?�G9?�M�>���䄿���+��>��[?؉N�Kc>���>�J�>���{��[�*�]N�������`:>�������,�i���=���=���>u�v>��]�����J?�(�i�v��̾+H.�rq��.�K�?�k��,>Ƚ>��r��Y��C8��{����)����>�{�?��|?4�>�I��\�Xl��N�:�N��^�>h{x�:����t>���>Q�,����q�7��1�>6��?���?�8?	��n+ο�Y��!ܮ��L��:��=秱=�a@>���ϛ=a"�<���;��V�>Z��>�RQ>T:�>}Â>c&L>��/>UH����$�Pܨ�8���C(;�)����~�v�����e���%�m���s�Ҿզɽ}O��Kk@�S3S��17�+=	����)<m�B>���>�s�>��>��>{i��G����n+��6�\W�����{B��
��+|�r|A=l����k2�Y^�&=?���<�H�>�?�U��"&>��>��;b��>�X>`��>Y��>ʰi>5bj>���=��1>h>p��> �?>�؁�r���B���#��u>�1�?$�J��[��;��������;� �>�<?��>�#0������J��E�>��ǽ	Q��B�̾��=��>�ϥ>��=��<�=�H����,��B>Fܽ>;�g��Z0���x�W�=�$>~��>����̚>x!�>�1N?�q�?F�^?�����3>��>�6�>�1�<�W(�w��>��>ԩ/?}�c?b�+?{? ��=��=��">��]�`,;��E��i�������g�'�<x��.=Kf�>�p�=�/	>!N�=�<�p<�|n��&?q�??��>��?��۾�q���q�k��2I>�3���y�>�?R-?%�>lA!?�˱>{�g�H���7���>�>Zӂ�5�d��Z���Lz>o��>"�y?q�C?��U�(�y��2�>��t>< �>��7?0�*?"4>3�">)�<�������{d����=������G	�kBb>L?���Zؾs�(z�=�D�>�5>�Ǿ>*u�>�>'g�==v�>%��=s�����=��>�&���>2��B:<�'\>����.=W�=��5�k/�=XnȽ�~����������?C�?�{����Ǽ�?�����y�f�>jZ>s��>$��>[�׽]/�;Lw��C��|b��Q�>�5x?�M�>���} �=h���h���?��>^Os>X����S�eš�<�����>!E?���>�K��#C���I���:�[+b>@eK�L��a��?�|9?
ϡ����*�iEZ��T8����BO�h�Ҿ+�����;���s��0��L��սg=tT�>Tt�?���,ٱ<���[��yZt�5��5�yܶ=�f�>[g�=罾����:��B(��������c;�=�u=9�=�;7?��+?��?zd?��P?����>G4�>��>K�>�>܇,?S��>��?C
?!�˽�h(>U�1�dݯ�<�A�<��>���>��)>_=�O �D{�=v�=�����[��YX��DC�AuU��w�<\m�>��>�{?V2?��<���=�m�`ө�i3Q=*	9<��> 6������	��>�<�>}?�{?=K�>���<J�s�"����g+;�%;?��0?63�>)�#�0\�>Y����엾���;�4>�=��H��퍾�5����I�&�>9��=k= >Y#>���?R�W?J�3>���fe6���~��PL�a֒���>OmC?�~N>*X�ٮ徦L�o�l������4���W�}�ݽ֗}����<�33>%��=�>�;RG>>RQ=y�(>sK���É��.<Ġ�>{�?��?���>�f>nʫ��5�TZI?�O�����b#������	�����>ù>��1���>F��}�������HY��;�>�8�?G'�?�6w?b(�ڰa���>��n>���=�Ĩ=_R�P��<�cֽ5,>�ta=!���}��{ƽ�y>Az�>����M����4��f�w�ÿAT�����'�*�p�8�! ��	Ӿ��0=Y$>o�X�8���b�﹆��b�;· =\U���/U�2����g���d�?p�?%�|���):A��پ�� ����>�v9���=�%W:y&��U���Tξ|g��n�C�Hg�SSҹ>̓���A���_���/(�>pV)�9�r?W��Ⱦ�r ���_>;�Y>
������3��򦞿N��Hjg?@Ti?��<r'��[>Li=͙?k�U>�W>����%<ʣ?: ?wJI?Њ�����[�� x�����?���?ҧa?� �P�\�pr��{X��?K�>QV&?C'��ʾ�b8���?D�j?ܯ�>J�پS�~��� ��4?ב:?Δl��'�=��>C�>������9g�^�پ�g��es>�m<�'� ����`���޸�B�>R�>�~K����;�>�#��9q�_�����tp3��佽��>�վ9U�>�>�Z�;	�	�⍿f�N)Q�׊(?q`�?�Ai?ǵ$?�2��f�-���hp�E�>���>�P>� ���n>���>��	 ~�X40��\?���?CN�?�{e?p�O��Ʒ����bH��+���H�>�w�=9�_>��:��>ʽ>YC.�����ӑD=	��>.��> k�>1��>�<'>ܖ>U���ȋ��֬��'���w3��3��:?�Lӽ��پL�p���&��֚��]��֑�tB7��䯼����;`�ц�6Q־-��<�ߚ>�Ǆ>�?��>>���>��������;��R4�{E&�W�s�� �n(���>c`��.�#��j���M�>�<�<�O<�y�>Y �=�Z�<Ҏ3>��=��>|�p=:�0>�v�>�'R>]>�=��>�v7>��;���=I�X�_�"����#�~t�����XG?��.��@k�ICM����N��/w�>0?�Ԧ>��U7���x��w
?2-
��þ��ƽm��[�>�ޡ>��!>�弽�'/�k0Z��o����R>�ʎ>�>[�&�\�ԾN�����=��><K���=]�4>� ?м�?�^1?ӪQ�I܊>R��=��v>N��+�>��>���>�?�4?x2?�/�>K9
>�rS��A�>Z�o=�h��L�ݻ�b��[
"� �E=�ݽ��ͼ��<�BG>}�)�[��=�ڿ=�-W��V�k�\���>I�5?�_ ?�-%?��޾p6�V&׾;����;>0��=#/�>.�>Ϥ�>	?��>0�g> 4�<��־�Q��#�>��>�P�)m��y��2�>�.u>�Xs?=�J?�k�=:/���'=��>���>>�?��9?�r�>~e>�1=}��!�ʿ-�&�EG&����=	� |#<�&��m����2=[�]��D�S���i>o�k>S�K>Hf�>,+>�Kj>V��>�Z�=w��=��=7�Ⱥ)~�=;�5�������߻�9�x|����1=�8������t�r�n;C�@6�<����`��iA?"$?��@��e�L��b��緾Y?��0?��I>w�?��>_歾(�h��sE��1���>9�U?7D%?t�v��Y
>셸=��J>3?	 #>2��>E�%�/Ӿ�t�����?�>�]�>lS�>cD:�o�FpN���%�8�*>��ּ9���ۍ?m�W?�� ���#�J޾|�3��K��4���wỞY���U��f�Ծ=v)�����J�������ս_�?nݯ?-}���7�=C��r���zz�<7�@V"=q{�>
(-?���>%H���Ӿ9+)�L�CRn���<٢�>i>��>L)-?�n.?�}N?�m?p>?����� ?���>Q��>���>��?	&?�8?98?��>*F�O�Ͻ��������K=��м�d�>��~>��~=�7>o�>y��=P�=�᜽�2E��~=��=ڹ<w:q�=>c>Ͼ?
�-?Nּth�=r�=�㏾�>�
>�>��z�;<��/&6>u�#>\�>?���>�+�=�C��
�������D=�D/?&�?���>K<J<�k>�:(��4Ҿ�=i}�>TI�BÓ�bH��yO��2�>����>�F�=�m�<9&��4�x?�^?%��>3����B���^�I�X�I�վc�Žxî>A*�>�|=�c���eﾳAI�~�s���Z�Y^�����rh	�ć>_e�>��>�`��� �=di=0�=���<6I��L���w�>*��>U}?M?d>=J0>�c��ҾF�%?r�¾�-(���u�x3��3Z����>���<}�Ž��?BTH��'���5��9x�@?M��?�\�?텍?�?s�����ݏ�>̌>Ę+<���=��b���>"X����+��Q�q�X�l��A��e�/>>ؖ<P�B��k0��#%�9��'���a�c$ҽ���6"�oVl��\���C⽌=��f�:��\B�� _c�f�q����:���g�����@�Rz?���?L��<ֽD6�,���	���=)���~��5y��G��b���Zw��U�r�z�O�c�:�dJ	���>\�žq9�����������!>\��/!T?�x����|��:>�N�>:��=�*���+������{�d��tE?%�J?`뾓��[S9��|>u�<?7�>8>S��~���ٿ�>�?ò2?���j���\���?�%T�?K��?�Vp?���'C��~3�6����?��=�J@?PLR>���sd>��?��q?�"�����O���Q�g�!?UȆ?bP�G�> Nr>'Su>��;s��&�t�<C��~aU=�DF> c1�I�A�F���������=�>�>X�>�"軜N���>f���q��<c�WS�өE=�ws��?���g�9>�1>�Dz=EC^�m��wd�N�@?�Y�?B{?��??�����xľ��>d^���>��>�O绔�+�$`�>O?��$�x1-�+A'��� ?5��?�_�?[��?��g�b]ÿt���ž�"/�aG�<�">�J>�����=@��	��!=8Uc>[��>G�_>\�>?�>h>(@�=����<%�-G��������P���%���C�b� �⾴V0�,�ھijA��=���=I!�:f����?�Ϣ1�:������=_>}��>�]�>f?�<�>���>9q��	����Ki������򾓋��}.������̢<
��<YG�JF��6�=?�����A���?t(׼��=�^�>*��N >ߏd>_��>?;�>��>��=>n��=
9O>�G�=:ys>��=�����!���7�hU��ؐ9�C?�V�����G6���޾�^����>��?�;T>�?'�����Z�x���>�x1��Ec��:Խ��'�Њ>��>���=p���9�"���|�])����=/z�>�l>7����钾�6�^�=5��>�u¾��o>�ʏ=�R�>�ڀ?�H,?���= ��>!mc>�p>,���Ww>8�>?��<?r5@?��?��>@-(>u�?��zZ>�=���:��:2���Ld;��#>��e�;�_=p)�E�j>8!=�&�=�==�-�;��������>��??9o�>c��>h���\?���)�6��W>
'�$i�>E�>��?���>���>�"/>���� �߾���?�>��1>��K�qml�1���vQ�>�v>c\M?q�+?��H<�@^��:�<��=z��>�?��4?�^�>��>�ǌ�����Pοxg!�&0����F1*�p=p�K�W����>�B�>Zپ��<n:)>��>�.�>qˑ>��>�M�=/�G�4r�>]xX>�k�=���>,V<<_�bc=*�$>�c�<c��;���?���~GP��z.�:�𽀍��]˲�⿆���?�($?�1���7=/�f��������>�>gl�>��>��6=���t1M��I�2�D�I�?	�F?��>��Ͼ�T�<Ѕ�=��Y>�K?�M!>��>��ƾY���׾���<7ف>$6?pq4?0����k��A��V)����>:s�<Zk$=���?O�a?�<�qP���K�,�v�0�����=s@��B.����ZJ6� 澌���bپ��
����>Iߡ?��'�� >y%��������M�3��\�����>c�?�Ð>t������\���)�����ӷ��U�>���=%dY>��7?xm�>��6?�EY?@�,?mȽ!��>��>(��=�R>��?hrg?�/R?�b2?5��>&ݻж��B�ɼa^��+xX��� ��ꍽ(��=�	=���=�=>�(�=�;>��/=.ǽ��R����=�M�=�<�=`�;>�v>D(?jB/?Ќ����a=���CmV���<k>�Fg>��ν�����w�:9>�S�>�g9?D��>2������F� ����lg=b�?"9?�m[>qaԽ
��>�
�X�O����p�<>� �!T��/��e���� ���p>U�B>>rS>���?�`?��	?�W�;��4�vmо�Z��n͉���8��� ?.>��载x���J �O�h�rv����g��o��Ѝ#�)Z�<Is.=
�#>b�r>|�<�p>񤽏��=��j�ʜ��_����=>�2�>τ=?͇>;�d=q}��� �t�W?����S8^���<���7��đ�=���=��ת�>�̛����
7��������=�?��?Rל?ZW�9�{����>���>׼&=��D�|��m��>�I4�v��=�t�=���6N�O���S>z\�=�;o�l]��I��p:� �����T���I�N��y���w��%����	U=3:U�ͭ	�Sh;�jcs��=����
ٴ��/b��﷾�[ɾ^@�?,��?J��=�SD����[�U˾×�>ޅ�%����?	���~>���*����۾- 񾢡P���E��ٮ�|,�>�a����l��to��I,�|m|���<�gT?(+w�/(�&'��A�m>�>������գ��ܚ�|��9b?�z?��ԾHiS�T2̾c��>|�d?�a�=�?о��ǽ�'?q��?8,?`���ヿc��h<�^�?���?�2�?����.�{7�r����A!?g�->�a�?�����:澯j%>�0�?�҂?��#=�3���oj��
� ��>��?�:�U5�>&�>�֓>��==V˥�2�?�ꖾs�o�r3�>B�0��Р�$��Z�ƾ�tk>��*?k��>�����+��Y�?�*���}������<����=$��"D?�p��>�`�=���<,<��-��ʀX��ʛ�S�+?j��?��?`'?#ھ�ㄾ5Z�=Pݭ��9�>"y�>���Ɍ���\c>��>�T%�ps���:�nF�>���?��?��?����ʿ�웿  �������2�2��=��Y>�[�M�< �a>텤�.R�l#�<�C�>�~�>t��>�Wr>o��=�Z>��}�1�K̖�_���/qb�b��A��~H���P����O������&X�g�����=�92=��S�آͽz�<�?��P�<>f>�Z�>��-?�^�>��>ѹ��%���X4�u,�T�8��t��>����=�3'>�b�*Ӵ����7C#� �.?�b;��=|�?���=5>6=�o�>?�ƽ�v>л�>e��>f�>y,�>^�e>�p='QA>6q�=��+�w�C�y�p��⦿57������:��F�M?�Oe>7�A���c��������>�,?xh,>�M��x��"���`�>D�'�@�H�>�=��8���R>��>}ɻ�9���=ʁ/�Ѭ��ǋ�	�M>0w>9��ݶ;�4������>��¾�Y>�=>�v�>z:�?�?�q�=$��>��>s?6�6=���>s�<��h>�3?=�?�!A?��>o��=���)-�>Dmb>���Rr$�`����1B��r�=�w�<�t�=���Eo�=T�	q�<RB[>2���eݽj$=�!?��1?��><G	?�Sﾯ`��m)��ϵ=d��>�tn�<�?���>�?�>*-�>`�z9�������F��0�>^��=$}��}����ּ^��>�q�=�Wp?0�D?a
��>��nX>�J>�.R>���>��?V��>nhw>+>��"oԿo��Ad!�RuK�J��������"��9� �������׽����Ğ>;��>��>	�+>��=ga;>�>�t>Q�X����<D�=� �;��6�(u=@0�<$�̽���8ѳ=���=ǌ_�t�r������t������%?�u2?�7�����Cb�$s�ǫ^�2��>S��>�?˙?�9t>�T�6�_�}��\�)�>5�A?/?qѾ�M$>|佐�S=R�??
�7>���>��]��ͅ�9�k�� �2H�>��9>�n?�<ӾTXo��G�n�@��I{>�<��Ԛ?'�u?��龤�]��[��F~>�K�̾�����>�����Ty�8��
�;������ͨ�&C����>F�?����}@�<�>پ����IK����=�l<=5ɽ�y�>���>�%�	��2�q�R�{��@e5����>(�=�sJ>��-?D	N?�S>?�%	?׆~?d�����>m��>�>��>:?�^?UB?0+�>OY`>5�h�_;�A9
�J-���.����=J��=�-=MV>�3=����Y=�м2���A��<�e�=0�-��Q�=�TZ>�0V>��=m	?�_&?�X��u�W���S%����=��=N�\>��}��u�~*�<	:@>�&�>Ee*?���>�\
=)}ݾ��侐p��q�=��?�x1?��>���&�=Z�뾋�o�hjM=�4?>���P����eྴL���xӽ�Y�>Γ�>T��=��=6G�?��q?T�>��B�H�ӓ+�	OV�E���L3���H�=�G�>р�>�q�l+�i��"����OW��O�����T��?
>��$>�d3=x7
>�
x>m%��'��?Z�=s�R���l;�U�>G��>��0?�֞>N/�=�D�����LW?� ��;�v��'[��~0=|k>z`*>�־��r�Sƽ�ԗ�~����������>k��?��?᪛?�6޾����>���>�����վ� �<vU�xF�>��(>����F��>�<M{>3��=mT�|Q˾���+�������B�R`��ׂ�1�*���߾p;��x=�F��#bu������̼�>�r<w�W�z=�����'�6���g��[V�?ޑ?��۽�4¾�/�^m������>Z�:�����=��T8W��h� ������PF����d���	�O5�>���\����z���ܾ�8�=���H�Z?-Ҽ��� �)�G3\=G|f>@��=� ��E(�������-	���F?r?���w(8��u�=f�u>��6?��=�݇>,���<�a;e��>Q�L?eI?3z�� 掿F�q��;?��?��?�W?b ���<�gU������!�>;�>�O?]?�;t���ҝ=��1?��C?"�>x���Hp���C�>�Bz?���֬d>0�>���=v��:�hw�J\:�l񲾇V���>c��,I��Q{�������Q>l��>�>�+��ya��Ib�>��HO�w�H����.����<��?���((>��h>�,>�p)����������� �&�M?���?OzS?�`8?���������}�=���>���>寱=Gl�ܑ�>:��>�f�[�q�Ҿ�8�?q�?���?��X?/ym�[ҿV���0b׾9�����=XE6>��l>8+�<���>��к~�\��L���9>� >�=�>	�>�{�>h��>�#�>�0����$�/������h�>�j���
���4��o���d�r[��&ؾ�2����Z�qƴ���B�Ὑ�ͽ>U�\��>��=/�?}�?[��>�>�(> t���Ӿ� ��R�����6߾6�*��L�:g��X$l�Z�Ô^�1@��{�|�?
ڕ>�}�>['?��=C>��?K۽S �<s(>�"�PS�<;U�>��<�׿>L��>5C>�ͻ>M1u>�.i�{�{�ˢ�1�w �>d�+?)h�vF����P���*\���U&?!a
?:�e>Z�:� "����a��#�>t��K�վ~�4�u���c�&>���>��>�N�#�>	ޖ�2u�e0�>���>'�=����l��ʱ���*>pa�>z���!W>l��>��D?��t?mR?֛>��>��=h9�=�	=kGh>�>��>/��>i�N?6s?���>�>�?�zl��Ġ$�D.��)�����.�=�1>ti��g��=U�3>�X@>]�=c_<>�ƥ=g��D|���?B�U?���>ͯ�>j�w�K%��S��r�(�>b"�cZ4?Y�?R��>���>���>f�=ф=�n���f���]�>n�w>��t�c}��z�ڽ�l>�ɫ>{\O?0�?�s�ʅܽ�O]�!���g�>�?r�#?�|�<�XB���=bn�z���I�L$3��B�=G�(>̥�=�<�v�>A���?<�Iw�iҽ��h>�}�>���>���><��>�� ?���>��!>�i"==z<�"�<�)���1罘��<�[A=�|�=K �=�z�=�D9��ٻ�C�������-�ټ�Z�?��2<?�M?`׍�|^���i����~ں�I´>��>o��>1�>W�>�l��S�E�E��e�PM�>��i?��>��5��6�=W��=�;�@�>���>�{	>��I�"�	�x2���=��>`|??��>���jX��l�P!�Ø�>���=(b��j�?��K?Å ��b��:<I��j�R��>+K>1Qy�H.h>�;n����"���+���p��s��P��" �>4�?l��T˼Qھ���������޾�4ʽ�ȯ>��[?�?D�t�Mv�9V���"�8�＀^�>�3�>yqX=A�>��)?�L(?`0n?�"?{?}��w�
?tG���w�>�ٲ>z��>��>�y?�fE>�o>��)=�z�����ǐ�)��<\�3��=�a:>̠�=Ի�?K=�Ǡ=�����F�<d����=>�=�Ԩ=�w�=KL�=F�=��?��?НD��㼘p�������\>?RۺǨ�ԑV>@ר����_�>��>��?��?�b���O%����@'�������^?=�@?!�?�>Ypt��>�Z�4��zw���=�㷾b����4��J�78���>�>��k>�3E��҄>�Iq?�V?�s7?��u�
=5����p(��s��OrO=yC?��?*
>*� �8zg�Tჿ��%��{�D���S4��f=a�5��=�O`>0��=b
�>�?�>�V��0z��M�Q�2m��j��>&.>�c?)a�>`�<�G޾��辔G?����X�O���9ɾK�=��>��A>����ر?���|�)+���:��%�>@��?���?�7c?B�H������-Y>YyS>��>	��< �>�<q�.G��-:>E��=�z��	��.6A<�S>-�~>�����Ͼ�e�M�b��H��A[Z�=��
�NV!�	,��~�:�)��<�]��Gf�<�[]�Z�����־���F���A��T��<��<�#�����?D��?��8>��S\�ҩ@����-�=E\"�����5��v�m=�\ �ǀ��'Zr�t��� P�ŝA�OT$�Wß>��P�Wc����|��u,���:�S�P>43?�;Ⱦ�&����u�S=�@=>=M=��b]���
���;���S?�4?	pﾈ�����=�Q?�&�>4�>!	��]���>��4?��/?�x��`��Ʌ���3:�3P�?j��?�9? �#��hB�MY�D�ʾ�*_>)?W�>�ा핈�m���@
?��_?3��>��ƾ$�g�_eK�ڔ�>v�X?df���+>
\?*��>�A�&[x���T�վ�z;���>�g<o�3��H|��=����>@T�>��.>�_�F�a��c�>����<O�A�H������fi<]?���Q~>�c>n�>�A%��_���Љ�X�����J?C��?�R?Uz8?f��h~�ڱ��/C�=��>[��>0�=�
�o�>���>Sl�ͤr��q��%? ��?��?��W?�p�M������R�Až��l>�i[>)7>��J�DM�>��=�,>A�9��<�=���>�ϼ> ��>��>��>���>�����c&�3���au����7�1����ξOF��&��������;���cb߽�8=)�:!n�.�ʽ�d��� f�nѳ���0?���>�+�>$�+>�5�>z���`���Ј��gھ7���.�����dQ;�x`�yD��P�G���w��ݽ��,R?���=��>��>ܺĩn>�O�>h����i��%��=��n;�s8�'>Q�>#�<��>��=���>g�>F��Z���۶� ��R�=�B?K����������L�Ӿ�tξ7
?��>̤L>Q@����}چ�e��>>���G��q��o�1�Q(���>a>'8����9>a�<��r��>\ky>�*>�;=E��9����߽y²>�f���*)>X�D?>�p?��?�P?Ko>��>���7�E>Ys ��]�>�7������v ?��z?
>L?.J?-|	=�)��WqC��ф<��{����=zI�L_>�O=��<�)x��py0=���<�Yܻ��]<ԡ�=����L�.>%�g>��>�<?�6�>�)�>�N�G���>.����~�(����=T��>p��>��>���>⛒>4�씨=䩩���|�^4�>T>�
|��"K�nѸ=�>ć�> {J?+�8?��Ǿ���?@z��G'��@�>y� ?;G?�T�=F�c����c�)Bο68�_�(�GP=������^���b=X	�<-Cѽ{~���>�c�>֋R>Wx�>��>>���>=#�>ԣ�>C��>ah>W��=�	�=���<�۽���;��G�i@5�>/=o{�<�����d��q=S�x=�<����W�I��=?�?�̼[
}�/6o�5@������b��>[��>�|�>��>��=����S��FB��`S����>��h?P
�>;�7����=��=����;US�>�Ȣ>�>�i����������<(o�>��?}��>u�&lX���j����ń�>�"�=}C�~ݛ?=�.?#�����Y�*��=�������f>�ґ���<�l����%������x����i�����>ѯ�?訜�� a���9�G���	��0U澒b�K��>W�?L�?P%�=<��=�y6����a~>3s�=4��=���=��>j_?��%?�3h?Q�?�6?�U���?c��=���>3��>T?E��>�s�>���>p��>X}�=�w"<s�ny��;m��sr=��#�=>��>�<�?�<H�=�X=;8c��1<��<�tμ$1=ϲk= ��=�>�?>?ND���q��;����8k>�z�>��=[DD�����6̽�I$>vR�>�5?��>n���!��EL�'7�@<k�:�m?�=S?���>��>�%-=y�$��=���~=�:>�?k�{��N(�T�N��{�Hr�>���>�R�>��>�Sl?�^o?�B?��?�c����R��܅��=�>�4O?F�@?�C�>���ݡN��o��U9+�jh
�K�/���!��=�s���*U>62�>�5�=f�\>dqb=D(Z��N���I>j����؎>V�>��>1IV>���=���^h`���I?Q���{\�����[о�R�g�>+�<>Y����?�s�}�/���L=�Z��>�}�?`��?�/d?ɤC�,���\>&@V>�>��/<%w>��Z�`]����3>���=�~y�6����;�]>�:y>_ɽ��ʾ����G�Oʺ�f,h��+þ�9#�_"�SR���]��3����&>�{���ܾk��X�[��^��_=y��"x���7�����%��?l�?:h>^�@����ڤ>������/>�ý����
�ƕ޽O�'�pX�����w��GU0�uG��5�IN�>��[�%E��G}�P
(�x4��oh=>��.?��þ�0���e�8�u=^�+>Q�<���-��G���*��5�W?sm:?�+�i&��xؽ�>�4?�J�>P� >����rm��b�>�4?�E-?��м�ڎ�!����i�냻?�e�?V??��L��A������i� ?oy?]��>ɳ���ƾZ���	?�X:?&�>�F�}<��{�����>"EX?�lN�C�^>oz�>�ٙ>�	������A1������L;��<>[V��I���h�OZ:��E�=�1�>��u>:�Z���Ib�>��HO�w�H����.����<��?���((>��h>�,>�p)����������� �&�M?���?OzS?�`8?���������}�=���>���>寱=Gl�ܑ�>:��>�f�[�q�Ҿ�8�?q�?���?��X?/ym�[ҿV���0b׾9�����=XE6>��l>8+�<���>��к~�\��L���9>� >�=�>	�>�{�>h��>�#�>�0����$�/������h�>�j���
���4��o���d�r[��&ؾ�2����Z�qƴ���B�Ὑ�ͽ>U�\��>��=/�?}�?[��>�>�(> t���Ӿ� ��R�����6߾6�*��L�:g��X$l�Z�Ô^�1@��{�|�?
ڕ>�}�>['?��=C>��?K۽S �<s(>�"�PS�<;U�>��<�׿>L��>5C>�ͻ>M1u>�.i�{�{�ˢ�1�w �>d�+?)h�vF����P���*\���U&?!a
?:�e>Z�:� "����a��#�>t��K�վ~�4�u���c�&>���>��>�N�#�>	ޖ�2u�e0�>���>'�=����l��ʱ���*>pa�>z���!W>l��>��D?��t?mR?֛>��>��=h9�=�	=kGh>�>��>/��>i�N?6s?���>�>�?�zl��Ġ$�D.��)�����.�=�1>ti��g��=U�3>�X@>]�=c_<>�ƥ=g��D|���?B�U?���>ͯ�>j�w�K%��S��r�(�>b"�cZ4?Y�?R��>���>���>f�=ф=�n���f���]�>n�w>��t�c}��z�ڽ�l>�ɫ>{\O?0�?�s�ʅܽ�O]�!���g�>�?r�#?�|�<�XB���=bn�z���I�L$3��B�=G�(>̥�=�<�v�>A���?<�Iw�iҽ��h>�}�>���>���><��>�� ?���>��!>�i"==z<�"�<�)���1罘��<�[A=�|�=K �=�z�=�D9��ٻ�C�������-�ټ�Z�?��2<?�M?`׍�|^���i����~ں�I´>��>o��>1�>W�>�l��S�E�E��e�PM�>��i?��>��5��6�=W��=�;�@�>���>�{	>��I�"�	�x2���=��>`|??��>���jX��l�P!�Ø�>���=(b��j�?��K?Å ��b��:<I��j�R��>+K>1Qy�H.h>�;n����"���+���p��s��P��" �>4�?l��T˼Qھ���������޾�4ʽ�ȯ>��[?�?D�t�Mv�9V���"�8�＀^�>�3�>yqX=A�>��)?�L(?`0n?�"?{?}��w�
?tG���w�>�ٲ>z��>��>�y?�fE>�o>��)=�z�����ǐ�)��<\�3��=�a:>̠�=Ի�?K=�Ǡ=�����F�<d����=>�=�Ԩ=�w�=KL�=F�=��?��?НD��㼘p�������\>?RۺǨ�ԑV>@ר����_�>��>��?��?�b���O%����@'�������^?=�@?!�?�>Ypt��>�Z�4��zw���=�㷾b����4��J�78���>�>��k>�3E��҄>�Iq?�V?�s7?��u�
=5����p(��s��OrO=yC?��?*
>*� �8zg�Tჿ��%��{�D���S4��f=a�5��=�O`>0��=b
�>�?�>�V��0z��M�Q�2m��j��>&.>�c?)a�>`�<�G޾��辔G?����X�O���9ɾK�=��>��A>����ر?���|�)+���:��%�>@��?���?�7c?B�H������-Y>YyS>��>	��< �>�<q�.G��-:>E��=�z��	��.6A<�S>-�~>�����Ͼ�e�M�b��H��A[Z�=��
�NV!�	,��~�:�)��<�]��Gf�<�[]�Z�����־���F���A��T��<��<�#�����?D��?��8>��S\�ҩ@����-�=E\"�����5��v�m=�\ �ǀ��'Zr�t��� P�ŝA�OT$�Wß>��P�Wc����|��u,���:�S�P>43?�;Ⱦ�&����u�S=�@=>=M=��b]���
���;���S?�4?	pﾈ�����=�Q?�&�>4�>!	��]���>��4?��/?�x��`��Ʌ���3:�3P�?j��?�9? �#��hB�MY�D�ʾ�*_>)?W�>�ा핈�m���@
?��_?3��>��ƾ$�g�_eK�ڔ�>v�X?df���+>
\?*��>�A�&[x���T�վ�z;���>�g<o�3��H|��=����>@T�>��.>�_�F�a�Ib�>��HO�w�H����.����<��?���((>��h>�,>�p)����������� �&�M?���?OzS?�`8?���������}�=���>���>寱=Gl�ܑ�>:��>�f�[�q�Ҿ�8�?q�?���?��X?/ym�[ҿV���0b׾9�����=XE6>��l>8+�<���>��к~�\��L���9>� >�=�>	�>�{�>h��>�#�>�0����$�/������h�>�j���
���4��o���d�r[��&ؾ�2����Z�qƴ���B�Ὑ�ͽ>U�\��>��=/�?}�?[��>�>�(> t���Ӿ� ��R�����6߾6�*��L�:g��X$l�Z�Ô^�1@��{�|�?
ڕ>�}�>['?��=C>��?K۽S �<s(>�"�PS�<;U�>��<�׿>L��>5C>�ͻ>M1u>�.i�{�{�ˢ�1�w �>d�+?)h�vF����P���*\���U&?!a
?:�e>Z�:� "����a��#�>t��K�վ~�4�u���c�&>���>��>�N�#�>	ޖ�2u�e0�>���>'�=����l��ʱ���*>pa�>z���!W>l��>��D?��t?mR?֛>��>��=h9�=�	=kGh>�>��>/��>i�N?6s?���>�>�?�zl��Ġ$�D.��)�����.�=�1>ti��g��=U�3>�X@>]�=c_<>�ƥ=g��D|���?B�U?���>ͯ�>j�w�K%��S��r�(�>b"�cZ4?Y�?R��>���>���>f�=ф=�n���f���]�>n�w>��t�c}��z�ڽ�l>�ɫ>{\O?0�?�s�ʅܽ�O]�!���g�>�?r�#?�|�<�XB���=bn�z���I�L$3��B�=G�(>̥�=�<�v�>A���?<�Iw�iҽ��h>�}�>���>���><��>�� ?���>��!>�i"==z<�"�<�)���1罘��<�[A=�|�=K �=�z�=�D9��ٻ�C�������-�ټ�Z�?��2<?�M?`׍�|^���i����~ں�I´>��>o��>1�>W�>�l��S�E�E��e�PM�>��i?��>��5��6�=W��=�;�@�>���>�{	>��I�"�	�x2���=��>`|??��>���jX��l�P!�Ø�>���=(b��j�?��K?Å ��b��:<I��j�R��>+K>1Qy�H.h>�;n����"���+���p��s��P��" �>4�?l��T˼Qھ���������޾�4ʽ�ȯ>��[?�?D�t�Mv�9V���"�8�＀^�>�3�>yqX=A�>��)?�L(?`0n?�"?{?}��w�
?tG���w�>�ٲ>z��>��>�y?�fE>�o>��)=�z�����ǐ�)��<\�3��=�a:>̠�=Ի�?K=�Ǡ=�����F�<d����=>�=�Ԩ=�w�=KL�=F�=��?��?НD��㼘p�������\>?RۺǨ�ԑV>@ר����_�>��>��?��?�b���O%����@'�������^?=�@?!�?�>Ypt��>�Z�4��zw���=�㷾b����4��J�78���>�>��k>�3E��҄>�Iq?�V?�s7?��u�
=5����p(��s��OrO=yC?��?*
>*� �8zg�Tჿ��%��{�D���S4��f=a�5��=�O`>0��=b
�>�?�>�V��0z��M�Q�2m��j��>&.>�c?)a�>`�<�G޾��辔G?����X�O���9ɾK�=��>��A>����ر?���|�)+���:��%�>@��?���?�7c?B�H������-Y>YyS>��>	��< �>�<q�.G��-:>E��=�z��	��.6A<�S>-�~>�����Ͼ�e�M�b��H��A[Z�=��
�NV!�	,��~�:�)��<�]��Gf�<�[]�Z�����־���F���A��T��<��<�#�����?D��?��8>��S\�ҩ@����-�=E\"�����5��v�m=�\ �ǀ��'Zr�t��� P�ŝA�OT$�Wß>��P�Wc����|��u,���:�S�P>43?�;Ⱦ�&����u�S=�@=>=M=��b]���
���;���S?�4?	pﾈ�����=�Q?�&�>4�>!	��]���>��4?��/?�x��`��Ʌ���3:�3P�?j��?�9? �#��hB�MY�D�ʾ�*_>)?W�>�ा핈�m���@
?��_?3��>��ƾ$�g�_eK�ڔ�>v�X?df���+>
\?*��>�A�&[x���T�վ�z;���>�g<o�3��H|��=����>@T�>��.>�_�F�a��c�>����<O�A�H������fi<]?���Q~>�c>n�>�A%��_���Љ�X�����J?C��?�R?Uz8?f��h~�ڱ��/C�=��>[��>0�=�
�o�>���>Sl�ͤr��q��%? ��?��?��W?�p�M������R�Až��l>�i[>)7>��J�DM�>��=�,>A�9��<�=���>�ϼ> ��>��>��>���>�����c&�3���au����7�1����ξOF��&��������;���cb߽�8=)�:!n�.�ʽ�d��� f�nѳ���0?���>�+�>$�+>�5�>z���`���Ј��gھ7���.�����dQ;�x`�yD��P�G���w��ݽ��,R?���=��>��>ܺĩn>�O�>h����i��%��=��n;�s8�'>Q�>#�<��>��=���>g�>F��Z���۶� ��R�=�B?K����������L�Ӿ�tξ7
?��>̤L>Q@����}چ�e��>>���G��q��o�1�Q(���>a>'8����9>a�<��r��>\ky>�*>�;=E��9����߽y²>�f���*)>X�D?>�p?��?�P?Ko>��>���7�E>Ys ��]�>�7������v ?��z?
>L?.J?-|	=�)��WqC��ф<��{����=zI�L_>�O=��<�)x��py0=���<�Yܻ��]<ԡ�=����L�.>%�g>��>�<?�6�>�)�>�N�G���>.����~�(����=T��>p��>��>���>⛒>4�씨=䩩���|�^4�>T>�
|��"K�nѸ=�>ć�> {J?+�8?��Ǿ���?@z��G'��@�>y� ?;G?�T�=F�c����c�)Bο68�_�(�GP=������^���b=X	�<-Cѽ{~���>�c�>֋R>Wx�>��>>���>=#�>ԣ�>C��>ah>W��=�	�=���<�۽���;��G�i@5�>/=o{�<�����d��q=S�x=�<����W�I��=?�?�̼[
}�/6o�5@������b��>[��>�|�>��>��=����S��FB��`S����>��h?P
�>;�7����=��=����;US�>�Ȣ>�>�i����������<(o�>��?}��>u�&lX���j����ń�>�"�=}C�~ݛ?=�.?#�����Y�*��=�������f>�ґ���<�l����%������x����i�����>ѯ�?訜�� a���9�G���	��0U澒b�K��>W�?L�?P%�=<��=�y6����a~>3s�=4��=���=��>j_?��%?�3h?Q�?�6?�U���?c��=���>3��>T?E��>�s�>���>p��>X}�=�w"<s�ny��;m��sr=��#�=>��>�<�?�<H�=�X=;8c��1<��<�tμ$1=ϲk= ��=�>�?>?ND���q��;����8k>�z�>��=[DD�����6̽�I$>vR�>�5?��>n���!��EL�'7�@<k�:�m?�=S?���>��>�%-=y�$��=���~=�:>�?k�{��N(�T�N��{�Hr�>���>�R�>��>�Sl?�^o?�B?��?�c����R��܅��=�>�4O?F�@?�C�>���ݡN��o��U9+�jh
�K�/���!��=�s���*U>62�>�5�=f�\>dqb=D(Z��N���I>j����؎>V�>��>1IV>���=���^h`���I?Q���{\�����[о�R�g�>+�<>Y����?�s�}�/���L=�Z��>�}�?`��?�/d?ɤC�,���\>&@V>�>��/<%w>��Z�`]����3>���=�~y�6����;�]>�:y>_ɽ��ʾ����G�Oʺ�f,h��+þ�9#�_"�SR���]��3����&>�{���ܾk��X�[��^��_=y��"x���7�����%��?l�?:h>^�@����ڤ>������/>�ý����
�ƕ޽O�'�pX�����w��GU0�uG��5�IN�>��[�%E��G}�P
(�x4��oh=>��.?��þ�0���e�8�u=^�+>Q�<���-��G���*��5�W?sm:?�+�i&��xؽ�>�4?�J�>P� >����rm��b�>�4?�E-?��м�ڎ�!����i�냻?�e�?V??��L��A������i� ?oy?]��>ɳ���ƾZ���	?�X:?&�>�F�}<��{�����>"EX?�lN�C�^>oz�>�ٙ>�	������A1������L;��<>[V��I���h�OZ:��E�=�1�>��u>:�Z����?Y谾T����ۅ�#�'��$��>'.>�id?��Z��&���l>��?N���Ӭ��+��#`�ހX?ɵ�?yn?��?޸˾լ��%>��z�6Ԁ=T� ?����䢾�K?Z
?<`۾�0��$�%��?�o�?ۇ@�:?CTU�O^Կt�B/��ǅվ��g�̂�=/�#>����Rv=~(ʽ	�4<�\���i=\��>���>��>j�.>��x>�n1>2����`%��2��r��W�0����-�͘��% ���T���P׾�ٵ����9Ľ��2=�i����"�Y=ޚ���&>�N�>���>�Ĝ>d�E>�9>��e���Ծ-{|�����:�%���L� �`�ھxꐾm�/���m�c�G��M��QY�Υ?�+M=5S�;BE ?"R�N%�=�ǎ>}g�;p$�=oa�>��=6[+>�H>Q�>>��>O��=1��=-8�=Ci���e� c���Q
�군������HV?�i�k|��j��3/���Ͼ��>���>I�5>˺,�@3���9�����>�=���ʼ���[;�K�/>7T�>:�M>�,%��� �N�F�=�V�k<�}�>度=%�?���
���3�K$�<��>�2��ũ<���>��D?�T|?M�9?xȼ� �>�Ț>ю�>��ڽ�P�>���>�L�>i� ?�q5?$w9?;�>�}>�2���B��A�=�n8���{�m#�!��S� 1׼��Z�.\�=��7>���=M��2Ӧ<�B=q���ea�<�;?(y3?� ?	�? 1��.�]�G��W�.Xt>�켾o�>I�>��-?4�?�� ?РT>��=Ag����>��׾>�(c>�D���o�$��;��[>i�=0�?IH?�&��Aﾛ�Y=7�w=���>�W?��>?f��>&>C���,���ʿ.f۾���(��<�-T�%^�2_������1�_�UyQ�Vr��3�,��K�>z��>���>F>�=���L��>���>��:>:t=�-�>��@>�u��* ����=^=�{P=�w_�Tď=:=��"*��6��	�}��}�d���0c�<��?��E?6���n��T���q��\=���>U\Ž�K?%~	?ea�=�$7�₿���������['?���?o��>sõ�:��=a/�=�>"	?'�?Tc;�M_�&��>E�ɾ$:?>B��=�?0.�>;a�=zv&�u�j��(� ��>��>2�=�-�?�>\?�yF��A������+j��R�DN��|9�;��=K@վ��;��pV��@A�3�3����i��>��>s��?�4S>��>{�ƾy+������������:>t?�@b�[=d��#ͽI?'�8��U2ʾ�yP=ǉ>げ>��=<K?�"?Ynv?�Kt?W�+?�J����9?V/��)�>�p�8�*?�8?M}A?�t?�ng>�jn�+�ʾUֽ������m�<�R$�=�%>�K>[)��ٰ�:��="��=N����( �'xa=-�/�;��4>��>��?<�#?TW�������4(��ϽP!�<�
>�e>q�����f��ɹ1ރ>�?�"2?#+�>]��=�侦_��Q��ZI�=�X?�/?�^�>f�X=�}�=&d��2�z�o�=%^>:L��I��)����������j>8�>� >��>ww�?�=�?5X?�����@������T�NTN��B�>��I?(�x=�d��*��u�2����c m�����;>n4�y�/�ȵ>��8=Z�>��>�P>��=(%=ɏ==�����t|�>�	�>�rF?n��>��>��h��(���T?���)0�T�龯����W���t>�l�>��:�?�ཹA�7а���c�1Q>�ΰ?�>�?_H{?��9���(����>H�>�>S�ؽ���|��)=^�Vʁ>�m>�J��AU�����9�g>)��=z��ѹǾ@�վ� 2��ܯ�͑a�tb4����[����l�r�2�4pD>�y<������VW�m�B��y�������I�@��������K���ap�?�h?Vz�=���B�8����`��>�S���R<�<پ��=�M�����g�R��X' �����^6�{o�>H6�N���'��]J�I�E�F��M�u?:x��Ճ�=R��[~>쬅>���F�������G�������?Go?K�n�5T�~Q���h�\?�?ok�>Z�՗��� �>L?�f_?rP��S��������>���?��?7?�N�k(>��P����P��:	?	�
?.*�>rXM����mk��ĥ?��!?g�>��	�e���f��kk�>-_?��,��->ʮ?��>>Pk�/!z�˴2��iξ�Aн D>�}ӽ��%��t��Vd��h=�x�>��F>ɔk�����x�>�꾆�S��/K���
�~|5����=��?�]��><�a>�n7>t�'�s��k|��`D2�� E?޼�?* V?�q2?�i��־�r��D�<��>|��>�=�U����><�>2X��>y���oW?2v�?|�?�W?F�i��uԿ~����ľ��ƾ@Α=c�>��|=3��	#>�M>���<���*J>��>��v>���>�>�u>��i>�����'��b������Sq�1B!�O�$���p�/O⾼�Y�S�$�NK��˾�QB=����������4����c=�|��Uw>�1�>��>��>�>�N>X���{�����I���-���%�e���㲾�����nG�)�7�Z̰�:��׸?���=O�8=0S�>�����ե=�!q>�[P=:Q>��)>uQ��G�>��>#�@>y�>�37>b�=��=O�$�Y-��qԊ�W!�L�x�۾��?�ȁ��	��$lw�Y޼��EI�" ��$?��>����S竿�夿ҹ??l2=�~��N��p3���>�E�>��>'���B�����L�'�'����>��>6�ʽg4�}�Z��H�=Z&?.�¾y>Gh�>��F?-^�?��)?��>�J�>�X>k��>*>�����>�>���>�a3?#">?��8?oW�>g?1>sXl�;�D��ab>�̼�I,=O���[�6=A�+�"�?<��[�2�/=h��>wX��cT���ه=zo�9Qѻ��9=J?�
8?1�>���>PfŽ�t9��{&�J���@>�ν���>�$�>�?"?]?�Ǎ>���=m����ž���>]e>�v��67p�X�Y�T�=���>�j_?CM�>�ꬾڈw���_>��=��?i��>��?&�>�ȸ>�+�����J俪y��|)�{N���.�<%��!X�P�=\񽽔Q��S����2j��r�>躲>�f�>Pĭ>7�>��d>K��>`6�>ݹ�=����s�&>�u�<1ʶ;7�=���W3 �-?ս�SQ>`���6��׼WdJ=K<ڽ`��=l�?�r?rH�Yν*�Ծ�^�����W��>�p�>f�?_��>�>����d��5_��"���d> b?F�?y����=2�=���=Ο�>��>��h�"vؽ��5=YJ��(T,�wy>1?T��>�iǼl� ��Pd���]p>mn�=GW����?g�U?�[�l������Z����i7=�����*a�:;�_��\9J��W�
�'��A��fJA>.��>� �?��;٠b>�ゾ1ܛ�>�v��@����Ľ�V<���>��\>jXU��(���b	�Ӕ��U>��F;ܱ�>"wq>H�>�A1?�:A?b*�?�ob?S# ?�I��sm??�S='�>���3H?��?� &?�h ?���>�c޽Q`^�K����䕾ה�=�Bu�Y�=�6T>�x=>i��N�R>�	{>4E^��������=�T����<�2>b�>�S�g�=Q?X?6B�Ӓ+=�J�=��_�B=���=���>�>U�e�������̭>��?Y<?�>�f>V�ƾ�߾&��}����b?��??���>���=I�=e1�֦�3P>	l>�\�l�\�G�Ӿ����of���)�>�"h>ŉ=�9k>��?��_?��5?# ���M���[�T.��yW���*>��?��G>Uኾ ���6�<�޽X���k�:Z�&q>T#p�#�<h�=qPP=���>���>T�V=��=�jT>�p�̞>+X�pJ�>;�w>�@&?���>Jvi>:ė���_�I?�����j�6 sо�S���>E�<>��8�?�����}���H=�d��>*��?7��?9?d?I�C��)�1�\>)LV>��>�(/<w�>���؂����3>[�=�|y����vf�;m]>�Gy>�ɽ8�ʾZ3�=�H�U���>BR�N�N��
�U���茶Xm
����WF7��]�{��)5�S�X�/ ����½��R�z/(�^Xƾ����֎?,�?/���ͽ*���)���w~�>����'�"<�ѾC��=򑖽)MӾE�Ҿn��Ֆ��5��i8��k�>Q��M����K����+��&� �~>�%�?�J%�����J��b�>�@�=P-�;��þ"'���C�����;�&?4?�';����PA�Z�ݼ�b�>T6P?����y��w�?�4?��>��\<������g�P[�?���?wF?:a�mN�m���[�4:P>ƜV?k��>ß�7ɵ�%o����B?��>�r>�HI�>p��<����B?�d?�Ⴞ��>8�#?	-?DM��:�z��
�����L�=bJ�>���O��F|۾�s� *�=�h�>mF->���پ��x��>�B��N���H�'�����7C�<�z?Z��a>�-i>B>�(���Q̉�����L?���?r�S?#b8?dN�����\h��]��=w�>AЬ>�w�=���p�>���>��fwr���,�?�I�?U��?UZ?|�m��Կ8����㨾���H	2>s��=p�=V�ؽT2�=��<Xͅ������>
�>B�P>�n>�a>)nx>��
>�̈���/�����!.���T<�������W����	 ��T�.��ܾ��1�ĽR��jя�Y�˽���N��@��K��>�װ>�$�>Ei>\�>{�>��Z�ʎ���ռ�y�Ҿ'lT��:��ʫ����	�����@l��bN	�iyt��~ �?��>GT�=�r�<q?�`�7l�=�ʜ>H�=s�>1#>�뽑�>*џ> Ou>H�9>w!>�|��tb=B �=�d��sT���S�'�Ⱦ�瓾2\�?��Y�l�X�s�������E�E��=�H*?��%>� ?�����	��Os$?�>�@�ղ6�;�F����>2g?���>�Y��'��@Ǿ�=���E�=]��>q�>JN��;��Z��=ua�<Sc#?��%�c��{�>�'?<�q?�[?A.�ɊO>Á�>���>�$�~�d>i�켌5_>�Q?s�e?�M?76)?_�=J���[1�9��������r�����l��8�� ��$������=K z�H�׼E��=%�;=�v<?)�=�` <��>�=H?���>F��>_�˽Sr=���C�i�d��;>U���a�>��>^�#?��?|��>���=�Z����������>� )>�h��y���=���>���> *M?�g8?�	>
O��+��ѫ�>g�>_�?�7[?�,�>�H�=���<D>	�koѿ@p#�:�'�7�ZU8�7P��3��q�d�I<Z;A������n<k�<>�S�>	Rm>��H>�>��
>̲�>��G>�l=�>�=�N<��;����툃=�����<�F��'�<���j�ý蕋��9��L
�
�A�T���?�?�8�v���mn�� ���O�����>���>�1�>�X�>4��=���W���B��L����>�mh?.�>�<�&!�=Iy��I�;b�>�>sL>�v��R���w��N�<r�>�?`N�>����qZ��n�������>^d=�yJ<(�w?�;?�.O�F��8Q���4��r#���s=��V�s�n�l-�$����sq�U5��L2������,>K�>ײ�?�,�<��>���m=���'���-��f����=2?�,�=qЦ�/�*H����%���4�~<�n�=�z>R&�>R1g?C�?ok?&>0?��>�p���X0?�\�>��?P��>��!?�|?��?Z��>�X�>�ϫ=i�=����(Î���<�H�GC�<]��>DqO>s��=�=�9�`�7���۽�w�݃��Qy彄�=0�^>�y*=hj>?�b$?;��A7�k���H^� �<��=eON>i�F��z_��R8<�=g>hj?�<0?���>�y=�w۾2ﾀ������=D�?�$/?0�>�d�;}�=ٔ뾱�~��=�U>g�n����������:R���>��>��=7&�=��?��?|�8?��^�FEu�۞}��-G�ԁ��1}�I�>yF>![�����r�;����,V�����~`�bs��w��=x�=}v�=f� ?̟�>q��>g�=8K�>Ogc�Z��=]�N�T��>[ ?��6? 7�>�1>LPѾ���%�I?�:��#� ���Ͼ�c��F>��:>�W�=?b.
��}�"���̊=�?�>��?F��?�Fd?$6B������\>�U>M�>�<�=�h��,탽�X5>�8�=]{�������;4\>��x>��ƽx�ʾ ���K���ٿ��k�����Ò3�b�ݾ��о������<���c��G���Tɾ���Ԇ�Y���)q��W9�.u�\m��ǆ?��n?1�=e��R�?�(�nV���>$�n��;���ՠ����=gs2<v��Vj~�G���K&��P�4�%����>�6'>���������O��9��a�>U�?��Ͼm�6��L���>�ޠ=��z>�g���!���'���1��>�n?���
(=^�>�3}�?�l>�>��]��q��=k�=6<�>vB?���>�mܽ�˟�����-�/��?���?�8??��C�^�?�/��X�*�� ?z	?j��>�=��[�Ǿk
�	?6�7?�
�> ���ֽ�y'�>ִ\?� U�W\^>��>�h�>��������_��A���Mμ$�N>�����!�Ԉa���U�Hl=+��>��q>^Cc��Ū���>�꾆�N���H�����:�̉�<�o?���1\>��h>�>ζ(��!��Oԉ�\v�v�L?8{�?juS?�68?�J�����#����=FC�>��>5~�=�M�@t�>���>��辤Br�+ ���?->�?��?�MZ?�m���̿Z���M驾�������=k{>VQS>���1=
��=���<%!����_>c��>��i>���>f�v>�Y>ŐC>������%��K���Ԑ�7�D�������ϧl�<��A�P���	�q���>�ľ%.������27�����r��xμ�\����=X�W>�>^Z�>��=��S>��b����Vu��)G��U���o>���_�X�\���X:��eV#����Rv ����>��=����?���<nV�=�?�J�<�>�Z>e_�=���>[��>�1>acD>)P>$�>4�F>�)=�-��)����Z������(d<ᆊ?��9�v�2���T��#V�P����h�=��7?Y;�>��-������1�?�;Y�Ѿv�d=s{�ޖ1=��?F	p>����8 '=���}�ý�=�k��>�҉>�CڽŮ��Ƭ��Ӣ>�m�>lȾ�f�>��>��Z?��?�O?������>2؈>;u�>�u���ٔ>YU�>)��>�4?�:[?]�Q?lk�>]h=������:D�=f�����='b+��8��S��xZ<��q�Υ�a�;5ot�M��6>h�<>��=4d�=5P�>a�8?���>��>+�1�^x?���L� t�if>\|��T�>Ѡ�>�o?, ?q	�>*>D�>�����q���>׈6>��\��w���8��΅>��>�J?[�+?��Q���`���:=��=R�>Bi?��'?t�>��!>�	��HM�Q�ۿ�R��t(���뼈C7=��=H�m�������}= �C�)s����ļ��i>���>���>�qm>	=y>��>4��>C�p>���=�}�<��&���<wf���:>��>aL��bs���c�<J��=����V���P�ݽ]�8�A�R�z_,��?�?� /���hh�����s��Y��>4*�><�>�t�>'��=ĉ��U�d�A���I����>.g?��>��:��=��<"'�>r�>?>y�m�m�3����V�<���>��?9P�>����Z��8n�?Z	��Ҥ>��=0 ����?�ce?v&�iX���!%���_��߾�^>6н���������C?��H,����4���D�g>9��>ݸ�?�z�=�=�ֹ�3���Ë�/(Ӿ�=ct`>�I?�\->"׾F���.�"�dD辒���N�a<]�>�/>i%�>�{.?��?uLg?5,?��$?M�����>��=B��>��>A`?�M.?�R?���>nV�>=4�>D�=l꽫<����p���2���T> Q�>sc>`Ѽ����S��G(z�wSҷ�B=(�2=�� =�m8=r"���D>�Cf>O?}�?������D����A�f��v8>
��=윺7�j��B=�x1>_��>CT?6�>�{ļ�}�N�ݾT����=�?�RD?���>�wt<^�=��>r��m�=�|>͚x����Ts�s�ɾyl���>q+�>�>7o�>�w�?��>?HH;?�����_�-��=0#��k�<��G>�a3?�?�ꔾ�þ��\�����K�����U>������n[�<���=f�>��=ݱs>ݢ>D%�������>���< ?/�>�z?u��>���>�������I?ᘡ��h��젾/qо�I���>��<>�
���?�����}��
��2F=�,��>Έ�?h��?�?d?l�C�(��\>uJV>;�>/<*�>����|����3>}�=�y�^��G:�;X]>�Fy>��ɽ��ʾN/�ށH��J˿M�`��O@�s���G���с��ʣ�bCM���j�>����f��ڭ��(����S���#7ս��潏z����2[�?�N�?�As��д�L�7�:P)�>�.v�>[���{�������J�b=�I��1��������\��9�|Gb���[�3m�>��.��+��X���D�F����]P>�??�Q��
����*�3��=%��=:n`=cw۾�g��49��P����0?e�?��þ'8b��;��U>���>�>�h �IB��V<C>�u�>}0?d�?�C���`��2�ͽ�W�?\��?&A??�YB�;�A���Q<1�9��>�� ?���>�����^��t^��?A�,?���>٫�ǽ��ae&���>(X?�[g�S�Z>/b�>��>�;n�������R�Z���k���	C>��<��$�G�c�Ӂ���uQ=�Ŝ>�J>�`-�f����>�߾��L�yE�_	�$�"�]6�<:� ?�B�E&�=,R>�c>:�"�\Ќ��.���4��FG? ��?�S?T3?�o����쁽cO�=~8�>��>&��=Jiܽ!ϒ>i$�>�����x����?1T�?�>�?"+S?_�m� ��������X����u�/>�B	>��>js�v>q��14�ʔ@���D���-��>��>-�Q>�Hi>�8�>Ǎ>���z9)�������J"2�/�-�Qb �~h����E�-ա���"��Z��Ⱦ-���p��cα�zk���ٟ�'xz��M>c��>6R�>�l}>�>oO>ֵx��E��e��㻾�G�l�c��������@P��^��+z*�eFs�!L�rV?���<��'=��>@�ս>
�=c�> �6>h!}>��3>{���#�>x �>ݘ3>f�>��Z>�=��<c�>�Ot�r�� �"�x��%;[$X?B�_>J�ߤ:�53�"�'�A� �~w
?]�>贾������i�?��>2ᘾ�,H�n�\>T3�>Ȫ�>{��R����}��6�nu>��U>F\�>~������Qߤ�\|�=<?w����>��>R�X?�?}�C?�wt���?�r�>h��=� �M�>�� ?�>-Z?�^?��3?�y�>[�>R�_��!�	�ֻ<R��m?����T���0��BɽHf�=��J�Ľ��+>9>�`�=wִ=���=��=�9f=c*�>ye6?8��>X��>��c6�pP���8�gr�=b%���a�>���>[?{Y?O�>:�>�>r���վD1۾�K�>�>�<H��v������>�>��G?F�0?�9<�!���:�F���=��>u�?��0?F~�>��%>�]�b8��H߿h5�o���=T����=߭u�L�Ͼmy���)[��Ҫ���ǽ�ă>�C�>ԕ�>��>��>?��=&��>��>�=>����C�ƽ�Y<ő����=m��=�x�{~�:?�f>rk�;�,ؽ��o������,4�_�I���a?��?����p����k�����n1����>���>��>f�>C�=�����U���A��J���>��f?���>W�6��r�=�
�mQ�:Z�>��>��>e�m�X#�@��e��<L��>-<?�U�>��?n[�"o���	�v�>� �=<�ż�x�?U7d?M�*�ݟ���O�Z�0H��vG>��[���ջ�B3�f�9�����!� $|���O>��>�O�?h 1�up�>&�r�Q���������/_��N>+-?���>���H�ƾ�gԾ.0˾U����Ϛ=�C�>�Uh>���>�ie?��+?9�a?�m5?.ׄ>.�g���?b��>��&?]��=���>�&?h�?��>pW�>"t��酾�]��L��g==���Q�>��>�2>+��<쎲=��>%��+ސ<��4�
�:=u��=��=��>@�9>��
>x�?U#?����s����ļ����<��=�U>_��
V��X�{Y>��?�0?$��>�Q�=�۾���������k�='�?E�.?�e�>y\��n=|��_�g�ڛ�=�?K>�-p�AU���Z徎��}�ཹo�>���>9��=��>�V�?(�A?r]6?�N���r�������F���z���=L	(?�?d��=������G���o���W������n>]fD�]ʓ�������<r�?QQk>��%=.{>��K>�MҾ�ݣ=�8x�"?�>�G�>:��>��>2M�>V�%Y�3�I?����pd��㠾�Wо�����>��<>����?�����}�0���?=���>@��?���?�>d?2�C�j�;�\>�*V>��>*�.<��>���5�����3>��=�y�J+��K�;�J]>�]y>�kɽ\�ʾL1�k�H�A_��	�D��:k���'۩��'�����u��xA�@(�G��������ؾࢴ�B�j�9R���6��Ӿ����?⮑?�d�=���� +����Ѱ�_��=�ϵ�Yl��Ի�rND=b�]�"�Ҿ��վt�� �Ѿ�!��%3���>�Z�=�$��E ��K75��P׽��{> ��?��{�\RX�tH���>Ɗ�>:�%=di������}���=-�#?G~>?;����侗�==7۽��>��L?]��=W�������Cƫ>�(?T�>#�=>+��P���:�I�=B�?��?�E?���<Z�3������h �=I�E?
+�>[���O~�Z�`���;?R�0?;�L>�a�vN���!X��?���?Xݓ�d�G>g�2?iw?�?_�6Hq�o"a�?)-��>/���?D��
X�/����y������D�>�P�>M�ľ������>|�����Y�avt�=-�~e��TG�=�,?E���F�=%�>���>�8 ��C�����jn���B3?�ǯ?��?l�=?�¾k���W�ɣ1=�v�>�q�>G��= ��-�>���>�賾�����0	�>��?�3�?VDW?�\j��_Ϳ���1��0Ѿ��<��ǻ3P�=��J�)� >z#>���=3>C�q>OLz>� �=/�=ɨ�<�x�=0"�=�����"�8������~�O�?\/��H����pN������T��Q椾!9t��'g���'�;�Z�	���s��L�D?��N[���'?n��>Ew�>}�=��i=��&��C����=:�����*�Ir�����z�� �׼Fvy����ڡ��߽0��=?Z�1>&sX>1'.?B��=�,)>(��=
�Q=b�>I��>���=�!>
X>w{>�>��d>�<(>ٗ(=�1��uO����7��mE�Q�*��nA?fP����Z�0��L��Xo��I>�g�>Y$>?�2�H����o����>��:xT���T������̓>l�>#^>i�뼟���l�E�����Ff:p/u>d��=K��;_�K�z1��8V=� �>[����=)5�>��U?=d�?�6:?⛵���o>���={7H>q=7�>�> �>2|�>��?;��>�Ŷ>mm�=���X,C��դ�,2�ڇ�=R���/=����=�8>�#�<�7X�0P��l���������Yn��]�����>1�:?)��>�7-?�,��(o�m�R�w���#��>ٶ�x'�>x�-�TԀ>�W�>Y�>�>"�>q���D>/��>��>J2W�#�3����=d
>ʋe=�?�i?Y�Ѿ�-���>b��%����>��?�I�=�����=j��,Lܿ�$�o&�!���LA>R0�<�)���_����=6p4=H9��	~>sn�=-��=���=�\8���2���]>Q��>��A>��\=�/�=�;�=,P0����=��j�ַ��W�9����D�7�����=�S>i^�=�|=C��b���?P.?�H�=`�=j�x�g����1����v>\�>�F�>�P�>M�>-!׾
`�k���x��U�?�X�??��>��W�tq"=�>�>�|�>Ԉ{>%+�=��4�Bٿ��{R����[>�?o�?4bB��73��u>�ׄ��0~�>+��=GkA���?Pb?־��B�ڰ-���2�cC@�~��>�B;�T��X���׾_J��I���p>���;qe�>=ѧ?���>�U�TD����g�O���o�<��~�{�?�i:=Z���|̲�E������#Q��L�=���>�xG>�RL>|�>�U ?(�?��/?i/?��B���?�^�C�>6�>��?4��>k�?���>DR�=��������˽���x ��
۽jN�<�N>0V>��%=���=uM�=~M1�|�?=9�`=�ӽ��/�[��<�T�<Jc�=�?�=�
?y<?���=#�>�[���U�J}�����o�>��;��y����=)ě�l��>!)?zx�>:Q�>  ���?<=ǀ˾���[?D�?ل.>�P��+�>�پ�򖾙(�>�C=�.�}�;Aڬ�g#��o��m�p>�,�>�c��Hj>��~?C?<W#?���J�-��Nr�[�+�ۉżWl�f¬>s��>��=�Ӿ�O5��)s��]�/C-���&�w�I����<:��=ى>��Q>d��=N">)�=������;'dC�Rг>�"�>^�?Q�\>o��=R첾%� ���5?h^M��ž�����۾u^¾�>�W�>� ��_�&?���<�d��m���L�|��>�b�?�V�?�Y?5_žn��Y֔���>Fi�>6x>��.�i�˼x���l>�e�>�$��-����	���>���>؃l>,:�����̇^=�Z��Oi\� ��������J�$žZɱ�t�$�#NR�0��=D	�xbZ��H��c�tp�����H'�p�:�!��)<�?��?7��=�W�N���#��G��BD�>��b��������Ȅ�=����󾖶ԾW���$�Z���b������Y��D��#Ѕ�'���	���=�?�������t�(R>���>6Q�c�8�Tz��T������?��;?q��Jݺ�p��kr��(?���>��?BL���u>�� ?�?U"U��[�Pcm��_�>��?:��?7`6?�9��HZ��+�)PL�3p?R�2?J�<?�	k�sT�(�^��"?#!�>���=D���*��8��y�>^�>��]�>��>A�~>{@I�G���ֿ�j�0�b��=��>4���2�V�����kB��^[>�>��>��[��*�� �>� ݾ�N�`�K��O����#�_=�h?�y�>�MF>$#>��'�j���r��c3��mF?$�?��G?�E4?�S꾒u���z���uY=�ބ>�1�>���=�$E���>j�>������k�)�?�t�?~�?��X?�{g��߿�����7���Nƾm��=>m�v�:>U��S��<�!l=NV�<���-)��qB>Vn�=T�;�?���=$�6>����	)��
������:X��f1�u$��O�$g����L����Q�ѾŴ��a��ὗ�T��	+�}콣��K0�l��=��?6<�>>;�>�Cg>5�>B���5��aw�`ҿ��<�V��b��\bb��l%��ӊ���Iɀ��4��+����>X���)9�>3_+?��=ӂ>2:>�1z�~(���=d5�=^>�=p�>�>a����=�U>�I}>B��=�y���ς�K'8�M�5�����l"A?:gQ�9㈾�8��$۾�_��Q�>�a�>H�L>�o"��M��x���>(���m�ۥ���_��;��>���>��>KK����^���m��MĽ��>��z>1|�=����Ə�K��vT?=�=�>�R��%=`me>�G;?2�?U�? �K>��L>M)m>�0�>ޡ��iV>�v>��%>���>�O ?�?�9�>��=�"�ǳ�>v/b>N���҄��>߽�"`�����T����_�>�0l>���h���RA����#���=��= <�>�NO?���>>��>��x��d4��uc�Jz�à�<P��;N�>���>��a>�2�>�W�>V��>��>?	5=�@>��>>�U>tQI�6��<���>�t>T0H?kA?]]�;"r�qT�����=��==�>>z��>��>GN��Zx���a�޿6��w�l���0=���J
>�* >l)<u:I=5�Ƽy$��2�����պ _#>���<��<l�s��n�����>��@>ߢ�=�U�=N�=�Q�=.v��e�-=�[�f��=�ּL�g���V��M����m�=4Q=g�۽î�;3@	?I�?�<T�[���=�^[پ����(>��>���=S�>aſ>>��1�q�r�/�;�<�C)?�X?X.&?Ǥ	�/ �=�k��!�<��>Dcn>��<>d[�H؞<캠�	��p�>O��>��>�v�=�O=�5l�EKھ���>Z��=�$̽�ݣ?&a?�\�7��S�"��P�h5N��<�9���=0�\�Iv&�Ѣ��?-�t�{�j`���������=�T�>5ݥ?k!�� ~�=jϾ��z8m�_���{�<j�:�I ?�3�>��Q��[;\=�q߀�S�=bΎ<���>��=��>��?A! ?0�3?0��>�y?0>��&?��=>Y�>R�L>@'�>1[?� ?��>�=��<y�;�����敾�[*<E�����=z=O>�~+>=���<1�r�$큼ehҽ��\;R#�=d�t�A�<*S�<��>�%>�L?�?�m.>��]>pᨾ_
�a����ȼeû�L�>�p��S�=ۆ�l�>��E?�ݠ>�k>:������NѾ??7��*?r"?xv�>��n=�G�=��V��u�P>{�>v�����%��ɽ�U'�/�M�z|�=摕>H��<�&u>��z?�hA?�r%?�a�f2�Gb�6�0���<S=P�>��>9C�=K�þm��D�k�]�^���)��p���F��Q<w��=��>��;>���=��>|�<iI��;K���;*@6��+�>&�>%��>)�G>v�D=J�����>I?i.��]��\��h0վ��J��)>%�D>";�u�?,��}aw����L�<��,�>�?o��?׍c?e�M������S>��`>�k)>,�<�B�h$�湗�E�!>z��=X�q�1ʗ� <�X>��~>�˽�fž���a��ݶ�X�9�i�����4�B�醛��u��wnӽ�]���¨=�� �t���'쁾F����ͽ��}��	۾n��a�?E�?�A	;7M¾���Pq�y�:��L#=I)�K�]=��#����Y����Xm���Z>�#��΁y��ؾ���>%!�0���^��������=�oP>��?�����x��&��Q�<0Xi>^���H.�K�v�߂m�?;�<?�"?��=?3��O>'�>Fڗ��w?n-�>�ͪ>�$ݾ�"f�us�>18?asH?Ms����S���?�=U��?��?�&?*�m��Op����y:>H�R?�c?��C?�8>2��7zV����>3�\?��>�".�xo���2�-�7>�+�>f`�	��=��>�g�>m�3�����82=;����=��e>�[�=���=�󥾃v���dO>f�>&C��$W����
��>ᾈ�N�O3@�y����ϡ�{A�=���>Y>�'M>���>m�>:v+�'E��7���Gv�g|3?p}�?�s;?�M$?�$ҾS��z9>��>�	�>V·=�@�HZ�>+x�>{:��C�y�T@��� ?�
�?��?�?1`���ο�����!��̶�b�>�:�= �V>�z���=_ �=tT�<����Dcc=4ۉ>���>�:�>��S>@�>C�=���@)��]������uk=�8��Է	�;�b��&�7�\�E�];��m�ݾ�ϝ�����=��gG�
[���t���F��3��=C$?���>�jw>1B=3�=�Ƥ�ô��y|ξ��T��������*���R����x�w���������I%?.�>>q��=$.?{�޽�&����><佝
>#LJ>�j�=�	�=�_>13�>a��!w̼�N>���>�!�<{́�U�g�&Ǿ{��)y>kL?���0����C��_�����>��>�?v�>�D�qz��}%c��'�>̍���=Ѿ�����ýE�!>�k>t��f>�	F�=��3�7�s�;X�=�F�>�|<>nT,��ݾ������>|�>�������=�0j>��?��U?�n&?��>-ۿ>�Y>���>�;=�*>��3>' u>*�?t�.?Q�?��>�ѿ=�m��7�=�X�=�Yp���Y����N�Ȼ: ��M���t���ﻈ=|e�=#�X=Á�=��=�0���<c5=#�>�U?���>� �>��>==�x'^�ҲӾ�`�>T��<���>9��U�==���>6#?]�>1�>M�g���S�6��>X~o>kF��J`����,\>W_�>��4?{��>J�_�rB|�j���U�=�0�>�I>�vz>Ũ�>*���s�9�L���?m@�#��[���m=�=&>I�8=,Q�=�R�=Xl��W5�>��<��2=B��>ܰ�>&�UB-�r���>(U>`�=���>U�@�.>x�K�y�轏	>?|>��A���=v}4>��}�g�㽜��=s	�ò.>j��<%� ?&?nG�c=P�9^�zо�Dľ֊�>�`�>y��>+ϵ>m_��oH־�$��*��Q�M�?nM?G@�>�>����`;�y/�'+v�Ν>u��>ˮ>3�>K�I#�g��� $�>F�2?8�>G����C�V�i��jξ�v{>�-j=Ύ���?E>|?��%�޲>��v4�ieI�7&�M�+��Ps��=�il��W�)J�>���
�ыν�Y�=���>
0�?�Y�<Z?>�w>������咿����{�<I��,�?ֳ)>	H׽�HO�_�۾�q�e�<;�9� >{!>w�>$,?�� ?t�S?J�Y>K�&>����><;��<v�>'�>��>�B?`��>{"�> �?4��<���=�=�CϞ���1�]J����
>��>�LL>��<�ʰ=(�=�l=�U[=	Å���_=��B�2�P�=1Y<>�ݶ��W?��?��=��[>��ྉ�۾0r=<%O>z��=. ܽ��t��y=X�=�g�>s��>_��>ӂu�Y^�� ����Z����?��>5�>�=�='�>M��줅��> du>��f=��Ӿee���ʢ=�d�<��=��=}�����>��u?F>?��&?0&�xC+�ߠU�5m'��^b� �ȼ?��>�a�>=8=&WϾ�E�v�`���_��,�m�&�sS���u<n�=Z��=}?�>�f
>؀@>
�;�7�N��K�.��V^=� �>���>�G?(C�=}�5=�泾*����C?_����X��韾�TľX�h��}">ȫv>�^��A? 2ݽ,
o�L.��jgC��T�>�ֿ??i�?S�Y?��J�mT!���/>���>~#>�]=!�-��ן��.:��l>���=��������(�2���a>I��>��D�=D��u+徼���Y����?��;��n��\�*O��ޏ��u@#���<��U>�T��e�)ʪ��5�6#i��=��S�	���Z��\��?)԰?v}w>�:��	@���W�B�d^��?�����=R ̾���>�Q�sܰ=��Z�?��}�[Ӿ���y��>a�<�jȒ�VYh�;�Ӿhl>�5�>Ƴ�>�����?�3d�(	����>S~>����A�������������U?R�!?�R�2꾨dJ=T��1�?2 �>�^>� x��o���6��i�N?��a?֪&=ˊ����:�-;�
�?*��?�W2?���&PP��ؾ���;K?fn<? ?�_����޾������>ˮF?q��=o�c��6�����N�>3,?�;L��i	=(? n�>#�����f�\�O�>����(�=�ak>�\{���Ҿy����2�ϭ�>���>-=Ս۾��>|�����Y�avt�=-�~e��TG�=�,?E���F�=%�>���>�8 ��C�����jn���B3?�ǯ?��?l�=?�¾k���W�ɣ1=�v�>�q�>G��= ��-�>���>�賾�����0	�>��?�3�?VDW?�\j��_Ϳ���1��0Ѿ��<��ǻ3P�=��J�)� >z#>���=3>C�q>OLz>� �=/�=ɨ�<�x�=0"�=�����"�8������~�O�?\/��H����pN������T��Q椾!9t��'g���'�;�Z�	���s��L�D?��N[���'?n��>Ew�>}�=��i=��&��C����=:�����*�Ir�����z�� �׼Fvy����ڡ��߽0��=?Z�1>&sX>1'.?B��=�,)>(��=
�Q=b�>I��>���=�!>
X>w{>�>��d>�<(>ٗ(=�1��uO����7��mE�Q�*��nA?fP����Z�0��L��Xo��I>�g�>Y$>?�2�H����o����>��:xT���T������̓>l�>#^>i�뼟���l�E�����Ff:p/u>d��=K��;_�K�z1��8V=� �>[����=)5�>��U?=d�?�6:?⛵���o>���={7H>q=7�>�> �>2|�>��?;��>�Ŷ>mm�=���X,C��դ�,2�ڇ�=R���/=����=�8>�#�<�7X�0P��l���������Yn��]�����>1�:?)��>�7-?�,��(o�m�R�w���#��>ٶ�x'�>x�-�TԀ>�W�>Y�>�>"�>q���D>/��>��>J2W�#�3����=d
>ʋe=�?�i?Y�Ѿ�-���>b��%����>��?�I�=�����=j��,Lܿ�$�o&�!���LA>R0�<�)���_����=6p4=H9��	~>sn�=-��=���=�\8���2���]>Q��>��A>��\=�/�=�;�=,P0����=��j�ַ��W�9����D�7�����=�S>i^�=�|=C��b���?P.?�H�=`�=j�x�g����1����v>\�>�F�>�P�>M�>-!׾
`�k���x��U�?�X�??��>��W�tq"=�>�>�|�>Ԉ{>%+�=��4�Bٿ��{R����[>�?o�?4bB��73��u>�ׄ��0~�>+��=GkA���?Pb?־��B�ڰ-���2�cC@�~��>�B;�T��X���׾_J��I���p>���;qe�>=ѧ?���>�U�TD����g�O���o�<��~�{�?�i:=Z���|̲�E������#Q��L�=���>�xG>�RL>|�>�U ?(�?��/?i/?��B���?�^�C�>6�>��?4��>k�?���>DR�=��������˽���x ��
۽jN�<�N>0V>��%=���=uM�=~M1�|�?=9�`=�ӽ��/�[��<�T�<Jc�=�?�=�
?y<?���=#�>�[���U�J}�����o�>��;��y����=)ě�l��>!)?zx�>:Q�>  ���?<=ǀ˾���[?D�?ل.>�P��+�>�پ�򖾙(�>�C=�.�}�;Aڬ�g#��o��m�p>�,�>�c��Hj>��~?C?<W#?���J�-��Nr�[�+�ۉżWl�f¬>s��>��=�Ӿ�O5��)s��]�/C-���&�w�I����<:��=ى>��Q>d��=N">)�=������;'dC�Rг>�"�>^�?Q�\>o��=R첾%� ���5?h^M��ž�����۾u^¾�>�W�>� ��_�&?���<�d��m���L�|��>�b�?�V�?�Y?5_žn��Y֔���>Fi�>6x>��.�i�˼x���l>�e�>�$��-����	���>���>؃l>,:�����̇^=�Z��Oi\� ��������J�$žZɱ�t�$�#NR�0��=D	�xbZ��H��c�tp�����H'�p�:�!��)<�?��?7��=�W�N���#��G��BD�>��b��������Ȅ�=����󾖶ԾW���$�Z���b������Y��D��#Ѕ�'���	���=�?�������t�(R>���>6Q�c�8�Tz��T������?��;?q��Jݺ�p��kr��(?���>��?BL���u>�� ?�?U"U��[�Pcm��_�>��?:��?7`6?�9��HZ��+�)PL�3p?R�2?J�<?�	k�sT�(�^��"?#!�>���=D���*��8��y�>^�>��]�>��>A�~>{@I�G���ֿ�j�0�b��=��>4���2�V�����kB��^[>�>��>��[��*�� �>� ݾ�N�`�K��O����#�_=�h?�y�>�MF>$#>��'�j���r��c3��mF?$�?��G?�E4?�S꾒u���z���uY=�ބ>�1�>���=�$E���>j�>������k�)�?�t�?~�?��X?�{g��߿�����7���Nƾm��=>m�v�:>U��S��<�!l=NV�<���-)��qB>Vn�=T�;�?���=$�6>����	)��
������:X��f1�u$��O�$g����L����Q�ѾŴ��a��ὗ�T��	+�}콣��K0�l��=��?6<�>>;�>�Cg>5�>B���5��aw�`ҿ��<�V��b��\bb��l%��ӊ���Iɀ��4��+����>X���)9�>3_+?��=ӂ>2:>�1z�~(���=d5�=^>�=p�>�>a����=�U>�I}>B��=�y���ς�K'8�M�5�����l"A?:gQ�9㈾�8��$۾�_��Q�>�a�>H�L>�o"��M��x���>(���m�ۥ���_��;��>���>��>KK����^���m��MĽ��>��z>1|�=����Ə�K��vT?=�=�>�R��%=`me>�G;?2�?U�? �K>��L>M)m>�0�>ޡ��iV>�v>��%>���>�O ?�?�9�>��=�"�ǳ�>v/b>N���҄��>߽�"`�����T����_�>�0l>���h���RA����#���=��= <�>�NO?���>>��>��x��d4��uc�Jz�à�<P��;N�>���>��a>�2�>�W�>V��>��>?	5=�@>��>>�U>tQI�6��<���>�t>T0H?kA?]]�;"r�qT�����=��==�>>z��>��>GN��Zx���a�޿6��w�l���0=���J
>�* >l)<u:I=5�Ƽy$��2�����պ _#>���<��<l�s��n�����>��@>ߢ�=�U�=N�=�Q�=.v��e�-=�[�f��=�ּL�g���V��M����m�=4Q=g�۽î�;3@	?I�?�<T�[���=�^[پ����(>��>���=S�>aſ>>��1�q�r�/�;�<�C)?�X?X.&?Ǥ	�/ �=�k��!�<��>Dcn>��<>d[�H؞<캠�	��p�>O��>��>�v�=�O=�5l�EKھ���>Z��=�$̽�ݣ?&a?�\�7��S�"��P�h5N��<�9���=0�\�Iv&�Ѣ��?-�t�{�j`���������=�T�>5ݥ?k!�� ~�=jϾ��z8m�_���{�<j�:�I ?�3�>��Q��[;\=�q߀�S�=bΎ<���>��=��>��?A! ?0�3?0��>�y?0>��&?��=>Y�>R�L>@'�>1[?� ?��>�=��<y�;�����敾�[*<E�����=z=O>�~+>=���<1�r�$큼ehҽ��\;R#�=d�t�A�<*S�<��>�%>�L?�?�m.>��]>pᨾ_
�a����ȼeû�L�>�p��S�=ۆ�l�>��E?�ݠ>�k>:������NѾ??7��*?r"?xv�>��n=�G�=��V��u�P>{�>v�����%��ɽ�U'�/�M�z|�=摕>H��<�&u>��z?�hA?�r%?�a�f2�Gb�6�0���<S=P�>��>9C�=K�þm��D�k�]�^���)��p���F��Q<w��=��>��;>���=��>|�<iI��;K���;*@6��+�>&�>%��>)�G>v�D=J�����>I?i.��]��\��h0վ��J��)>%�D>";�u�?,��}aw����L�<��,�>�?o��?׍c?e�M������S>��`>�k)>,�<�B�h$�湗�E�!>z��=X�q�1ʗ� <�X>��~>�˽�fž���a��ݶ�X�9�i�����4�B�醛��u��wnӽ�]���¨=�� �t���'쁾F����ͽ��}��	۾n��a�?E�?�A	;7M¾���Pq�y�:��L#=I)�K�]=��#����Y����Xm���Z>�#��΁y��ؾ���>%!�0���^��������=�oP>��?�����x��&��Q�<0Xi>^���H.�K�v�߂m�?;�<?�"?��=?3��O>'�>Fڗ��w?n-�>�ͪ>�$ݾ�"f�us�>18?asH?Ms����S���?�=U��?��?�&?*�m��Op����y:>H�R?�c?��C?�8>2��7zV����>3�\?��>�".�xo���2�-�7>�+�>f`�	��=��>�g�>m�3�����82=;����=��e>�[�=���=�󥾃v���dO>f�>&C��$W����G�>�}꾹N� �G��������<M�?Rr�T>+�f>�>�E(�|����Y��e��PL?G�?\�S?�7?�.��񾅔��S�=�>�7�>�,�=������>V4�>* 辭�p�<���?@ �?@��?��Z?v,l���ؿw?����ʾ}�׾(@�Q�=7>#��IA�=��`uԽKȽ��!>��>���>z'>	�,>#�/>&�>@T����'��5�����J^��V��۾��������nB��о�I��q·<�>�:����K��D����5=����t�(>33M?�� ?��>�]�><&^>XLȾ�p&�C��w齴��:�ɾ��4���3���1��o��+~�����2�a�J�3��0�>������>��?έ�<1�>��>X,�Q5� ��=Ó���<�zI>f>�gJ>XZ�>x�?�+�>h#�>�����:��缽�z����*@�?�i�Ӣ�"�b�{�����-�}��>�]-� �.>&^a��������z��>�2U���C�p>Z��Z��C��>4� =Ro��m>31�k���D�x=���>��.>�Ⱦ�~����]��ž�A�>	���H�� N���G?��?�hn?8���)>I=P5����>��r>��>J�>�&d>�U�> �?�>�?�-l? �=�~½�p���	��P�I����B������%��G�=�:=h5=E# >S�=��<�J��+:>�]N=[O=f�?�_?��>�?w"�<<ဿ��M���>���>�D?{�5?��=(��>�'�>��G?��z>QXg=�ܾ<WϾ���>p��>9�<�	�{����=J#V>(�>�9�\?�ri?C��^����=t��z�=���>���>j�v>'}z>�&>�,��a޿�7�P� ��&,��8�=4YE�w�8��G��?S8������b>�_�>q�?z�!>C�Z>:��>O��>sI�>�G4>�[>Hc:>�Uo=!��s
�m�w=���<����l���t�<c�H�����@4�6��?w{��U����Z�, ?��"?]=�W�=��󽦜����#�s)?(�?r_E? \�>ds�#4���:�3�����:[��>z#Q?}� ?9�V�L˼��E>���>���>��>��Q>:�Ѿ��ª��ڤ>
��>�4?h��>,3��sK��Dz�`(�-I�=�1�=�v_��;�?�b?���>[�:��;�����7��#��YN�=\hg=(C�*E{�K~������H3��@���RJ��4�>�J�?	 `�h}�=B�[��勿6�=�'џ�EF>��=']�>~͡>���<}J�,p�5��iѽ���=�V�>��=���>;�?ZO?�`?!?N5?�X^���>1��=���>�Ъ>ޫ?�?���>N��>}�>�w�=d5�<���<����<�k&����= �=/�=��b=��=�8�<$~�<������ɼ�Τ�)�м��U=L��=ӵ=��=
�
?�{=?�.x=��z>2��=�.��W�=w7�=)v�<xi>=�9>j��&>�~�>�`?���>J�<!ھRR;�0㾢�
��c?4�;?��>XU�=s��>��׾�Խ����>�y�>�eǾwtھ�Ӿ�������<��>l��=�"#>�͋>�~~?��I?tx.?��I�����-u��M��L}�����1?)�:?�,?�Q�/u���,�Y����a�ɾ�eν�|>CB��4U<���>�V$�D�>�ۑ��_5��-���S>��=}�> _�>��>��X=�>@Y��U�{��4L?"�I�F]�>���?��'Wཞ�=#�>�I�=�.?����y��9I���8�f�>���?:��?�Y?(Q�E���G>"�4>��>�q�&���=0W�<'� >>G/~����'e��p/>�h>��ҽ/���1l��z��<踱��H����iT��xƽ|آ����ME�=�L�<�����"����^G����j��h����2��麽U�����=�f �?��?�1�k��� �r�I�Ѿ���8�>X]�<�-�D*���/=�����v�������(�V�+��B����GY�>Ԏ��n��^pg�X�1V�kx>Ͻ"?O�����x���������t�=f�=8��gk��_+��;���(?<�?]����:�j�}�_�=3+?w�y>��(�s��2�<ˮ>��,?�3?��`��t�b�������`�?50�?��??S�#=��Y�&��Q?��?���>&Ǒ���Ⱦ���7?�R<?Lc�>d��~���h����>�Z?<%G���O>��>|S�>u&�
��azh�+	��O�+��s7>]�^:���^�W�6��9�=٫�>/ۀ>�aS������u�>��L%N��WH�Ç�HP���<o?�	�#�>�Ve>�>Xb)��쌿!\�����wL?F��?�ES?n�7?b���,��������=>ץ>���>B�=�	��1�>}>�>Ӫ��s�,���i?���?�N�?��Z?��k���п]���� ���̾��=;�=XϽ>��f���)e�<ud7<����=me>��=]4P=���>�0x>��K>�Ą�,�%�k��	����R3���U���N�n��)|���>���׾k��� sJ��T.��u�O���hb�+_s=ۃ�<% �G�*?�q�>�|�={��>ǘ>��~���Ͼ�'����1�]�_�ۦ'�_\4�x�H��v0�/�*��j}��ؿ�o���6�.�?^��<Д�>�,?�e�=�m>4�>�Eս��>��H<t�l>�'��U̼��s>-�>I�?��s>Fެ=�E=�Z��LGm�z����zѧ���|?�
6���`����SWĽ8� ��h�>p�>��,>�G������؅����>r������2%4=�ľ��6>�?�,��I�㻨��=�c�*��b�ἣ�~>=�={�~�vז�Ɲ��.r?�n�.?%s��/�<S`>.�
?Û{?Rz3?���O�>��>d��>�A�=��W<�g�>`0*?T�2?�+?��a?Ѹ@?#�1=�ye��:v>�e>����սT�����8<}^��W��=�0�=EQ�<EB�=`}E;:��=��?<��3>M��<���3�>-�a?���>&��>hm�<�p@��QK�H����c=b��:��>�-?(?�e>t]�>Ut>�bk���徳ϱ�/a�>>��>۫w��J��h�n>?�>$[��,� ?3]s??W/�6`ܾ���>6L߽�w�>!\�>%�>Q��>@�B>�c�>b���zԿ�W���I���ٽģJ�j��=*�ʃ]��=�����v����>���>Fќ>�)>�L>��>?�>��>-�->'��=~˾=�W3=`�j��ps����=���=�ج=�Ҫ<��>��=/8c��I=�q>��d�� ������?�?�!"��1�*F����U���NU�>���>-�>�]�>�|�=���?J��=6�O�
���?�]?U?�D����=��<��=���>�ٙ>�$>����G��?<�� =x�>��#?6��>��-��U�o'b�5��9��>	=="2���?��J?"%�}+�;��<�j�0�i������&��=�����o�:`��L6��J�UD�EI�����>�p�?gPe�7�j=zj��ƚ�%���[�������g�S� ?���>��P>��_��O����0=��-��Ab��O��E>�^�>Py?)�+?	�^?ݿ�>��>`s��M��>;�>t��>Ɛ�>�k?��?�9�>�g9>�w�>�����^�;�\�f�g�E�<� Ҽ�c�=m�>ޣn>�Qq=��n=�LP<��9a��vm���������R�<��<Ó1>��U=�p?�1/?w�� ���㸻x(P�G�ɼH�,���>_���(�9���Z=6e>�B�>�n?�~�>���=�đ�o�Q�/�Ͼ�.��e'�>�O?�ؼ>>��>�(޾�D��dcd>FD�>l�$�ʬ��@�w�z~���/Z�-I>�|�>7�k>�.a>5vp?1M? �V?�
��(��7C��I��A�-��<?�>�q]>8��Z# � �O��=3���/����S;��s)=�~�=�y�>c�>����M��>��;�)���K�=B�N<��뼭ҷ>�=�>Em�>c�=>˔�=U������L?����0�al�����qx�J�!>D&�><�{����>���s(r�?����>��\�>���?���?F�b?��	�_��P�E>�>c�@>fZ���U]�ʨ^��ֽ��>P�0>�]�i���,�=�bu>H>Yt��M���r⾡�������b?������i��y��h��uc߾�b�=U�n��0��	��œ=aUY�1�l����$F�=I޾V����=f�5��?V'�?Q<>�GĽT3���,��$ ���]>�+پ�8���{7��{^��������=�_��� ��+&��2B�1�>�}C�-���~sh��B�(>�=�2>2�?�ξ�Ǘ�aE3��P��ZB=�q�<�F���W��_���T�p�Uj5?��?�r	��i��d����ю>�.?���>~�5>=��x���i�>�!?��&?�V-�i������px�=�ݽ?�d�?�C?����x<�����x�B�?���>��>&.$���ݾT���(?�'(?|��>�����w�O �)X�>}\?]KC�GmC>�)�>W�>3��+���K=;�6�kE���=��<=&��Q���\���?>�Y�>C�i>ƍ�����G�>�}꾹N� �G��������<M�?Rr�T>+�f>�>�E(�|����Y��e��PL?G�?\�S?�7?�.��񾅔��S�=�>�7�>�,�=������>V4�>* 辭�p�<���?@ �?@��?��Z?v,l���ؿw?����ʾ}�׾(@�Q�=7>#��IA�=��`uԽKȽ��!>��>���>z'>	�,>#�/>&�>@T����'��5�����J^��V��۾��������nB��о�I��q·<�>�:����K��D����5=����t�(>33M?�� ?��>�]�><&^>XLȾ�p&�C��w齴��:�ɾ��4���3���1��o��+~�����2�a�J�3��0�>������>��?έ�<1�>��>X,�Q5� ��=Ó���<�zI>f>�gJ>XZ�>x�?�+�>h#�>�����:��缽�z����*@�?�i�Ӣ�"�b�{�����-�}��>�]-� �.>&^a��������z��>�2U���C�p>Z��Z��C��>4� =Ro��m>31�k���D�x=���>��.>�Ⱦ�~����]��ž�A�>	���H�� N���G?��?�hn?8���)>I=P5����>��r>��>J�>�&d>�U�> �?�>�?�-l? �=�~½�p���	��P�I����B������%��G�=�:=h5=E# >S�=��<�J��+:>�]N=[O=f�?�_?��>�?w"�<<ဿ��M���>���>�D?{�5?��=(��>�'�>��G?��z>QXg=�ܾ<WϾ���>p��>9�<�	�{����=J#V>(�>�9�\?�ri?C��^����=t��z�=���>���>j�v>'}z>�&>�,��a޿�7�P� ��&,��8�=4YE�w�8��G��?S8������b>�_�>q�?z�!>C�Z>:��>O��>sI�>�G4>�[>Hc:>�Uo=!��s
�m�w=���<����l���t�<c�H�����@4�6��?w{��U����Z�, ?��"?]=�W�=��󽦜����#�s)?(�?r_E? \�>ds�#4���:�3�����:[��>z#Q?}� ?9�V�L˼��E>���>���>��>��Q>:�Ѿ��ª��ڤ>
��>�4?h��>,3��sK��Dz�`(�-I�=�1�=�v_��;�?�b?���>[�:��;�����7��#��YN�=\hg=(C�*E{�K~������H3��@���RJ��4�>�J�?	 `�h}�=B�[��勿6�=�'џ�EF>��=']�>~͡>���<}J�,p�5��iѽ���=�V�>��=���>;�?ZO?�`?!?N5?�X^���>1��=���>�Ъ>ޫ?�?���>N��>}�>�w�=d5�<���<����<�k&����= �=/�=��b=��=�8�<$~�<������ɼ�Τ�)�м��U=L��=ӵ=��=
�
?�{=?�.x=��z>2��=�.��W�=w7�=)v�<xi>=�9>j��&>�~�>�`?���>J�<!ھRR;�0㾢�
��c?4�;?��>XU�=s��>��׾�Խ����>�y�>�eǾwtھ�Ӿ�������<��>l��=�"#>�͋>�~~?��I?tx.?��I�����-u��M��L}�����1?)�:?�,?�Q�/u���,�Y����a�ɾ�eν�|>CB��4U<���>�V$�D�>�ۑ��_5��-���S>��=}�> _�>��>��X=�>@Y��U�{��4L?"�I�F]�>���?��'Wཞ�=#�>�I�=�.?����y��9I���8�f�>���?:��?�Y?(Q�E���G>"�4>��>�q�&���=0W�<'� >>G/~����'e��p/>�h>��ҽ/���1l��z��<踱��H����iT��xƽ|آ����ME�=�L�<�����"����^G����j��h����2��麽U�����=�f �?��?�1�k��� �r�I�Ѿ���8�>X]�<�-�D*���/=�����v�������(�V�+��B����GY�>Ԏ��n��^pg�X�1V�kx>Ͻ"?O�����x���������t�=f�=8��gk��_+��;���(?<�?]����:�j�}�_�=3+?w�y>��(�s��2�<ˮ>��,?�3?��`��t�b�������`�?50�?��??S�#=��Y�&��Q?��?���>&Ǒ���Ⱦ���7?�R<?Lc�>d��~���h����>�Z?<%G���O>��>|S�>u&�
��azh�+	��O�+��s7>]�^:���^�W�6��9�=٫�>/ۀ>�aS�����G�>�}꾹N� �G��������<M�?Rr�T>+�f>�>�E(�|����Y��e��PL?G�?\�S?�7?�.��񾅔��S�=�>�7�>�,�=������>V4�>* 辭�p�<���?@ �?@��?��Z?v,l���ؿw?����ʾ}�׾(@�Q�=7>#��IA�=��`uԽKȽ��!>��>���>z'>	�,>#�/>&�>@T����'��5�����J^��V��۾��������nB��о�I��q·<�>�:����K��D����5=����t�(>33M?�� ?��>�]�><&^>XLȾ�p&�C��w齴��:�ɾ��4���3���1��o��+~�����2�a�J�3��0�>������>��?έ�<1�>��>X,�Q5� ��=Ó���<�zI>f>�gJ>XZ�>x�?�+�>h#�>�����:��缽�z����*@�?�i�Ӣ�"�b�{�����-�}��>�]-� �.>&^a��������z��>�2U���C�p>Z��Z��C��>4� =Ro��m>31�k���D�x=���>��.>�Ⱦ�~����]��ž�A�>	���H�� N���G?��?�hn?8���)>I=P5����>��r>��>J�>�&d>�U�> �?�>�?�-l? �=�~½�p���	��P�I����B������%��G�=�:=h5=E# >S�=��<�J��+:>�]N=[O=f�?�_?��>�?w"�<<ဿ��M���>���>�D?{�5?��=(��>�'�>��G?��z>QXg=�ܾ<WϾ���>p��>9�<�	�{����=J#V>(�>�9�\?�ri?C��^����=t��z�=���>���>j�v>'}z>�&>�,��a޿�7�P� ��&,��8�=4YE�w�8��G��?S8������b>�_�>q�?z�!>C�Z>:��>O��>sI�>�G4>�[>Hc:>�Uo=!��s
�m�w=���<����l���t�<c�H�����@4�6��?w{��U����Z�, ?��"?]=�W�=��󽦜����#�s)?(�?r_E? \�>ds�#4���:�3�����:[��>z#Q?}� ?9�V�L˼��E>���>���>��>��Q>:�Ѿ��ª��ڤ>
��>�4?h��>,3��sK��Dz�`(�-I�=�1�=�v_��;�?�b?���>[�:��;�����7��#��YN�=\hg=(C�*E{�K~������H3��@���RJ��4�>�J�?	 `�h}�=B�[��勿6�=�'џ�EF>��=']�>~͡>���<}J�,p�5��iѽ���=�V�>��=���>;�?ZO?�`?!?N5?�X^���>1��=���>�Ъ>ޫ?�?���>N��>}�>�w�=d5�<���<����<�k&����= �=/�=��b=��=�8�<$~�<������ɼ�Τ�)�м��U=L��=ӵ=��=
�
?�{=?�.x=��z>2��=�.��W�=w7�=)v�<xi>=�9>j��&>�~�>�`?���>J�<!ھRR;�0㾢�
��c?4�;?��>XU�=s��>��׾�Խ����>�y�>�eǾwtھ�Ӿ�������<��>l��=�"#>�͋>�~~?��I?tx.?��I�����-u��M��L}�����1?)�:?�,?�Q�/u���,�Y����a�ɾ�eν�|>CB��4U<���>�V$�D�>�ۑ��_5��-���S>��=}�> _�>��>��X=�>@Y��U�{��4L?"�I�F]�>���?��'Wཞ�=#�>�I�=�.?����y��9I���8�f�>���?:��?�Y?(Q�E���G>"�4>��>�q�&���=0W�<'� >>G/~����'e��p/>�h>��ҽ/���1l��z��<踱��H����iT��xƽ|آ����ME�=�L�<�����"����^G����j��h����2��麽U�����=�f �?��?�1�k��� �r�I�Ѿ���8�>X]�<�-�D*���/=�����v�������(�V�+��B����GY�>Ԏ��n��^pg�X�1V�kx>Ͻ"?O�����x���������t�=f�=8��gk��_+��;���(?<�?]����:�j�}�_�=3+?w�y>��(�s��2�<ˮ>��,?�3?��`��t�b�������`�?50�?��??S�#=��Y�&��Q?��?���>&Ǒ���Ⱦ���7?�R<?Lc�>d��~���h����>�Z?<%G���O>��>|S�>u&�
��azh�+	��O�+��s7>]�^:���^�W�6��9�=٫�>/ۀ>�aS������u�>��L%N��WH�Ç�HP���<o?�	�#�>�Ve>�>Xb)��쌿!\�����wL?F��?�ES?n�7?b���,��������=>ץ>���>B�=�	��1�>}>�>Ӫ��s�,���i?���?�N�?��Z?��k���п]���� ���̾��=;�=XϽ>��f���)e�<ud7<����=me>��=]4P=���>�0x>��K>�Ą�,�%�k��	����R3���U���N�n��)|���>���׾k��� sJ��T.��u�O���hb�+_s=ۃ�<% �G�*?�q�>�|�={��>ǘ>��~���Ͼ�'����1�]�_�ۦ'�_\4�x�H��v0�/�*��j}��ؿ�o���6�.�?^��<Д�>�,?�e�=�m>4�>�Eս��>��H<t�l>�'��U̼��s>-�>I�?��s>Fެ=�E=�Z��LGm�z����zѧ���|?�
6���`����SWĽ8� ��h�>p�>��,>�G������؅����>r������2%4=�ľ��6>�?�,��I�㻨��=�c�*��b�ἣ�~>=�={�~�vז�Ɲ��.r?�n�.?%s��/�<S`>.�
?Û{?Rz3?���O�>��>d��>�A�=��W<�g�>`0*?T�2?�+?��a?Ѹ@?#�1=�ye��:v>�e>����սT�����8<}^��W��=�0�=EQ�<EB�=`}E;:��=��?<��3>M��<���3�>-�a?���>&��>hm�<�p@��QK�H����c=b��:��>�-?(?�e>t]�>Ut>�bk���徳ϱ�/a�>>��>۫w��J��h�n>?�>$[��,� ?3]s??W/�6`ܾ���>6L߽�w�>!\�>%�>Q��>@�B>�c�>b���zԿ�W���I���ٽģJ�j��=*�ʃ]��=�����v����>���>Fќ>�)>�L>��>?�>��>-�->'��=~˾=�W3=`�j��ps����=���=�ج=�Ҫ<��>��=/8c��I=�q>��d�� ������?�?�!"��1�*F����U���NU�>���>-�>�]�>�|�=���?J��=6�O�
���?�]?U?�D����=��<��=���>�ٙ>�$>����G��?<�� =x�>��#?6��>��-��U�o'b�5��9��>	=="2���?��J?"%�}+�;��<�j�0�i������&��=�����o�:`��L6��J�UD�EI�����>�p�?gPe�7�j=zj��ƚ�%���[�������g�S� ?���>��P>��_��O����0=��-��Ab��O��E>�^�>Py?)�+?	�^?ݿ�>��>`s��M��>;�>t��>Ɛ�>�k?��?�9�>�g9>�w�>�����^�;�\�f�g�E�<� Ҽ�c�=m�>ޣn>�Qq=��n=�LP<��9a��vm���������R�<��<Ó1>��U=�p?�1/?w�� ���㸻x(P�G�ɼH�,���>_���(�9���Z=6e>�B�>�n?�~�>���=�đ�o�Q�/�Ͼ�.��e'�>�O?�ؼ>>��>�(޾�D��dcd>FD�>l�$�ʬ��@�w�z~���/Z�-I>�|�>7�k>�.a>5vp?1M? �V?�
��(��7C��I��A�-��<?�>�q]>8��Z# � �O��=3���/����S;��s)=�~�=�y�>c�>����M��>��;�)���K�=B�N<��뼭ҷ>�=�>Em�>c�=>˔�=U������L?����0�al�����qx�J�!>D&�><�{����>���s(r�?����>��\�>���?���?F�b?��	�_��P�E>�>c�@>fZ���U]�ʨ^��ֽ��>P�0>�]�i���,�=�bu>H>Yt��M���r⾡�������b?������i��y��h��uc߾�b�=U�n��0��	��œ=aUY�1�l����$F�=I޾V����=f�5��?V'�?Q<>�GĽT3���,��$ ���]>�+پ�8���{7��{^��������=�_��� ��+&��2B�1�>�}C�-���~sh��B�(>�=�2>2�?�ξ�Ǘ�aE3��P��ZB=�q�<�F���W��_���T�p�Uj5?��?�r	��i��d����ю>�.?���>~�5>=��x���i�>�!?��&?�V-�i������px�=�ݽ?�d�?�C?����x<�����x�B�?���>��>&.$���ݾT���(?�'(?|��>�����w�O �)X�>}\?]KC�GmC>�)�>W�>3��+���K=;�6�kE���=��<=&��Q���\���?>�Y�>C�i>ƍ�������>W��,�P���M������S=yo�>i��~I>c�X>7I>�p,����Z�������CF?�î?�O?0�:?�y��p�Y����<D�{>�d�>���=O����>�T�>a¾��b�4 ���?�9�?�U�?��[?�i�U�ٿ+Х�����f�pR�=���<C�c>hR��z��=���=�N=�螼�:�=,^L>�a>k�>sZ>U�>�E�=M���'�4������$8�A��p���i�� �>�]������Ѿ%�Ӿ��꽓^�=��@i��<�j��f�j�[�sji=�PC?�.�>p�G>����+��>� �`Ȥ�� )���|�������U���i1��G����񾋕���(���8����q	�>���=:��>�0?�;��ca>�y�>���:*C=.o�< �>d�ս�VW>��>q�'>B�>5�>���>���>*�������v[�Q|u�@������?x�>�ɑ�>�����2`>3|���?ʒ?�5;>��0��-��NY���9�>�����~���>a�[�g��<���>��^>���e핽O�'����w>��>�Ā>������r�z�]B�<�\�>%%y�3<=1e�>g8?��G?��d?�ʽ#h�>!�>.�?I���y������ם�>C�d?9�7?NV^?�rJ<̦T�X�ʽ�Y���g��Q�����=�+>���pΫ�������=h�4����Z�	d>�UW����^��=�m�>��>?P��>k1?��P=7^����X��D��{k�>SK����>��>#o9?�a�>���>&��O�=?ך��*����>�$�>�o��	��.�X=@r�>�=i�?6�
?��>~����9��oc>��]>���>���>���>Ȩ�>���=h� ��ʿj{A�n2��b��?=c>�=�(�6б�<1=�ꧽ�P��"�{�RLx���=�Q`>F��=|�==~X�=ny?�X�>0�ڽD2��y����.=q
�a������H�>>0D��d@	=zQ�����:��)=��<Ϡ�6�m=K=�
?�V
?F��Q����n���򄟾�e�>�á>�}?�W�>~ >d	�xfI�rp=����N��>�]?���>N��d�=]�M�<���>͠>��>�@M�Uw������Yٻ�o�>�#	?��>�<�)�O���r�E�� �>h�z=裳��K�?�dH?�|��>_������5��������`>*C��K���Ͼ�ȾL����h+���+�Z�==h�>h�?g����n>oe���ۂ��颿ʖ+�ak#>'��fq?�D�>,���>�ܾ�F^�I�žԐ�=g�#>;߂>�Y	>���>�@?�"N?�Z?3q?���>����?��4����>�1�>� ?��>��?wç>6ظ>�O�=��=���T����sϽǊ'=ݷ�<�?>	k>4*;=n�ܼ�����
�=�.$���������I=���=���=�
���%=Uq?�G#?{��;���<N����z���1��;�����=��Q���l���=C��>�p,?���>��=/=��lv���L��Y[��.ā���b?x�^?�>��)�>�>�����3=�ݗ>(�����H��r ��(m���E>�U�>*��=�[�>��?�\?�8?+/8>�����n�|�"�_ �>�� X�>{�>+P?�M��$�+�(W�O5�����d���q��'뽊t0>_R�=��!>~��>eUz>���=��>7L=����(>��><�?��:?Vf4>)�$>Ą��W�ξp�G?�ˢ�r�����>�Ͼ-?�>e89>�l�ג?[$��z�Ω��]B=��d�>��?0%�?jNc?l�7�ya���5[>�+T>��>�*�<��;�^�+��{��;/>�[�=?�}�;����ĺ�R]>I-u>�2Ľ�4;|����S�4F��ϩ-�^�ҾZ�%�vo��S��ɾtj���?>���B�:�	��杽c�R�)oL���U��z/��}�.$�?��?BD>�r�`j�����LK � x�>6�t��8�Y���Ny���$�����
O����
�h<�o�
���$��,�>�)
�������q�>bL���:��uD>�B?�v�����|�o��=�r�=v��=	��:ꍿ]���1S��*0?۫?�i�A����c�<A�=�V�>K��>Ȃ����������>z?
?3�.?�j��ה��l���ż7��?s�?�A? x̽��6�HC����&5�>ŧ�>?�>
�x�𪩾�P4����>�4?���>Ѱ�tχ�
[���>�CN?
l^��'J>�T�>dy�>>Ӽ�t��a�=e��܃���Z>�wK<_�Q��vw��;
�Y����r�>���>i�m�����^į>;���N�n`I�,���"����<)� ?w��>z�}>i�
>X3'�^%��I������u/L?n_�?��V?�7?7�ӈ��޽�q%=�z�>"�>�0�=���ũ>^��>	쾥r������?���?���?K�R?'�g���Կ�d���н�YK���0�=�'">7�`>�P�Y=�� d�����g=y��>k+>�@o>Hʡ>d�>��|>�V����+�n������{��@M�8��cTT��#�3��<��f��[��ĕA�"��fG����N�����<�u�a�1��=�� ?�>���>]]L>�O�>&"S��H���'z�=[J���N�X���q[ݾ�)������>��E������٥�F�>𨵽m(>J��>��9���G=z��>^2>�nH>W��>)�>v�7>ҳ�>V��>R��=7̡>�#�;Z��>��]>�ϋ��V=�iht�s����f?2��T�>�ڌ���)��̾O]�>�M�>��<`�O�WS���#l����>�&��难�H��@X��~!>m �>�`�>�����o=2�ɽK��=��M>	Ơ>�P>:���ϰ��Ј<�v>w��>�@���ܼ=���>��;?�{?A?�-�b�>��̽�=��E�v;�<r�=���z>�B;?�%I?��9?�7�>���=�����\H��pýg-��ը���м G������>�{����<d� =���<��>k>��`=��$>tZ�>[��>��[?Po?Cu?�
>�� ��v��,�����<G�����?���>��!?84�>0�>���>=8�=fqپd~X��HZ>/!->L�X��N�g|>}�?�;�>�5??b?�<��	����v��=��!?���>��>c�?��>�J�<���jE�2�)�dD��U��(������=e}��͎F>�<�=�a�=��ͽc'.���ѽ)�E�w���E\>�W?�&?5��>���>�;�����H����Q�-��r�=/>=��M>�{6>���=�$�=`��<eB��Y2ý2�|��>����=F|?B#?�A���}��	X�h���q����>Us�>z�>���>�2�=Uo��oS�U�B���=�xE�>ie?���>P<�&�=�d�/ }�7�>QM�>r_>����jG���U��<F��>?��>Ղ��QY�K�o����ۨ>��=IW۽gW�?3�i?�|�(C������P�~��C�v>��->k�w��6�)V�܋8�>X�����ƾ^�l��c�>��?}�1r�>���/l���W��]�ܾ/��G��p?ٛ�>*�k`����������>�ڽ@�_=n Z>J-�>e�	?��@?�S[?�80?%��>	d�a-?{��Ի�=���>U?/?���>���>��?��>Q��������F��g`;D]�|J>.�>�"�>]��:�i���W��ۚ=Ǌ���6�|)��V��+��=��	_��g�}?��"?@���Z�=<[;"��S�}�%=���=�^>o#�ڢ	��=Z��>��?:?÷>�Lr=#뱾A�־V��`N�<^:?��L?���>����>"& ��ٵ�R׼�)>�����2��{	��/߾?`�;&�>��t>���=��>6y?�sL?�`?Ց��G2P��8��J�Ca<ڂӽâ�>�[�>��> ���P[&�2oi���X��z/���ý���m�&�]x�>}��>��>o�>w٨>�@B<�Y�8����X �r��PV>��S>�d�>n	y>�+�����a���9I?�͠�e��W���
˾���w>�S8>���R�?`\���~�_C��z�>�yd�>(�?�?�c?;�A�p����W>�~S>4�>߯M<�E;�����L1>9��=��y�[1��ՓS���T>�4x>�OԽ.Nʾ���M0��,��(�2����<�6�����q"P�`N����r��\I��m�>Gp$�����)��~ݻA�K�r}���HF�e��J�z=���?�%�?�g>.a~��=��o�������M>�8��t���2��, �奄�}��Sc��d�˾�eO��Hi���C�t��>���cp���Չ�݉S�c�A
B>r�?�#��j<�5��	�>y�>�܄>��%�=D������0G��K?<�?�Ҽ�5C���#9<�Nٽ��[>�?��e>Ani��&�����>��?��/?��0=��A����Dq��(=�?t��?�S?�H���=�J�����W�>��?W1?��p���~�o�+?�p-?�)�>m�H�9���FL���>�b?���9_k>o�4?3�?4o&��򾋥�����+�=�"�=�;>Q���1���}�:_��L>ց�>HN��b��2!�>E,��,�0�l>��޹�9�ܾ�W�<�m�>�=���>Ũ7>'T!>��J�W?���5�������C�>���?�Sd?�@�>�.K�R�=�i>A>��/>񈘾I�Թu��>�>�%��:y��"���>�f�?l��?�.�>>o���Gڿ����I�����t�W>_��=�;N>����,T<�y��5�;L�<+�|>{b�> E�>���>0��>���>�c>D؄��S��V��h������i� ����NW|���-�k��
B@�L���C���C<�T$�A���xO��}?'�$<@��.k������%!?���> ?�>��^=�=��5��L���p&>��'%����H���i�˾M������-��,H,�1bD�u���ľG�=?�Q>���$?���=C�x>n�p>9Iǽ��"�⩐=ą�>X>�^>m�Y>_]>>�,=}(���P��j>�j�v
��hP�b=RPm�j�2?������<����Y�����=���>lT<�!־{}��M�A��-�>���;v��b�dAͼ9��>X?F>�o>4����=�e�[> C�=��t>�>y;�6b��Z���sj�>s��>�ɾ͕�=��>p�8?=tp?w!2?�xz=p:�>��!>�s�>9a�=��(>zw>���>�%#?L�D?a	6?�e�>�ks=Vƃ���ʼ��o=b�0��y9�P�꼙'=���<�CL;�KK�C�a=�B�;������=�M�=�|�����:Mq@=Ua�>.'3?��>.�>B���.���K�>���Wt>П��/�?�Ӓ>�9)?ŝ?Ӗ�>>��8>']⽃�����>v>}5j�Hۑ�Q�B=�<m>�<(���>��>j�=�b��\��n*�>Xo?OY ?���>_�?���>�G��9��[�տǶJ�w�+��]�����=m��=��~D��G� �+�}�ƀR�b��=��)>Y�H>G~a>Q`>�*>��>�!�>4�W>�=��Z�_�A�����I�!�a�i<���@E>���=����,��E��j��)
��H"��H�s0��!�?��?�)��݆��rb��a��1���\M�>���>���>d�>��=I]	��EW�OWC��J��+�>ݑg?��>��:� ��=�Q�4;}�>��>~�>ƊE�x�?뗾r~{<q �> ?I{�>��ԳZ��n�:W
�D$�>��=WF�ѡ?�?|?ӏ�{�����5N�3�Ծ��P=X��
��g��N&�&=�7*þv�"��h����"����>w��?�оh;&=q��������%s��^�����_̢��1.?Z�>����ؼ��þ�:�t�������#�=e^c>s��>D�?�*0?+��?Kb�>Ƀ>�l徹�"?,��ΜJ?�E��)�>y4?z!5?dw?N��>z��>�m���O�������ΘZ=b��=��S>�C�>�Q>�=����Ov�<z�;>G~*������9�<���=��>�>?��>�?D)#?v{�������g=��
�~����=?!b>N����� �e=��_>�Q�>�>?.Z?�!O>������R����X=;m?T�:?�@�>k�-��Y>4¾�Ex�B�Q=A�t>�ԼK��������)��C����)�>Z�]>�K�=�[>�<~?��M?(�)?ZBR�4���v�3�C��� >	��t��>b�>dl��g�D�0���n ��qh�c�M�㤹��	8��>���<[`Ҽ�`�><�>>�H�<�Ja=�?�<g�����=@��"�>��?N�,?Eu/>"�	>>�)�N���I?ɔ���6�����R;о���|�>��<>�����?�����}�g���cQ=��w�>Ly�?���?;d?i�C��4���\>WcV>�>k*+<�>>��~�iJ���|3>���=�y�L-�����;o:]>��y>��Ƚ��ʾ�1��+I�ZǱ�l,��ɸ���p�þD�5�5#��� �D�8J=�߾m��t¾�*��R%޽U<�n8���4Ҿ��x����?���?L�|>c7g�_Y2��> �L�� 8���b��"?>����Gk���5���Ƚ�x6ʽ��j�kz#�[��w`?a��� ���#n��=t�?��>.A�>���?�E½7���M	b���?Y��>O{>>T>��^$����e���[��P�?3�#?����۵���>b��=���>#?�Rz>�s��j�ܾ(ą=MD�>��>�U=EU�������X�:�?c��?|�O?��+�شB�/`���4�yH�>��?!�?8cǾ:ξ��)?�?�B�>�4��g��tH�C?jW�?�큾�S�>eL	?k��>o2>�[�&����߾[Ƚ6>�>&>hh�t߷�������Ƚ���>��%>I*�*���$��>{�ܾ�	<���@�w ��b�!I=g?�	�u�=�UG>[!>N)+����+��� ^���0?��?�_?�\ ?=���Ѿܯ��+��=�>�Ǽ>�J�;�즽E��>G�>='�PYo��
��?@;�?���?��9?Hy��o�%~��<tǾ�ں�us�=d��=�.Q>���b�S=�=�2=�� =�f�=D�y>��|>u��>�EL>�5>r�V>k���a �j���4��4�K�Fg&��4�bc^�s �4��V�
�1-����¾3�罙�5��tT���v����o�����=Kp?��R>E�>�o�>͊1>�SI ���6>�;����(�iT�.D�?r
������O��8�ӾN�k��m&����y��>kws>)�=%{�>G�Z���">N �>1�1>|�`>*��>� r>f�_>)��>z\�>�Dw>F_>��:f�=��F>�}g��X��}zD��0�=3�c�?D��C��>�"k��(��o;��h�>��
?��;6x(�1����f��?���=W��� +�0M���(>�>q��>���=$w}��&�5�M��l�>��>0&>�4���͢�����-�`�]Ü>"�v��l
�>�m:?E4m?�Ut?�+ļ��>�{��,�>u��x)6=垝>w+�>��>9�?s�?/1?(��<4՗�ذ�� ��L�8<{0���3>�L�1�&�q��=�$>#5�=�+�=��<��ռ��1����s��%5?��W?6��>y6?��1���X�����q��<0�>�u���2?�?+��>�\�>_��>�V�>/�>P�A�)�7��R�>��f>LeQ�8v���C���=�Ͻ�*?��r?N��=X%ľ��GO�=�������>��F?��?�?�C>o��ɡ��[C����̽[,ٽ���<?S�3��M)½�"˽�½�?켇	x=Y�G>F(=>��A>D��=<�=k�?S�>G;�=�=k>ia%�q��[�Ͻ.�> <���<�D轶�^����=NN�����(Z���.�ký�)��(?��H?Đ�=�!��	t&=���A����=Y��>���>���>^�=���x[�� �?�>8#0?A��?x�?�پ%zS�(�E>#MM>#�>х�>��?�p����� � �Pީ���>>��>`�U>T{�*lG��{2������>�H�=�,����?�5�?��ʾvۥ�1���L����=�C>�ሼ����Ҏ��b���>:��ݭ��U���E���٧?���?9<ܾ��>>�$�~���Ɂ�7� ��{���E�� �2?�0�>?J����={	þ����$�ڽ������^�C|�=Ri��[T�>_�&?��y?^|&?;�0?^D��0�>��z�D*�>S4�=_��>�) ?J�>�l�>�=�>�MJ>�8>#�k��͛��˅=�Y�o�=�7?>h�=ӽ<~2�~�W>┉=H�W=g@�D(���[	>3=?<=17���=p$?H6?�;
=��0=4�=�\�"h��<<�T�>��T]<�{iH�	y�>�T�>�*$?SX?Vn�>�Ƨ�/���o�A�?�9'?@x�>��>O|o>�~�𱯾�㾼s>�U�`�0�>����u���O�%uT>�kI>�F�=Xli>�,h?��S?�m?d�;�|	V�|y�E������<q`>;�y>��7����b�?�r��<l��6�QT����u��<J�v>/�z>w`R>�=1>���='I!�x�=��mӯ�-m���Z�>�>>hM?�m�>H�>hV׾9��p5I?E+��������s���;L���=}.>����s�?Ue��|���ڤD�=�>���?Q7�?��o?K>����ݒs>�OF>���=�:=�#E�o��+�ҽ]�%>k�>� ���ē��6<>�)>#�6>D���������w�Oɵ�ʠM�����[�����G��� ��?�.�����R>��ľ�����ƾ��r];#���4�����7��I?�?i�?�^�=vo�P{,� �����4+ �O��^��=�C��N������b��/߽&���E�/j5�dv����%?��b=`g��U��(o����O�N7>,Ѥ?ӕ����s��AK��2'?��<?Q�>yPȾDȥ�97��N?���?|8�>ta�����p�3>�2�>M�K>��>�R����ھA��Y?��2?C�l>CF5�������w�0�o�Ye�?&U�?��G?�D�S�,��V�Ӌ���>��?��?%i���¾F.�t3+?�,&?Ņ�>�@+��N���!D�ML?m?*��`�>��>K:�>��=`R���.��彾r����>�F�<.���������:��;{��>�*>�Y��!ž!o�>sb�"�G��bD�'x��p5���<W ?f4���>�j>jU>>�)��΋��5���%�ӦE?��?D�P?V'3?����:辽)�����=�Ϻ>땱>m^�=�B��,��>r��>�l��"�v�o��WE?[\�?K��?Q?]�m��9տV���l�оb7���'�=1�=QbR>6ٽ�k=HZ��0Y�;v�;i=Tu�>�P�>͵&>K*>M�U>32>uƉ��L)�����2���E�g2�+����Q�)�u���w��C�þgq��R�%��Ž��ֽ�)�`Ua����v�t����=2i(?���>g>t�$>��`>+�,=D��9�z�2 p����#)��� ��׾痾�M��sK��>�y�� ����90�>���=][�����>Hҍ�xt>�>��>�V0>�D>��>Pn>���>���>�v>��r>���m7�>��?�e|��웿�j��B�;�B���4H?�2 �?P�>���9Q�>z�#���>&b2?)G�_q7��$��ܑ���>��m�|����>�K���O�WB�>�Y�>��[>-�&��1k���>��p>^��>�4>B��=YiA�	�:=cɼ�>=ƹ�9h�=�1�>S=P?��I?��2?�І��.�>c��>���>��^�E!�>�X=`*=-J5?G]?ha2?B�?W��;��j�����}˽$����=#J%=y}���ýV�ظI�5��}�= �>gJy=P���o�4�l���=�\!=6��>59.?�	 ?�?���F�,�O�\�o�b� ��>"���tP?n�>#=?I�`>�LH>q��>��<e�F����L��>0	'>��|��Yf��.%��5�>w�+>��0?��4?7ϣ=!���v*��7^��%�>��&?@�/?���>r�>Xo>f���O�0�e��6A��� ��
��U�p^d�V��VEa����F��|7���;�=��>��C>jK[>r0>¨>U��>�Չ>�}>������r�=>�ܽ=��f<�ϖ>t���N���S���4�qr�y��/y<m���S�Ƿ?�D?�#�S���%�
�������>�>��?��>��>�����8�XC��/c�x?�d?�D�>��c�f���Yo�=�e>z��>~o�>?s>��k��6Q��ʋ��ýE�>y1 ?�e>������B��W���Rѭ>�{�=�A+���?f3k?�B���þ�3����pw�ߌ%���<��i�C���	�5���7���� (��Ӂ�d�
�y#�>�+�?��`�`�=���7��f��闿�g�Awսf���~?��>	"���ʾ����%���E���7����=��>��=�^?�%<?^Vf?�f(?s�W?v�,�3}?#�X�Y�>�o�>��?#�I?Q�>'B�>���>n>t�?�"��톾$�@<Z�s����=��9=���=��><2[=�\��|=G轌�C��m���K=�(>�ah�Rs�=zG>�?"�?�t��Z*�=VX�������2�tF�>��>��4��I���<�'g>��>]?.�?<g�|7ѽ���Q�����@�@�*?10?,�?k�<��|�BXϾ����xi>u��=5?I���J�\�+p����8�>~�>�D>Vpy>L�e?��U?\~?����K\��NW�c���\���<�>�B�>��ӽ�,���j�p�w�2�l�)��p��i�r���n=�6=��
>k	�>�5�>��N>��M=�>�����TI:��O��/>�=U>��?��?B	=7b����B?cP�2�����lџ����<��">�!�=��$�{;#?Z��T��`꘿�$F�!i�>�q�?��?��i?�%ڽ���̜R>d�>�=�~>E���=�Iڽ��=�#>.i���W�o]�T�>��b>�#F����뾲��:qM��whE� ���>b�Ҫ}���μ:＾��ǽ�����<�v�h������H���f�=�¾�ӥ��R���d����?��?Uk&>�����㾰j���?�=�^�zD+�eѾT���OT��%��}wf�8|(�}-8���I�,5����>X3D���{���_���Z�V��+59>��e?�i˾�����|�#�>��a>{r�>{�+n���2��$�E]?��>g�����ڽ[�M=ᇦ>q?>��>l�Խ����a�<��?�z&?���>�*�r���7:��o���5��?��?�+A?�p.�5	;�D�n�K���>?��>u/��ow������D?�D7?�q�>��(K��?����>�	R?��c���Y>�-�>"��>y����ۙ����Z��4�;�9=>��<R�º|���]�οx< ��>b�_>�
;�����6J����+���2�CF��9&��)��v*�=��?g�Ͼ�T>��&>'�Խ��S�@���.]i�v(�=�hy?�}�?`�_?�N�>U$�}����3�+a���Y>wu�>��=���|6�>�r�>c��KƋ����?K��?~�?�P??d.P�Z�Ͽ󪚿�R��R���b�b=8��=J\W>�H��9s�=-�f=�/ѻx_Y�~�=�c�>�Mi>M�>�(�>ӿ�>a�b>F1����#�(����5���L�f��M�
�#]4�d	�k�y��������5 ���.�k��7�<����ňĽW���Ҫ��.��!�?J<o>sy?y�p=oݕ=V�'���ؾt��<�G��O������q�����ze��F&o��S�w���n ܾ!��>� �=�Ɔ>�� ?j���B��т>�Ӗ=ubA>ǈ�>�pk<��	=�!�=�Xs>l*F>Let>�K<>�\�>��^>�0��������נ�kU��z!g?��v=4�����@�4�U��<��b>D�?�^�<�C���y��D~�,��>s����Hq��=x��M��=N�?a�>5��D<I	r���i��)y>S�>�S�=�G=�����$;��f�� �>����<�q�f>��?c��?�&R?�7>�y��>E��=0w�>
����-��P�q=/k�>��?3~Q?�NC?UA?2� =/�B��>='�=�z���2��sr��n���	H���(>:�>�g>��>�ZJ>���=�+��;k����r>�n?=U��>�A?i�g>Ы>iS��X׾�'������>�ڊ�p�u>�T?��>MN5>qU�>\��=̆��5Ͼ#�����>�@�>��q��톿�==CY�> ��>LU?7?�<�K�;�Uk9=l9z=�k >�>I�V?���>��i�\�⽾��4Xӿc�#�!�!��ぽ�	�kQ�;�=���L�|*?:Z�-�`��7�<�Y>�Ӆ>b n>�)E>	">.Z5>!$�>H+J>W�=@�=�U�;�^;EJO�igP=Y0���2<crY�T_���q��b���l6���'Q��K� �x_�?b�?4��b��Cq_�^_��a����>��>t��>m��>���=���KT���>���B�&��>�zh??��>yF9�➶=�
��% <$]�>��>�P>��i�NZ�>T��O'�<�k�>��?�{�>p��6�[��n�$�Fͣ>?�=�[��R+�?�c3?��U���r�m�#�д)�ǩF�Ͱ�>�}Ӽ�>���ξ�(�=�O�\���#�����â=2Z�>y$�?�s��[O=j��A������x����T7��Ï�9�?���>%X�������m ���I��P����>=�Ğ>%[??Uyr? C
?%� ?2?2�m��>R8���:?��>@?�� ?�?i0�>�7�>i�+>!�-�\�+�d�ž&�u=�_�=�����X>��>�Q�R���ɽS�;"�<� <�Jt=C*<���D�>��=�Qj=�J?�x?��ݽ��=7�1�ojĽ�!��J��ޟF>f޽�>�c�P=M�>j��>l�?a�>X���a�T;`3�]a[�*�,?�V?��>Gs����H>�{�v<Ͻ6��>ó=9����j5�����V�>�����1s�<d��>uP>⩂>j8v?�m.??J���%��K���`��<_�ב�>���>�������#>��6��I��D��u��)����2>L����>��<>r�r>G�(>\`>:Y�M>6T���ƽ_έ<�Y�>ɛ�>�'?M3z>�>��Ⱦ?�;*�I?�=��t�������ξ���~>Z<>��Ս?����~}������=�ۣ�>!W�?���?�c?�x@��Z�d�\>ϭS>��>�#_<�=�?C��J��\�4>��=�`z�
"��gm;�Q]>�x>��Ž/ʾ�1�"(@�QmĿ\@��O��]��J.�!ӥ�jE���H���5��[��R���r��p��>������־Aꂾ��þL�s����?�+�?�����{���������C,�#�C>=[�����<��H�<���mq�>��������2��Y����>��>nγ��UU���Z�����7����B>L�C?p7�^:���Y���>E�p>>_�����������	��$?�
 ?����ڽ�)�FV�>F�?�s>媀=&�$�
�z<��j=�% ?��>0�q������w���"ީ?FL�?(?M?�Z���[�T����ľRύ>ߊ?;�?�걾iÀ��u���>�S?9?�C���e�L�iI�>+H?�Cv���>"�?r��>	戽���2ú���,������>�o6=�1_�g�+�۽�5��I>+|�>P����Ӎ���>c8�"�1�e�>����I.%���=�d?�6��p>x�~>�1>@(�9���F��i�F�t�8?�ȯ?RY?+c?@������]�ν�'>-L�>=�>f�=��ܽh>#��>�bþ�XX��f��U�?�@�?���?g�@?�w���ҿ�e����
�N�-�(�N>�˶=�[�>�����I�=�+�>̎U�"dϽe>Mϧ>�p�>1=�>� �>)�&>^FL>�����(�ҡ���[�oO��$=�����������z�(�~�1�~뾵��P:��æ|�8[�=�μ�{���Y<��;��	�Bc?���=9F?}��=tDz>t�9���"�+��Dd�sd����<���ž\L���5E��:`�A������ڠt
?ſ7����=ZT�=K7���<M�>ޞƺ��/>7�>�=���=E�=��M>��>�>#>Jy��ؘ����I=O�`��f~��B�^�ƽ_ )=�LD?N��������]�H���S:a�2�:�+�>�`>8���ʧ�9�2�И	?�/�=��I�t�{��8��>$>bS=?b��Fl��Ml�����=B"����[>�D>��̾cH`�Ά�<��"��>�>�ǵ�H#>��>L�9?��}?>&7?�ּ��>��y>�Ks>��<u:>7��>�>��?�@?#� ?��>W8�=~���z=��=R��:3��T=������9�">=s�@�}��=AJ�=���<8��l�=��-=v�ļ;��;k�?�I2?���>�:�>ˤ���P���B��>�*�>����'��>`��>Ag?��f>�O?6�>TG��ƾ0N�r��>��=�~�E����>c�{>���>�J?��+?V��=gξ
ɀ>J{(>�g)?���>��?B�P>���=i�f=W���O�fCk�n.����I>w~��-��=/�����>4�	?�;���~�!(��Y�>���Z;6?9b1?3h9>y4�>�
�>%�>���=ל$�@=�/��)���	�>d,�=7�� %�.4�O'�S��H�N�TV	>�'�y�ݻ�<�?�w?�fa�ϊJ�H-H�n����;?��>5�>@��>�
�>�)Q>���p{F��|>�ⵊ�A��>� Z?;�>�W˽�g(>�䳽����a6>$>�>P�(>��=���&�����=���>�+?	��>��W�ʉ?���V���޾G�>d��=��E��?L]?����� ��&&��羈@�*�=
o>`��ZM�H�>�	�>�I�^@�,�
��:>���>r�?����%�>�۾r5���O���Pڽ�?#>>Q>Ӏ?�">�J��r�ɾֻ��(m���д�w=}=��?�E�=���>Z�&?�{7?��?d�5?�'?�eǾ��?"��>�)�>4�U>�
?,W?�?�>t?�>m��>�����t�#��	��%��<��>=c|=�w�=���>~������p��=-^��W��|)�=M�=�xW���>�f=�4=�O%>�U?h7?_hh=V=0>&w">��>5�>G
���>�ew��ۑ�˓��TR�8�M?f�?���>vb&>$x�#	K�"�Ͼ��=��?�E?/,�>V�>9��=o6 �,�!�c|,>'�4>�&��}��\�]k�� 5&��ݺ>�5>Fޟ=�G�>ʋ?F�:?��C?aʾ�6B�n/�����d�_=��o��H?�h�>��k��9����ܾ��åC�63���� ;��W��F�[ >5>�"�<O�>��
>�{!�hQ�=b���h2�������>��Z>�O/?ᨍ>�O9>�ڧ��44�6�I?w����e�⠾�eо�����>#�<>: �ѡ?����}�
���<=�N��>(��?���?Z:d?t�C��+��\>bNV>(�>��/<%�>����|���3>��=�~y����=��;]>�*y>��ɽU�ʾV0�x�H������K�Nȃ��ѾW�A��:�xLV����<ٍ�!���댩�����+|a��pϽ� �=�l�K>�U1�8�?���?#�!>�00���+��{Ǿ4*׾�aM>M���G-@�wp��T��<�.콲����LW�����{O���=�5�ؾZ��>!������l،�gGG��>8>��0?9�b�ٻ޾���$l�>���>4�����퉿=Ў�KK��q-W?T8?>�*eվl��=��vE+?{�	?�o>\�־�]I����>�?�\�>�\ǽ�(g��A��jC��J)�?�)�?�VV?�:G��F�f���
D�CC	?� ?H�?s��P���\�F>�q�>��>Ӹ�>��;��៿9�^��p?È? Y��1K�=��?�˶>��&>!���G�4��+,�5W¾�Ŏ>��=0r��{Z������=��>��>}�-��ڒ�0��>2^꾱�N�դH������ ��<"u?X���k>	i>J>�(�T���׉�<���L?���?��S?�]8?�A��"�������=���>���>Sį=X���	�>��>0J�6Lr��p�? ;�?���?�PZ?�m���ο�*�����9���>�=�"7>��>�R��;��Ơ==�뱽��>p@�>��>>cQ>	�>�3�>Ь>M�>I����O'�F���m����$=�H�γ(��AԾ>j1��
����-�q�z������k=�R��IL�<`<��V���i�wG������	?/�:>�c?�{����>a�m�F�־ZＮvξ�@@�MS.�����FվJ���"2�ʎm�4�����Ĥ?j\��|�>�D�>`��=�{�=�{h>I�(>"l=C�l>�I�=�� ��Si(>7J�>�ܥ>`��=H��>�|�>)�{��K���9��x���o��v?���>w⸾d>6�b�`�9�����X>F47?�K>�EF�Δ���c���H�>��%�(�Ծ�,=�h��#z�>�3(?�{�>��q�����tG��aҽ��/=l�4>R��>f�,>�S��K�i�	�+��M�>Ѭ��s�%>�;�>jp?v|?�G?+�h=+��>e�=>��>��X<�D>}._>���>KW?�i5?��?t��>�`s=D�F3=�X=}4��E˼w��v�ӽ��	<��==���>�̋=�ZR�+�=s�	>�X==M���O�=��?�%X?�>�*�>"쵼_J�d8_�[�8��9?�{��
�>_�#?k�?'.>���>�5\>;:޽$Ѿ|��?�|>��p�o^����>#�>>*��>g�?��=?���K�ľ�׆>�,�< ?G�?�)?7��>�*�&����]�ڿg�4��.��U�w`�>C!�R$�����3{�L����[=L�U>�?m��>��(?��3?<�?F	?� �>��o>�u�=��=�Y���/� MཆgC>�fg=y���1��=X��_�f��Y��:{�綐�����v���A�;~$?�?��=MH�n綾-�ׁྴ��>=�;>�F!?܊7?ÎJ>*����B�L�W�	��֍�>_!r?\?�5½I2q>V̻X<�=�1c>v=?������=�V�6�,= ��>�ʑ>�=(�
�/�K���h����ۧ�>�a=�]�7�?�C?G]����־&� ��C�%�>��>E��=p}�6�����
�Y�`�!�x�Ǿ����ۙ=�#�>t��?�]��<X>���}*���k����
���<j�E>{Q)?9o�>���=#�������a��y>Y��>n,�=3��>R�,?�)@?��F?��I?��C?�d�VF�><s\=Un�>��I>�^?#?�U?���>~��>Jdu��h:=?X4�����w�w;@�J�م>�	�>�{;>F����$=�U>K�<��<I�$<�_��ZY<s��=c>3��=��,>�V.?�?4�1���;>�O�~A >�t�>�I�>��=xq���aK�y噾�'����>E 0?��>1}q;��%�6����G��fD?!W?�b�>�Ź�Pr�=��8�+�Ǿa?�=je�>�J���lK�������mS��y^�>�n>���>��z>D�a?1_?��=?l����¾o���-$��+<M]�;�?׬�>���=�22�i�"���l�B�V�^���>����NR�\0�=�h>.~1>d�>-��=��
�z�<��a��T�Y+b�9`�>��>��
?�n�>�z�n���q�:���I?,l���_�Ê��N6оFq��U>�M=>���P?fE���}�����?=����>��?Ŷ�?`�c?}�D�Z��T�\>W>c�>�B-<�>��D��(��}�3>���=,|x�Rc���O�;�3]>�fx>"�ʽ�ʾ��}{F�
7����=������S���w�=�W��>����6�6�ǽ+��������:��վ�=�u�L�g���9�쮴��5��$t�?���?�ը<�W��'I�Pj9��O
�d}8>�W=��X=m$���y0�0+���3��~K���yqj���z�%�"�>#��(���y���;���Fh>p�??肰�Ê��A�["�=�S>��=�����Oz��'��m1]�n�:?�."?y����N޾��ļ�=��?���>S'>i>�,��=[�>#� ?�5G?��=/���H�~�2��=1��?��?�W>?�#*��vC�����sx�}R�>�@?��>�ѾTMQ�Ho(=&��>�ID?K��>�d��{~���#��߹>'Y?xZ��4�=��?淀>��;$ľ�I��I(⾾�ѽ�M'>�8�D�� 霾b|��݀��jf#> ��>ζ]�{ե�fZ�>��Ͼ�g-�3.$�ɧ����K=EY�>��ξ[��<�&!>�W�=F~1��m�������'�� �\?R�?�H?%43?���j/�HOȽ@�:= ��>	��>���=� �_z�>���>��{�M��?�9�?C?�?&�T?��k�v�ۿU���/�a�N8���9�ı�=QTE>ZpH�v�!>/ȉ=mu'�`4#��_�=��=��>0g�>r�>P�(>E6>����%%�U���u����6X���L��x9����a܏��}.���l�Ⱦ�� ����8Ac�<K�>���e�Xo��M�&�r���?U>y
?h�>��>�츾�E�m�n=�m���U(�V3����s�¾Oa+��D*�������3�9�^�о�� ?��a>K|>�-�>e����a>%��>�e�= �>p_>b�H>�=(8"=��=$DH>nL�>7��>&��>�\�>�X��%���t��x�$�۾�Ƃ?�7�>]�-��4�w}�_�����>=�?�X�l/���׆��({���?��
�p�J嘼eǾ�>rg�>�<>��������M�=6��� >�#�>�ٟ>ZI��oT��E���$	>��>,S��է>�6�>��>�zq?��Q?�峾�i�>オ�2>\̊>�O�>p��>���>��S?�?Lt�?�\?u��<�2�;\���x���~��j�=Ѧ̽��>(�9>S�=f����=�p=!W���Q���=J�R>h3w>}k�=��?�"d?�J>u)�>�E����c��8>��
�=��>�t���9{>�R?�m#?���>xJ�=�p�=멿��\ƾ�݂����>�*l>�4S��m���k�>��>�*)=��u?��f?�"
>�w��;�ؖ�;R�>�U?��`?vR�=��}�z&$��X��F޿X���]�'��������=�۩=(���+~�=�=1c־o������t��⃚>tЍ>�-�>i&n>M��;ե�>2f>����>=��>6��<�Hݽ�}X�7Y��U�=��>(`>�|���p߽cN"����#�Ž3y>���?�`??����uA���~�쾜a��$q�>�U�>�{�>Ps�>٘�=����k�N�6�G��gj��Z�>��d?�2�>Od2�r��=�yK��F��l��>�/�>��>>��y��'�~M���� <�
�>�?r��>���3Y�?qh����uڜ>��=(�J�:Ք?�<)?�����K�3��&��d/�G�B>��>%U���⌾]V?�j�]��0.�l ��rx����>���>s�?�Z�W>(��I�w�����录#�=�]E��	?�k�>��̻*��y.� L�)m¾A�d>�?%��=���>�OL?:~N?Lvt?1�?�Y$?cN6��"�>V�ؽ�%�>uz�<<e�>��?>��>�85>�Cn>8)>8��=��:���4��.>WZ����=��0>I4�=?�L���=%Y���F���L�=��ֽ[�üx��=�-����>naX>1R6>v&?k�?s}v�>.��z�C=u)߽J3�>�L�>Ja����]�t����ͽ�=/=��?�|?F��>p5��_�,�	@3����D�;�,&\?��?�P�>lp>`�>[�@�����P=86-=%;����r�6`ѾL7L���>g>[�����>Uـ?I?8?��.?�0Ҿ��}���tѹ��/�C;>RoU?0�?<v�>����D�V5����-���þJ��>�0ʽ�E=��(����>˯�=
3>`��>������/ԾG���!N���>�V?�K�>�N�=;��>�@;�}k5�+j:?�<�����C?^�o����[�=�I>:��;ڲ�Ǐ�>��=e�Gᨿd�8��h�>���?���?Űr?!i��z�!�Z=0�C<Jzp=m#��ƣ�O��=����������>"O:�@Ƚ8��>%��>���>���=�J�#��Z�'=BԷ�o'2���ƾ���*ؒ�}���s׾�}������R=��վ�2������5���d���k�ۇ3��9	����;�?���?,�,��tL��%���A#�F��ǘ�>t�=��@O�sN��j���F�H:��@^�����MPV�'o�3ƾxR�>:�\����\f}�;.�t��"=>�i2?Ež.\����[RQ=��(>!=�侎���7K���
���S?R5?���o��G^ܽ��>�C?؞�>f�'>�t��Bq�����>c\/?��+?U6��+���j���73��<�?\��?��@?5�d��.V���	�w�ȾTg�>�?
?�hݾ�yq��| >H/�>�L3?�?���ıt�[�*����>Q|J?6�I>^?��>�̜�������	�d6̾��<�Q�>B��=N�ǽqg�~Һ������f�>��>�h����x�DR�>M��\��B��Y��ҾB.>�A	?��2��v�>�q>?��=�Gξ)c������汨�'�)?��?�x?���>�_�Gн9�o�x��>ШL>�ݜ>X >��K�Ӌh>e��>?����[�����?)��?���?h?�&u�KӿV��g���2�����=�O�=��>>U�޽�ĭ=�YK=Z���5R>�Æ>#��>��n>�2x>/�T>��<>+�.>����J�#�%Ǥ��֒�=UB�������_g��u	��y����(̴���������ַ����|G�`��w7>��� ���#��=?w	?*��>�A�>�`�>���!w��`^�A�s<r�?��Z�c��A̾�n�y����М���U����pɾ9k�>`�c����>~+?:l�;T��>�>^>HYO>X�+>�:�;=:^�>��>��>_�">c�Ϻ�c�=��U>�Or�=���-��⒌��F����.?`(���@��V�J$�<�L�~75>��?+<�>�#��-{��?���o�#?D]F�:����;E��	��7�>���>�F>���;������*��<���>�c�>�>l=P���&��:��b,��Ǵ>N��?{>\�>��*?*�|?�<?��= ,�>�E>K&�>a�=b�>��>?j�>��>_7?��<?�V�>��<�HT�"_�<}c�<��/�{���IP꽛ZY�t�RE<��=���L>o��=+w�<|��=��Ѽ�~�<'D�=���<HO?"�N?`#>�5�>�����B8�jkv�������>%�0>R�?Q9?���>��>.D�>�.�>£'�kU���p�>愒>��O���`�;�ڽ��>ɪ>S"?;I#?�x�/��'���Ob>%�#?�'�>�?��>�78�<M���2O߿�%�3��ZX>;2�=���<펽�=QO����isk�х�=il>�p2<T�y>�z�>gWX>�w�=��>7/�=�&�=��;�� �pf�ӴW=��>rM�=�4��z
j�tx�����Ĭ=�M�0"�=�62�}���D
_�vi	?h�?�tT�����?�a�����Oz���3�>c�>c�>;��>�=�� �:W�n+>��K7��*�>ae?��>ڐ@�YM�=̀���μ<)�>S`�>�8>I昽_"��Z���<���>�x?�c�>d"���[��%h�4K����>U=z<W�[�s��?��,?��ؾay��}��T�,���
���>敾;���=����>�f4����Ē����.��Qb>���>KĦ?1b�t�S>���dΣ�-������M��>cX�=-J�>���>+�=:Q���S���ɮ�M�7���=��_>�4�=���>��'?��3?��`?rR_?�� ?>��iб>c�<�zf	?f�>_m�>]q?x�)?;z>9�>��>�� �ߌ��I3��~�=Ӈ����=�9=�5>�5�=E�<�i"����=
;|>�M��w#=�>�s佭 V=��>�S?>�i)?Q� ?ҥ��R�=b��=�({<��D>T-D>	�>�������+ܽ��<``?�?#�>QT>*�M���t��R��[?��8? �w>�@`>��=�)ƾ�G��_��_�>����0�VN+�z���]�����=�B&>��!>cAu>'�x?,_6?�2?��Ĕ���u��>�����c#=���>t��>7V<����p�+���S���Z���1���л;3�j=�פ=�u�=?R*>q�=c�=��=��f.����<_Xf��;�>h��>�=
?��H>�=�����k�a�I?�t��3k�@���yJо���%u>Z�<>�����?�?���}������C=����>��?���?3&d?D�&K��k\>�qV>�?>�|0<�a>��F����j3>W��=�jy�	�����;��\>?y>brʽ�ʾP&侰#H�B����w5��)���Y!�?�0�۾�`޾�Ov=§=v���+.(�Â7���a�;9��U�H��;����⩾4־C��?�?���Y���� ������� �=��>�?弼|��>�&=�L����2�
팾�&�h ��m��yT�>2Ӵ��i���[t�ݐh����=��>X^D?$�����ɾz��(Q3>���=��8>C߽{l��F���cT�C;?��?���]{ɾ':=WS��q�>��>��%>E+���tC���?��>��>H�
=�����4����k���?3�?�C?�D�O�E���ܾCF��Օ�>0�?���>:ؾ�;����=E;�>tl?,��>��-�Y����Bf�)�0?�w�?��ľ5�>Y &?v�?8�":?0�#v	=Jä�j�Z�M��>{!w��B�+݆=;����WǾ�c5>���>�	���jk��	�>������2�L�X��m2����	}>���>m��"�>3!>�ɷ>Nuj�˨��%X���}��*?�د?}�i? ,C?�ެ��Э���x= �s=R!?[�?�g꽊'*���8=��>3�׾�{��|Z3��?���?��@G�r?��w���ڿ���z����g��S%#>p|><y>�&���:Q>���=[�����9Q!>�O�>?�h>�~>o�@>��>��l>pr��$�,�t����ȏ�r�(��I0�9)���Y��`ƾ�%����k򆾿����[��0D��>�:����	�`�b�^b���i�P6?���>U�|>8�>��꽶o��)C��w��<��G侃����X���1�=/]�)y���!��g������~>$z7=&�>g~�>=f�>�&�>�O���V5>[��=�A�>���>�`�=�`����w�&�
>�V=�&�>��=z��������4��:K�$�;
�B?	zO�.放�2�$Ӿ�o4�>��?qVG>݀)�u���w�S �>b�<���g��ǽ������>�~�>H��=�������cr�r�󽬠�=��>bh>p��:�q��զ"��=@=���>�:���mo�!�>7?'�{?�iS?(�>?Hu">���>��[>�>lq�>���>�{?�A?��?x�>U= >�Z���<��WT��#���M:ۼ�`�=b�g=~;�=�=r;D���[�=�ff>�I�=2ɑ�a�;>�X�=� ?X0?EF�>ee�>(�b�V���e���>t�=�S�<Y?��>�?�B�>o#�>pȽ����,Bʾ+�I����>O`>�ڊ�"������=�qK=���>3�E?�Y5?�Z���X���>�� >�y�>��>�}
?қe>��=>�
<B���係.z�$V
��&>�����o=҆��n�N�fh˽|����]y��@>l��=lE,>tj�>R�/>��2<ea>���>yT> �
>G�>��"����]p=*D�<C�c">�#��g�����&H��4�P�Ǽ��"�<�h���=J�>X?��A>+������G���9�b�>W�>�1�>h�?sx=�i��a{������4$?��S?�=Y>���5��a�A��5���M>���>t�;>���BA���Ӽhe=<C�>�8-?��>�'T�;�U�@E�H)����>�r�=�y��?Pti?V��w�N�ܫq�4u�� �9���}����C����
�.�ľK���/T��pt�&��>��?�O���$�=^b
��3��T2��V���5=��ӽUB?=Nd=d[�� ����$��z�h5�>��=>��Q>�R�>���>��B?�_�?��K?F� ?$@��M�<?V+�B��>� �>>.D?k�i?ľA?�_R>��3���ҾH�ž���>�3�W�?>oPz=�>G>��=�}L<�e�;Ċk���e>S<==�Ε��G�cZ��BD�N��h�ļ�gW>L[M>>�?6�9?%���v�=�?�>��h=�X0>FT�cm+>�R��*�-���>)��>`�,?�?�,C>����<�l`��l������}@?r�i?��U>��=ja�=���K�-((��?|>�|�
G{��垾�������U�>��>��3� Wu>=Uz?�N?��?<P�ݝ�>�s��� �l�8��Ǽ+��>F-5>D>�Qʾ�6�z|��YV�X�.�����I�'�6=��A>��M>;��=���=�)�=z9�<�cU��=��v��;��н���>��>���>��w>q�ƽs�Ⱦ�K����5?V!��g)ؽ���+q#�P�j��ğ>?�L��z��֎>��!��l��(3���A���>w��?���?��w?*����k�ڻ>~��>�����'"�<cl��`y�
��=���>���u�A`R>>� >;'�>��.�g̴�J{&�����!ÿ��V�e�@�2����R��@��l���X��pv�35>�v��ꇾ ���6����웾�`��?¾ډ�������?y�z?w�>>�|��q�+�J�$�� ���=W������G��s0-=�C���j~�p�پג�<'4�/����5{�=�W��_�u��Rd��!��_�����=��/?�V��G4_�����A�>]
6=;�Z=-<.�����ġٽdQ�?eX?����`�Gf�x�n�%�>y3�>nN�>A�i�!��5��=U?��>8=��zw��;����?T��?��M?�OV;�vS�vr2�{�;�>��>�?�iܽ�o����%�&2?��U?��>��̾�􉿀2A�@Ph>�\9?��O���b>�p=>���=�>�=����mpZ�ڕ��H��=�8>�"���T��♾��8���>o�>ܾ�>��۾�:����>e�ľ��J��pM��?޾P��ň�Pa/?�\ �t�F>�1F>,�>=Eg��承i|�y��=AwB?��?l�K?ǐF?��S���}>��򽸊u>�d?BIQ>+���)�I>AF�>G��T<^����?Z��?�T�?J�x?5mZ��FϿ^��������Z�>�t:=��]>�V��;o=� <����<󮺻b�>	�>@T�>�5w>x�H>p D>�">m)��^�+�Ln��"ґ��C��"��;��`�������j��B������O��W����L���3;��Xн�D9�������4�#?Uy�>���>f��>Pv�J��͕��y�h����;�2վD"ʾ� ԾZ/{�@{��<E�:G���Խ����G�>�޽��>=�?e"��_�#>���>����*}>�1>I�>��>J�U>5t�<o�:rT>�(=>7\�>@(0>`m��Z���.8���#���P<gn)?��\�����0"���ʾ�l��T,�>2g?��>P"2�ԉ�����dӷ>JS���i���ܽ� ܻ4��>��>C"m=%�_��	/�X(��c�.�鯦=74o>j9�==uU=�I�lc:�=c�Y��>�ؾ`V>�Gz>��?�st?}B7?���=���>���>�Ά>�\�=�*>%>�3�>��?
ZB?9�8?��>#`�=w~R�����=<'�Kg����&�����$�w�ٝ�<���9Ƭ�=���=w+���<�=/��o)=mo�;�?��a?��>i#�>|%x��!�_�V����=���=[�I���(?��>� ?ܘ	?���>�]��d��bپx}�����>wπ>�j�6���� >�B�>֒�>aM�>�{?��H���y��$U>��:G?)�C?ü?���>��˽5ƾ��qݿݜU�zf����<�{�=�4>�q+��֎=)�k�>Fq�[$p�1��>rJ?���>�37>%>|N>�ک=�G�>Aȇ>�b�=4e�=$
�<���<��i�L�ҽʧ�<���=R<��H�=��Y�����'�=�m�=���;�0��xڽ�C1?��>h�L��D���H��Ŵ�^.;=� �>��#?�X?�q*?��>�G��d�L��>��ۅ�v��>�H?E�>�-��G\>LH=DMF=��>���='��L8E�"<��7�T��=3�N>�-?�e�>�:��zb`�pV{�/%��_�>k�R=װl��?W?o��	 ��a�3�V@�����b=�����a��.�Ǿ������O��\����$�H>���>�#�?��/��ȼ�����I�z�ß*��>��=��>]�>#4�K㽾�����ʾ���ѿk=�ʆ>��=
��>4�?{�9?,�?�B$?M�/?��Ѿ���>})�<j�>��<�%?�� ?�G?���>�(=C���躾!�?��O��>`�:J��=t�d>z�>>)�s>�UJ��=��=D�c:E|��c� =R��5���\=��>�$�=ڢd>A�>zR?�?��Gt�J��>��=l5>u�8�=���� %�������>{/?�[P?�Y�>�0��`M��n�O����h�I.	?(M?
b�>�3
=��>�"l���|+�;���=^�3�]�Y������š�(w=(��>�Y�>:��=��i>8�|?Sk[?˚5?	�=����S�[�P���j�K�=	��>��=>��ƾ��[�(T���u���(�u�>.�
{4>�¼�ң=L2M>���=$l���ĩ>:���پ��>����>���>�	�>Z6+<���^鑾#X� �;?Wr��D���G��=}���%����>:Z(=Z�����>8%��Z����֠O�Ӧ>J��?=t�?�	p?��=����F<1�慨> �y>�%�hO�<ɤ�=�找�
~�-�N>F��K����R�>ݧU>�b3>��>���þ�����#s��'����G�9�����t��>�׾�ӱ�R#��0��?��I���u �3rt�8���e罸�M��p�W(l��PC�럗?.m�?[`>�J;�R���m�Vr�
�J>{�#��@�=�.M�{��Ug0�*�>���<�s��Ү����_p�d�}>:�P��
��W��^�����u�=*?�K��z������=p�=����	�F�̓�GĽTo]?�j@?1ݾOJ ��}����=���>t��>F�V>���������>ƪ;?#�?˸-�	���ab��q~m�&��?�4�?vl>?���K?������"�?H
?Tg�>銂��ɾ���?�:?Kr�>Y_��7���C#�C��>.�L?hU��f>�L�>�X}>��Ͻ*��gk
�J񢾳 ���hB>Uj�"O;��7^�ޘ'�S�=9�>�>!���zӾ���>���~_��e �(�=��|!��2��F-?����!1?���>hT�=�S����K����[C�}�J?�̰?�i8?�3?����mh���M껨=��ߔ>�K)?U��=�V�v�>�/�>b���q�<���}�
?
F�?h��?%�y?�,L��ҿ ?���ݾ��.�>�|>vR>e[�<{�
>"�a�׏�}M=kX>W��>�k�>�Q�>���=g-�=z�m>�%��C*�"¯�w੿�QH��� ��F�K�����Ҿ��c��S� d������븽�=�p���<��"�����<]x���ޝ=�<=?�Z�>>��>OǨ>�{�<����=�#p#�4�߾��/������[;H|���!�J����i%����
	����u��>z,k=�v=#�)?�A���=WX�>���3xQ>��.>ʘ=��_z�>�r�=G	6>Z�>L?���U�>K�K>�䁿?���Q���߽��6�?�Fk��̢�,��'����/��'�>D�?��5>%e3�3B���숿�>@6�;�>"�������=HJ�>m3�>���=4	�<S�Y�����NJ�+��<TcC>�OX>��=��3���n��|�
7�>��о���=�҃>r�9?��?�-B?��r=�γ>dM5>e܉>�qi=cJ>ުh>��>�?��8?�q&?���>ޚ�=�cU���<��69TzO�w�������<a���=�=��w�= r�=�<�<��=w�k=z���.��kf=CI?�F?�YC>���>��T�L0�=�e��o�w=�D��?L1?�.?^�?���>��q?þ>{��=�����>x4p>�}�������;=6��>�m��?�"? L�=k�����>�>P1?S�N?}�X?���>�����o/��pǿ�F��Ye��S�=�֜=T+>�5e>a�.>�3����ɾw�ٽ�)l>�-�>�w?�ր>�F�<��g�4ڄ>�H�>j�m=p����>��л����h���O�Ū����c��2 }�������9��x���D�=�`�=W֕� �?�(?Ɂ
>�T����d�f��S ߾:U?��;?å ?A�1?��?Q��d��� �2�]=̚�>/�L?�Z�>�'��x>Џ��$W�7��>Q7�>|�A=LX��^���7���<}#�>��G?��>��L��y��U��Q�B����>�=�j9�cƉ?�?g?�w,�S�?�`e7��@�׾[b�=f�%�E(;�־P~8��'5������Ծ93ֻ�
Z>�
?�]�?�i�uE>��C������)7���˽�ɿ>K�>�p?ˌ>+���B�e(����� 2(�!�>s4�>��B>�Z�>Tu&?33?v�?%�a?pF?y���>�:>�����u�>�?q>��1?TLT?&��>�,>���>D=�������p ��vG7>��=;>>A��>\o&>ܽ�3���"������
�b�ƽ�*��v0��z����<�G_=�4>�(?�\R?��o��E�>�j+>��>p���a&�=v������K�=��>R@?�c?$@�> C�=��@�[�������)�(�H\0?��K?��>,�~��n�>r6Ѿ8>n��S=j��=�ϽH�[�V��򼺾\U��Y��>�0�>��j>���>�|?QB0?|�?,xP��y����/���������Q
�>��B>�Op><�����N�F�������.� ����>����M컞��Y�=M:#>m-�=�U�<Cπ=L�����3>�o���>f��>���>�P��ʶ�e@c�u��++?9e���@˽d��=�WA�]�t����>��r�,o�� �.?�Ğ�� |�З���iU�;�v=�y�?���?`e�?o�
6�`ܨ>Iy�>�R<@l�>'�-�󸇽��f��>ؤ�!����_
�,S(��>9X_>��)<�9��#��T�A�@��]��[��:��A�w�
̾����g�彸꘾(�G�`����վ%�v�����i����W``�����˸��^�?c)�?��l>�H����3��?�5����=�XH�ky�=�6��b��Ũ�O:	���[���e)����?���9�>�~Y�3��Wz|���(�B�����<>�'/?Rƾ7y��MI�Nyc=��">�u�<fj�В��	w���A
�GtW?�:?�뾥��|�὿>�V?�i�>�T'>�j��u�潆�>�4?�-?����%��H������s|�?s��?��A?w���>>�f�����Td?��>v��>�&��َվ�[����?c�>?���>���(&����#���>WcP?p�B�P�h>�|�>Ȕ�>4�������;��gw����M�>�)>A�ּ7�|jt�I(���=]��>��o>��|��?���@�>J��r:W��^�X������j"e�;?�<<� �
=3bi<Ũ�6�����xFJ��H�<r�f?g�?92?��M?0���U����K��q{�>�]�>y'W=Q�����>
V	?�Vܾ�0���X�_�f>��? @�6X?1�>���ٿm���0c�gw��q >�>>,�o>v��5�=��ٽ�Z޽=��<�S>R{�>2>^>��R>�+>���=�&1>�(���/�֡��N?����9��澷�辁�����	��m���D�/o����a�����������t�%Y������+y��6>.K/?̚>�]�>t32>��y�ݾ4�Ծh�K����X�iݶ�ǭ��� �
���k���k����᷾��Q�_!�>��=n�>h1?l����=>�>�ѽj�=*_<ݘ�=�5^>�^�>U2�=%�#��3�>�S�=�y>P��=�������/7��U���;�BD?wN\��㚾G"0���Ҿ�U���O�>[
?�L>u)������v�TR�>m�R�>e�#\���'ۼ�>�]�>��=c�ʻ��:��������_�=Yb�>^�>�;�*��6=$���h=X��>�ԾC��=3p>?,6?��?%!??�u=��>�xj>��>�� >�\e>���>MƠ>t2?�c2?S�'?���>b��=:�Q�#0�<-.=�<�p���U4��2~�;��̼˒�<e�c��'6=f��=]~f<66�=o��=H&�#��;u<q�?��I?���>�a�>����;�d9�ڰm=�`>�4`=���>�g$?p�#?�h�>�@O>�k򽘡��޾¾g�_����>�0?>������d�uV�=�R>���>�r+?��?4�M:Wł�	6�>:��=�?N�n?k/>?��>���=�����{��׿�>e��\���=��9=��J����&,���<�ʇ��Z�=ʭ>�H>;�>��[<&l�=()=D�x>�o�>��,>��<�.>��=���W3j�qF>X�X���>�o�=I�j=T��~�.'����La#�f�N=F ���?��%?8�>,:�=a%!�'�!�g�(�J�?�[??�/?��>#� �:�־�j��]�L�j�߽���>r_?�d�>FX��=>��>l��Mo�>�ڶ>ȕ�M&D�R�e��K�+>g?�!?���>�= ��������9���>>b�=��ý���?�a�?18��X�}�D���5�}����A���=��!�x�#��N�
:�r���S�=��A���?�(�?:%þ��>�d�h���D�(��`�VA=|ƽ���? -u=ܷ��Y��8־=v2����aD�>��>�(:>,N�=}�>���>���?!��?u�k?��"��>�i	>�,?^�>;?=TK?2�"?ÿ�=�F>ܦ��>nY�]'e�.��ύO��խ=**>�">+�>(��=\��<�b�=\֦=�к�v|<�3�=N�#>�._>��>��>��?��U?�P�u��=O3�<��k��>���`JD=����5�m����>x��>�N?'q&?�}N>"뙾�+R�>��� ���9?_�-?�B�>�U<rb	<��<����'Aɼ��=�U��xd����꾲9I�c�>��>P�����>���?
�k?'�+?�tN�����.�_ �<_��D�����>Ŋ>�ٯ>�����Ac� �����r�t<o���v��f��|䶼���=,QA>��>�,�<�>��:��z;;m[f=�Uؽ��>8�>��u>H��>�y.>��<K�z���-�@�0?����W̾�������oľ'�>P��>J��?�`	� -��UJ��<���1Ji>9�?��?�a~?���=�㡽/;�>�f�>D�#>�j)=~2>���1>=u-��u�>�u�>�+��������>��u>��=��z=G�����v��=.��󛀿S/����y�˽w{��,�Ǿ}O.>�x��?=`�Y��R��凾s�<���=P����B�O �bn�?���?���=��;�2K���J����Q�>�M��M\�p�|��, ��GҾ����1��R=��lOd���ξ���>��Y�r:����|���(�����W?>�:/?�eƾ�Ҵ�<��O�g=>h%>���<S�>���򭚿~��bW?#�9?bM쾹?����ུ�>��?݁�>�&>-���-��>C54?s�-?
l뼶
���(��~y��vb�?z��?-M?aUܻ��I�ĵ
�/'�?�>]��>�z? h�C�����g<��C?&Q@?�O�>j�n�[H}��7D�� �>�4?��@�>�>1�>ܰ>�M=�m��_)�=�,ž$r	��n�<���-���!՜��m�k�f>���>|�d>{���
����>r߾jZ���+�&S�b��!�t�B<?������?�^�>�=�;��x������ W���B"?ף?	b?�?Ԛ�������8�=~�>b?�� ��lF���>���>T]��Lj2��x���"?�_�?4�?~�i?�yQ��ӿJR���۸����j�=i�=T�;>r��>��=�b5=ϳ��H��d>�x�>�'r>Rx>ݷS>�>:>@�)>�>��7�#�����Qؒ��@�����+�ʍj�9�	�/�x�nK��k��罾j]��Y+��*���QE��-��v>�n����D3>U�??9
�>�[
?��>џ>>�ɾ�[���c���K�a� �Y��k�� ��6'�<��>�'��fv	�狾z+��D�>����|�#>).?QH��6��>j|�>�0����>ڽZ>���>Ts�>�Q>���=�r�=�>���<�>g��=�ㄿ޾���7���M��F<��A?d�`�M��ߞ1��H۾W�����>�
?:�O>�J)�@��O)x��=�>��I���b���½E���>���>)��='�ɻ��g�|����+�=�[�>�(	>�<ӻ����r���v=��>Cվz�=��v>R.*?��w?��5?�ɓ=mx�>%�X>	��>r��=	�K>�Q>���>��?T>:?�T0?r��>v{�=\Wn���=G9=�/H�\�;�Ő����ż��G
v<u?%�/�v=o|=��<�+}=��>=�ڰ��S[<�{�<gB?H�:?B7�>z��>0&`�o�-�5-�oA��>�M>[c<����>g�>�?�f�>W��>�OX=�X@�CD������[��>R�B>����v�����='�>MӔ>9O?�7"?�7R�h�t=�n>`�=B��>�
8?W#?%�O>���=8I��{[���Կ�h�S�^�)��>Wq�>h歽K<ϾCþ�Գ�����$�?��>h;?��>4K�>�*Y>p���ч��a�>�Qe<��0=+	�=��w���C�X�ٽ1>��M+$>p� =�t>e ���@��X��ˣ���I�<X"=��7>��?�)?u,�=K�=�ԭ��Ir��m��(?�n?āO?fcQ?Ϫ"<�)��� ?���ഏ�Q>hmL?��>Hr=��.>&����]w��@�>�ρ>N�=!Vڽ���b��������>B�?vV=
&dC�	T���;����>�Z�=?��֢?�lr?*��@/���<��65���x�5Ԭ=�k.�{����ʚ�m�	����7Ҩ��<��gP��� #?V۝?O����|>j������� W�Vi�>�a�>�A%?r�D���d��1��%����u��͔����>n�>�6�=2ػ>��?&$?"�p?�r??�%?�]w���>���<ϭ�>��>x� ?�� ?�` ?{ h>^�`>ݽf�f��C�1y��y�qwR�t�=%>V��=����0=0��<�	=�=��=���=-8.=�Qr=Ȫ=9 D>��.>=?�K?[bȽT�>鷼>0�i>��>&.�/u��0�ݾ<G���n�3�>,68?9�;?��>@Jf��>g��낿+t!���BD6?A�3?��>.;�=��=� ��
�������N+ѽQ����<��h-�6�¾	�2�A�>��W>m	��P�>���?�M?G$&?�T%��p���#���Ri&���Q�8 �>��U=�T>5J¾�k�+��޴x��d,�uF]>�2��#<1���j� �d>��:>��>r�%���9�g�I��'2�G��<�
�>0�?�9�>*������-����W��H6?v���;����ཏ��X@����>D�]�������>��ؾKE��Y����,q�f&�>ڋ�?Y��?�Hz?�R��o�o#�>Wa?B)�>��I>���C"F�>-˾���=��A� 
�b����蔽�p�>>z>>Xm;}Eʾ����d���s��v[�!�6�5&ྞ���[������5�=�v���ݠ�Hd��H��=�设܂#=�Ʀ����em��%�[��f�n��?z�?��=>k�ͽ�Z�ַC��<��>��O��>>�`��܍����+�{H���21�CoھH�����V�x��>��G��	���'p�Ok7��p�
�=��H?~d���������}�=�؝=��뼴n�@j��j+��y�ӽlNi?SJ?�sᾪ��t⸼q�2=T/?Z�>�*>{?���Ž�a�>ގ?��,?�2�������ɉ� ��S�?[�?=�F?���;�A�C��<��+��>�(?��>�楾�e��u=��?T�A?���><����E3S�J�U>��@?@�_���A>�+}>?]R>�� =;L�:��̃��Y�� η=&S��n�u/��� �b�}>D?@jW>>�̾o�"�t<�>1�`����u�Z�)��?�<��+<�	v?�Y�9�>�`>��c���e엿 ��q��tO?�=�?M�D?��2?k��u��^�s>5��>��=��>s�J>��W�Z�>X��>���I�m�8�2�-c�>V�@=�@��K?k���i�ܿAX��F&��yԾ�P�=���;���>%�2<���=�6~=��ĽP�̽|��=.5�>�j�>��+>�'>�1>�9> ̇��/"�kN���͎��V��e_����a�x�%���`��V󾨬�T�񾱢2�����o��o��%&:�sc��ߞ�,���!?���>"2>�c>�B(>�����r߾�1�^z�.
�����ӓ�]���F2����[����[d���,?��>);�=_u�>�w!��5�=���>a3=�:>^�:>@�P>դ�>s�\>�s�=Dk%>��>Pw)��~{>s��=ٗ���倿�[9��Q���7:�XB?N�Z�����LG3��M޾hA�� �>�?fR>��'�A���aLy�&q�>Y�I�'}c�y�Ƚ���\ԉ>���>���=	4ɻ���!y�4h��Ա=r	�>ǒ>U]�(������*�=�?����JϽ<J�=B?��??�t? �>�?˻V�;U�=��>ڥM=y�>�P?�Q4?I�X?��?�߯>��=Wj��B��<wE_�bb���̽ٹ=���;@�<�K=��ｒJ���=
�h=�}>��M=(1o�􊒽�M&=��?�tl?Ӡ�>+��>?��@�5����w~>�����)?�?�2;?�_?�?*�>D�2�1�����Lh�>	�>'��q��/Ѽ�S�>Z�����,?cX ?�(�Y���g#<}�>/r ?�s7?,�?龓>�<�'�����ɿ�J�~?��v��ˤ�}��������'�D�˽2��O[�qF���>�"M>KT�<
;91��=y�1>�R�>�:6>8�<�m�<��w=@�X=��Y��U�=C�<"�۽��	�&=F�<�7���Gg�cC��40�����U��h ?�x�>�iI��T��J��[Jﾄ�|�&ע>��>�&?��>v��<��	��Xh���D�������>ƅe?���>��J�R;�1�=�6'=���>���>�M�=
j���G�Ӛо�N>�>P�&?��>"$�ƀa���z��%�rf�>!n��������?�X?h ��>;�.t;o�����oL�=J�v�ǃȾK���&�"�g,j�� �����_|��B>l`�>(��?Q~�ܱ��#�S�}�/��1�:�5��=�r=���>�b=��mU��@�=��#����_����4��p-?ז�>�{z>J&%?�ZC?`�?��U?�>�=��>ė��ܙR>�e;?�?%�5? 7 ?��>�[>�x?�H͎���Ƚop�S���L�V�E>qێ>b�p>��\�o��=e`�=��N��H�����!�!�ӽ������=�+�>J(�=�?^X?ϡ�=�mD>��z>9��GX��Xb�=iX�>�о"]��`�> ��>?�C?�fe?rf�>���&�,�g�=��+˾y�;�� ?��d?�?Ҁ=| i>�2�)����BǼ�j�=-q>�+��+��������K�͛r>Rs�>��->�->���?�
?��>�$7������q�d�D�%��>�S�>�?�n>��w�B:��*�C_o���T�5#�-��>�O}�>��L�m<�Wx>O�>��Ἄ�;>�N)=��:�d�S�g�=	X>9�3>/�>�>-?���>D�<��Ǿ'�^?RT��Y�R�t⽾�P��Ӗ�5�>��>ȥ���c?J�$��?Z�u_���:���f���?���?�$�?������e��$M>�>?�v�<K�=��=���
�G� ����>c=�m㾎c��	��&�=rB>$���E
!�T�<==��ؿ
Jc�j�$�܅羛����*A�M:�����hп�,� �H�����*�rd3�'g˽�";�
׾�Ğ��X��X�?F�W?���e���E���� l�)?�:����7Խ��8R�B���x����վ����$�ږ�Y���b*[=@���ɑ��+��*��q+����>�(?�v�_]�}�Ӿ��}�4��=���<�����Sՙ�\����m?ЍW?�ȟ��E�3�����@T?鱠>R��>Rd׾��>�	>�1�>��u?��k�����2�s�Ez=Ԧ�?��?��??��O���A������4?5�?���>�����̾�N�I?��9?�̼>��^��s(���>�[?C>N�ځb>h��>F%�>�𽇲���'&��3��h$���9>�g�I���2h��>��	�=��>�rx>-]�&���~_�>z��V-���I�}��l�E>�H�<JF!?��?���>N7p��,�������Z v��0��s�J?�~�?kf?�'?Ik ��z���R>%۽�[�=X9�>�� >al����>��>���Y��Qt?���?�5�?{P@��U?������Ͽg�o���V���ź=���=�J>�Ϲ�i��=L�e=TzY=F���8�=^>�>��>��}>��Q>�S>3>|���T*����P���eG�������i�l�Z�2�w����
t��m�ž
*u�����`��=�l��K�&	ҼK���H�z%?�!>$�>I�>��>IG���-�������G�־�������� J��TO%�'����&�!��o)?�?>h5>|ұ>1���L>>hM>&�W=�\2>�:L�@�N>מ>ğg>E�>�:=�n�<5���Vo>$��=6��QM����9�c]]�,s6;�@?��_�8ڗ�2�������)T�>�a	?�eL>"+)��o��8Hx����>�AE�ae��˽��v�>g+�>���=��� ���r���ｬڷ=��{>�>{\�/]��������=n?���X=xr��??�O�?�DW?A�>��?�1�=�y/>�>�B>��y>��>_2*?�yF?g?/W�>S=e��H����'��'���⠽o䞽��<?d�<*�>4T=r挻���� %�?�)��#�����;�<|0�*�?�5h?B��>[��>�t��$�C�a���X&����	>-�/�L?���>%N"?��+?he?�K�=����]��f.��ɢ>R!>�'U��.j�8R�=L:>�h�=c-?@�<?�P�o2��?��=��=.?��4?��(?�E>�q�=2�y��A��Nȿ���5�"�*U	��XO�X�<�Nq��Y޽y>�<	R�K�]��	���g>u۔>�>���<��=�x�=*��>��M>_̋=��=���1�<����H$�=l�����=�v������ /<��ν3)�' �����������=�?O��>���e(Y�ξV�����7�=9a�>7�?n�y>D�N>���\�o��Ra�>_?���?.�r?��>,�;�h3��Q�>%�G���?up�>*��=z�꺈2R��S���F=���>.�$?��>��� <X�3���/�1�>�M<����A��?�?c?���]5D��X���l��y��~�>�7��𞷾v����+�/�l������᾵�r��<)>D"�>�k�?�1��=%$�GЎ�^Y��{������=,H�>���>L��=��+�t�=`���0
�M����OQ��%?Ӌ�>k-�>��?�1?_Ў?��*?n�>��	>��+?<����d�>�/L?D?�uK?��I?�D=?���>t6�����MX\��)��Fr+>���<�?>��L>Yw=>f�׽8��AO�=��1�@����<L�<�@:�իl=i�C>Lz�=���=�?|B?|�W��=3��=��ܽ�A�=�>�>,㒾z��Ji�=lH�>(?t�O?-�?f�������%�_����~�?׃F?\��>'�=L�]>x���O���l�=k>�� >�0�g׾�Z��
`o=�=�>�ߒ>�}> >v�z?�h?ח?<���pq6��]h��mԾy��>�9> ?3�A>&��3 ������a��9?����LF�>������sJf�I@,>9O�>َ|=tS�>�(>v���笖��C�<Z��=>?��?Y;�=mJ�=릡�{ �N�:?!i��._3�S㔾F?��+�>:�>k�5<�#�[�.?�Q��o�J�Ʈ����^�R��>q��?A��?
��?-�M�RJi���>گ�>�E�񠞽�ľ�e=b�Ѿ���>.��=CƐ��N=:d��f��=���)��ؾ�`�����忙Gx��fo���Ҿ�����C�����f �����7#I�Sb۾V����;A����|��Ȟ�7� ������Z�?��\?���&H��_�JQ'� ����
S=�޾�>z�ؽ������*��F�lP�{��-4���	�A�ʾ���=���s(���9��6�����<��:=�5?W�7�>�qO�&
־0��>p1	����a������7pƺ�<w?�Y?l+���O����끵=�l?�>_k�=Ħ�k��=��G=�S�>	�Q?�B������ſ��*��=�y�?���?h�??�P���A�#�W��F?з?���>����f�̾w�z?	�9?���>��W�����+�>��[?�FN���a>k��>�2�>y��ˎ���p&�g��ń�e�9>H�	����-@h�W;>�2<�=	'�>��x>K ]�����)C�F2��6��Йg�i�E��Y�gIž�*O?e�m�tm?|IP>�ƾ����㖿����������?��?2�U?�,2?!0�a]���>��>X��>�j>J�[��� ?`��>����J��Ӿ�L�>D��?��?@oZ?#����A��ݎ��wR��3����=�:=Q.:>(�!�I��=V/A�_=ᜈ<�>�މ>&�_>��:>�#>>�8>����I$��[��ߖ��yfS�]�?�����>
���+�t*��������3о'ɠ��!���Ҭ��#ľ��Q�7x�<e��s�*B<?��I>�N�>�v	=N��>	^�Ꜿ�����x3����l?"�R �� �_������}R�Ӂݾ�U�����?s�:�ѐ�>=��>�T����>/�>������E=�#p>��>Q��>���>��>��G��ڼ<���g�{>�c�=���=����$:���P���; �C?�\�����̕3��1߾R������>��?8�S>,k'�@����x����>��E�,Hc��̽O �Ϛ�>:��>���=��Ż�M��qw�~�8��=\G�>��
>��b�(���������=�H>?�Y��vA4>A���?t��?N)>?f̭>S�&?�u�=.w>�v>c>���>_�>V� ?��@?�$-?�>A��>�B�ƭ���9<�E��>zj��9�{�< ��=��&>��:���½,�0)=e=H=�I�M��� �=��>��Y?���>>W�>t�=���ApL�|*�\�j>y?��]�?�m1?��F?�I?<�<?�-�>K�ֽ��!��$�'O�>�Lv>�3;���3�X�>���=f���,�>r��>����q�
��>��#>���>[�?���>T��>G���#J�W��Pxӿw�#�~�!���������7�;�@=�[@L�����n.��������<�!\>���>{Up>�uD>b�>��2>�7�>d�F>�#�=���=�O�;�=;h�G���N=T����D<�WU��ү�U?��b㖽Ὴ��KJ�C�@����ټg��>���>c�B�r沽96���i��f"���>���>�U?l9T>x�$=���^d��?F�"���>�>u?��>O>C��>Ͱ2>-SQ��p�>ÿ�>B�>5'j���-�"��������?61�>P��>+�1��HF�$�|�q=�{��>x���xF�U�{?.;�?3@�|���?��d]����aT>>!���U���m���q%���F�#ξ�u!��F����>���>ܑ�?�J�{��>�8�Lߚ�V-�������E�,W,>�_?ćC>��Ѽ����<_3�.�־<�：^2��%?�>�7�>�C�>�Z�>�tp?�r;?�u�>iaA>��.?i$�*��>��?��>0,?+2?O�	?���>uzu�ZC@��������E�<> $�d�۽,�=<CX>z�>
��< 9�=>���k���;F���3��ܽW�>���	>��>ן�=��?ET;?�N��g=*7o>�<\��uz=E}>;�l�h��=��>cw>�!?IaD?�y ?)߻=��"�����HҾ�&�� �>a(?|��>���<p��=Wᓾ�G��N�=[Lh>}]������Sd�R�Ͼ��A�=�8>���>�3>ݷ�=�*�?��>BP8?𩊾[`C��B��[?�r�'�J  >�#�>ү}=<O�����N�S�����ݖb�
�5�5x�>��:���K<J/>M=�U?-�/>�<)=Qt�<9�(���y��	�Tnf=v:>�l�>�Z?��=��<�+��.�;�?
�쾒�1�Xt�'�,��j��-|I>j�O> �6� U_?�=��7�����]�T���(>
h�?�U�?�֎?z���T��aW�>5N?��i>v�-=��O4>5)�:M?�8=�-�m%d=�+(��EV>��>X׽��7����S�#=<t����|��Hi�����s��D�޾�-����������y�j]�N��M=�����J��.���z��e���U�����-?�|<?�|!���<_Q������Ӿ� >L�����V����Ѿ�_��`�"ľ΍"�~�;�sl�����HP~�Ծߙ��t���F�uܴ�8��=�,1?���$���������\�Ì.>"먾qH �T���t]���Ū��Xv?��$?�釾{����W���;c?��[>af�=��N�9�>��O>b�?�=k?��h�����Q��H>��?T�?��??��O�Y�A�����;-?��?��>���P�̾�(�!?��9?JӼ>/��_��s)��>��[?C)N��xb>I��>�7�>���o����(&�;��߅�N�9>�������`h��!>����=��>iRx>L]����>���䓿v�\�p94�pڼGs�'�"?�C����>z��>[����㾘ї�𩋿��E��`'?b��?H6e?�M(?�������Ë>Rn���=�w�>ݑ�>K���x�/>��7?�wW����"!	�t?�m�?���?m�_?e�{�T�ܿ+������"����^=
`�<!�*>����:�=ٔ=��L�_9�0�=,��>qSO>m�>s�9>uC>��2>�`���K-�hN���-��7O�?�	��SR=�����R��&��G羕h��J�ýM�潠I��Jz�x?h��ȼ\L����T�d��>��,>D�q>�.�=T�H>�@F�A���v��_=�kʾ�9%��5
�����;�8��M	��~��d�F�D���
?(\�=畍>��>��[�H�X>U��>��'<�y<��+>>�>r��>��?��%>Hc#>���>�>ҟ^>��=喂�����88�-�d��c"��??��@�{K���4�f來7��+0{>�?TxD>��)�C"����u���>�Q?�q�e�=Zý�ļ{�>��>J�=�*S�����>z�:ݽ�&�=vj|>��>�ܼ�Q��fw���=��
? �%����T���.2?���?'�_?��>?���9׭�s��>�%J�w�>'�?fL?EdD?w�?���>	J�<�`սA=>�c����S�-ٝ�.�G�i���OdǼWV>��u=u�=��A>���=@Q�=���"4�=�	v=�=�	?(�g?i�?n
�>�M���#P�ѽa��9��V��=;�J��>��>[�%?�l<?�-?��<���dz��5?��ҧ>*��=�S]�Qj]�-s=>��>{��>X&f?�C?��K������7�>��>,?��*?��>�&>�9��JB�#~ؿ���ߧ'���ʽjJa��R	�0��S2r��M��m�K#�.w`<^J>Q�l>�cc> �O>+f>�x0>X�>�u>�M�=���=1��<i�(;׸,����,�Z��<�_����Y����tXŽB�~���x�Ir���*�Ҡ�3K�>q�>먠�{�Q�S�	�~o)�V���.?0A��U<?��>?9�=�,J�����\3���{q�@#6?a^?���>������H��C�>�޽��	�>�{�>��u>AF��\�����j��;2?W v>� >�F��Y��Kp���=����=aY1=�p�=l&�?��Y?��'��B���L*�\PC�����>����ྣtm���
��r ���.�9��R[��Rm_>П?ߪ�?��+�<�>c
�����������?K;>�e�>2?([�=c'���\�V� �����;e&"��l?�ް>��E>'9�>�{M?���?n�9?*�;?O��j�>���Y"B>W�$?<uC?�S1?7	?Dv?�g>��eҷ���ν;n���K�E�$���=�mY><��>��K>>�Lv;�#4�K��ɵ�w ��c���D�=A�t=}�X>�a�>�F?�|??��A��
[>�׳=�(���k��V6<�/>�O��%����=3�>�:?��d?�q�>�.����,]]�0�Ӿ� N�Ac�>��4?k}?��2>�I�>o"��6��)r�=o��>ԭ�=�p콦uþ�㾀9�=��>X�t>$*I>�`>IN�?~u?OH>?�����2����[UN�Z�M��� ���>��|>:r��7S����)y��򅿺�O����=H］���<챁=�n>/��>�L����9=w���y��_ꤾ�VR���2>B�{><b?Rj�>�~8>oY������Z5��)?꽣���D��:��w����&���2>��?*ݾW7?��P>��j��椿SY�e�2>��?I��?�_�?E$��##��o=>���>��>���$�ʾ�8>`c����>�Dw>�'���=߼4�=n��>f�>'�w��[��/�i:�=D�ѿ�5�y+�<E�9�䓝��� �x�ܾn���<�>G5꽼Y��VҾd�p=�݂�D���7荾�-�������uU�\mv?���?+��=-.�	\������T�'�������^�4&Ѿ	s��<U��?f�G��� ���7���~�����2=���љ�+���$��3{h�3��.��>4�v�[�5��kX�� ��5�4>�c��\�6�Ux���혿�]ǽ::P?knV?>Ų�ByN����ٝ�rt>?��>�er>�QҾ� �>��>-�w>��C?�j�)�c���l��V�<���?L+�?o�??
XP�͕A�v��T��fr?|�?߇�>?"���̾%��t?5�9?�F�>/C�i�������>{L[?�MN��Qb>k��>Hg�>+��5���\&�����Ut�.�8>�7����)�g���>�C\�=!��>�[w>��\����.�>�����X�/@��!�¾�X�>y����>��>+��Z�'��V%�-���$��i�w���a?���?Hu(?!H?L����V���;�
(>'`�>��u>��?��ȾjU�>�c�>l|����C�qCk��8?>6�?ȿ@�Ij?=�k���ѿ�H���Ӿ����{>3�F>=|>��	��#�:Aj��e�j ��b>%�>��y>��(>4�O>���=R�!�A���Dz'��7��"R����&�������Hؽ3���4���D�վ9d��!���'���7�OSl�>"���?��M��+=� ?��>v�#>�3:��I>c����߾�{������7���f?���8��\�~ro�y����S���2���?l@< >�>�s��4x�<�\�>�����LD>��>��?G�d>F�	>�qN>�N�<�2�=V,=�}y>��=i儿�-���:�ZzQ�W
�;��B?�k[�==���	4��w߾�ʩ�;��>�?LR>�z'��R��(cx���>:�B�(�b��=Ͻ"��rˈ>5~�>�8�=e7��Z��9�w����g�=�>��	>Y�o��F��7���=��?���P�n=�:�>�/Y?^��?z�K?�LX>8�?{c��b�J>	z�>�	�>�<�>=�?~R?��/?j�'?���>��=V ��� w���$=���hH_�l��8X�=�RF=��=R��=���=�a`>fV>�R�=�v�=�"�=�J	>2���h;?��c?�?��>@�Z���9�	^�K���հ˼'����?B�>�w:?��3?�@?�d!= .�,I�I�Q�>}��=.:��J{��, >b�?Y�w>O�U?�
?����H��)x�I�,=Yj�>�$*?ٞ?�ؽ>`�����|��
���	��n,+�1�h�G>�*_>�v��1�M�<�;X�R�_Z��M%���IR>UI>tA�<$��<U���/t����>|3>p >�N��|/c=:���5�(�ƽ��>�U�=��¼i��gF��ԖV���O�+A�;�% �E�\>Ï>�?�f?�K���>�A�Ծ���B.��|�>�6O>��!?h��>ܺ:<k5�.f���6�}�0�`��>�UA?��>=i�����a�S>iؼ5� ?B��>�EI=�zٽ�������\p=��>��?��>�mZ�}�]��;��ؚ
�A��=S�=QG�c%�?�mj?��վ�؞��
�K�B����u,$=u#V��c�9+?��_$���a�C��Y	�����]N=)��>��?�����W>�����i��p��zʾ̣�>�͚=~��>)��<�z����M���V��o	��#����=-5�>�	(>�T.>j5?��?��m?��B?R�?H����?8�@��>e_ ?��?�V?�\?Å�>A>�C����8��A���3���-={�t=�9 A'>{�=y�Q=i�9�{�����<�5�<V�>���=2U=K5t=-�-=��=��N>a0?i�.?���=��;&B'�mz���iD���=<F�=��P����=2̸>;�?�.O?��>�R ����U �͈����<!h?�6?N�?p�=א=`��w��Ŗ<l�J=d�`�%�N������.��� �D>Dڙ>�3z=c�>1̍?`? \1?B3����]E.����+�>��=c�K?s9?5Q�>���\>�p�e���Y�����Z�>Boܼ���=��>��<���;X�7�Q=a�fh���4�� _>��> �c>~��>Hz�>�ʾ=xi<���9G��]S?���v�"^���H��($��?DC?�
��OP?��N������a���?�:�?��?#c�?TFB>c�����=@��>��>�Z��g�ھ$�>d�� �9=�>Z3��x��m����>�=�M�������6�+>Ų�4�K�x�-��F�`*�Iȗ���쾃_�p ����.�
"��Kt|��4���U��nr�l<o�CЙ��@d������5�?%b?�*/>W��� -4��$�Ω��3��=�D����=!��𖗾i�_���E�˾[�쾧q	��S��?�@�ؗ�>X�[��)������=�'��7�3�(>	4)?�*��K����E�Z0=� >�$�<@�������J�����wU?"�8?�߾�����n���=4?��>��&>�ޒ�Q#Ž��>�D,?�Z+?b����B���	L�:���?b��?#�??
�O��A�i�����'?�?��>溊�	�̾&�?��9?�>���a��b8����>�[?vGN�sxb>���>eA�>��d����y&��-��u!��x�9>���7���h��>�@w�=��>�_x>�]�B������>ӹ��,O�P�H�����# ��P^<��?K}�ϰ>��g>��>��(�9@��3�����վL?�o�?j%R?��8?�:������c͊=$��>�w�>�=Lu
��$�>[V�>d��Z4r�θ�ؙ?�b�?p�?ҐY?��m�Gӿ��ܶ�����+��=k'�=/�>>��޽�ɭ=��K=Nט��V=���>9��>�o>�:x>�T>7�<>��.>`���}�#��ʤ�4ْ�\B�� ���wg�|	�Ly�����ȴ��񽾮��������Г��G�x��:S>��̅�Ry>h0�>��>�l>���=_�D>R����$ �ꒇ������A$�%���Q���*������t���$d��͋����lR���C?��:�?�>�?��1>���;�n�>��
>���>��>���=�]�=F�>��>s�>V>煌>���>���=�������'���켾�=���m�?��o�m�+��9�*��
K����>hl??R>�Sd�����/���J�
?��s�`�A����=*UA��\B><�?B��;�<�g���:�������%>��)?�� >�y�<���O�޾+º=#?ض#��A>��;>8/D?���?Xe5?�K��;G>��?�Ӯ=���=���>#�=��>�8_=lNk?�V?)OB?��m<N����ؚ��!��Ք���E������F�;0�,��H=l����_׽?�>��?=~�>�	׽�@�=7�=;�D=�$�>i%l?�?��?������/�x4;��<��F�b��t�;j?P�?R�?���>.��>:�>�t<v�G���T�9��>��8>v�N�ZRD������=�!�>�mP?�RA?�ĽǙ���?�=����12�=��)?"�8?�J�>�c->���=�~�Լ�1&�';���ٽ��j��ܰ�ua����X=/�v�Ft��&�'Gӽ@���F+=�ޭ>�n> �W>�=N>�u�>z�:>���ͭ=�h}�^�s������ >���Ѽt>[(�>kf�=N�=<����#ֻ�P�<�8>{���<	?�K?���=a��<� ��n澕ָ���>�Y�>���>n�>��g>��j�J�^�6��R����>�[?a:�>�a����<��ּ,�<��>+!�>�	�>����VB�12��:���]�>q?q*�>l�A�O-r�3PX�n��	��>���<��6�Q��?@��?r��?S���ھ~�I���w�">���>N���
��}����*��	�u��0�`Ѹ=M�>�]�?J�=6q�>��O�x�j���|�m+��=�w��W�@��>+�ۻ�Z#=��������lp�8tp���=��<>��=���>�5.?�X?Sl?��?k?]'z����>��>>�P�>�*�>ݬ�>� ?`��>"��>��P><Y[<l��<��5���ʾ��<t���� >g+�>DG>���=�.���i>�b=SB��ν=��>��=vNļ�z >.�=�|w>߯?�X%?�����$༩� <�����>�n >_>]l�n�þ�5��?�=��!?�"?���>mD�������ƾ�,#���S���2?�A?���>H�|> J���{D���Z�>e��>�gx>R���C�2��*��UI�>i�>7)�=��W>FX�?�.b?�<?&��I&�Jς�^�?�T�m�?x��1�>�[�>Mg>����ńK�i�4�5ae���2���^��}T����=�a&>�l�<��F>D���ӄ���=�4e��z4����Vf�>ܶ�>��>U��>XĤ>���=s.���s����I?����l�r�Ekо�J�!�>��<>�����?:�O�}�_���B=�I��>��?���?�Bd?��C��-�\>�/V>��>r�.<ϣ>�(������3>��=�qy�����;<�\>�Ly>��ɽ��ʾ2�@�H�q�ȿ0�L�q�ƾL%��ƙ����U�>9ϵ=�Ǿr��'N�]$��@�Iؓ��鼽޽ͽ.=��p��?9,r?��<�*W���+��ټ���ᾲ��>����+���;�\�ZB~��`ܾX�����پ;��� ���:�u<�>M�X�����.{��)+��}˼�>>�H/?�:ȾK�����ݖ-=R�$>�V	=p�Q.���Ϛ����އS?W5?������BɽB�>c�
?0��>�>�C��)�ν�I�>��3?i,?���+���ԋ�}�����?x�?��:?�?ɾ�(������ż>(?�Y?�,�>[�n��'	��W��!�
?t:j?�Ŭ>C������Z�B(%?�B�?>n��9d>s�>��>���<iON�r._�VUI>�2q=8��=��Z�5fھ�T�i�=�=�>���=�G���Ͼ}�>���m�P���J�n���O&��!;�?�����=��^>@C>�'��č�W��2���kL?�T�?�N?��9?�4������%��9�]=Xç>^ӧ>�=6�����>�|�>$��r/q�?��)?���?[A�?�U?1�p��	׿�覿(����ؾW��=�n�=J�>���h�<���=�8>��=%�8=��>��>[�>,̓>�ϯ>�r[>Ւ��k'�Y/������
>�v�#�s��h�7��Ӿ<�)��ٝ�I��ɰν��ӽ�U��t[�@��2��QPþ�!�=��>��/>*!�>:��=v�>�,��������<���#	��-��5��c���U^���=��Ah���i����?FҾ�!�>c�=c';���><���F��=�	?Rx�=���>�q�>�">K>�đ>#	m>tt>���>7M>Iy�>��p=!�G���D���6��Zl��$0�?z���t>R�zC��2�Td�K�=b�>V�U>�u.����%��!��>P�ϼJM�ÁK>]&��z>��?��"������#">��F��=���3�XO'?��,>R�������c;7^��6?��?�/g�=�:|=EM;?0l{?W�??k!F�h�>;�>n3\>�ճ=��=��4���J��o�>A|q?-Y?�?@?��Z=t9!���m���E<c�q�x�<�$)�ز�eb��~T=̔˽�F\=y�v��ޙ�f�
=+P���1�=�0f<��;�>�Ok?v�%?��!?�r��&9E��L������m<�3��� 3?��?��O?��9?�/7?���>Gى��WԾ�붾���>N�=��;�?�t��0�p�z>�>[K@?HU?�r��/��M"�8�>�hq>��%>�?��>۝d>��6>���CSѿo#�������sc��ۘ�����<`q@>�5H���l�+�ǽ|\罉��=˝�>P��>m�<>/ >�$!>{�>��B=���=��>o&���ӽ��<�^(�q6�����e[���4=�=>E���sw	��1[���9����	|��?��?����ዽ�T����=��Bi�>8��>Τ�>U2�>p߷=-c���U��iA���H��>��g?�� ?�t4���=4�K(<�8�>X��>�>\�W�������b�;�N�>+N?��>�X���W��&m�\��h	�>b=�J���?���?@����z�"���U�+�F&
=ڣ�Lｏ}�����'4�_
���G:<�W�k=<��>4D�?�I=�4A>Zى������>����䁾�R��?���>�ˌ=Q,����!پ�T �9�!�1:���=a�>�6?�1?��L?�?��?:���� ?�n�>yL�>.r�>ַ?��?��?�ũ=o��=7'佐}�=�����;���s{<;k>��!>�G>�6^>�4=o�߻m�R����A9���U���=A�^=��(=��=�@>]�>���>s�+?�V��0w������g����:�+=��<���=��M�X��h��>B�?���>���>	�`�qv��i�<���5�=�e+?�t�>}�>?�R�>z�'>��!����H>�t�>}N�>��_�����;����`�>7y�>�ۯ>=�c>?x�?�T?�2?�α�P.%�9�m�
<��쎽ލr=!'�>��>,�M>�$N���@�m��^���4�����*'�2^�� �=�L>�`X>w�?>�o>��j=��������r�V�B�̼���>�u�>�"?zV6>d�d��������U�I?�^���`����$о2���>D�<>ۄ���?���I�}�^gR=��V�>���?n��?�5d?�HC�S����\>I�U>�>Q./<��=�������{3>q��=$�x�ɕ��F�;��\>O�y>>cȽ�PʾQ9�}�I���Ŀ���q�ϾdM������:$�������>¯�������,��u��e%������0����^���܂��y��
я?�_�?A=`��z�
�/��k&�	�? @���E���^�2�&�Sj���������0���оH���?�)͟>՗I������u���6���;��@>�w0?�ξ�:�����O7���>�2�=�/�/\��~��_�4�W�A?�6/?׌ݾv�ӾC��Ó >��	?�9�>�٦=Hi��V�$��ԑ>��8?��6?<|��� ��+��R��;���?ٿ�?�A?��὏�(�ݯ���h�Ej?��)?���>�(&�_�ӾG돾���>��'?��>���X0��.1��'?q6Q?�j0��>#Q�>�(u>w���yJ���ȭ��{�]�=��W>���<Qս�kn��Us�>`��O�>��~>6���-c��N>�pǾ��X�'�F���)�����c�U?X��C�o�+�>M:�>��%��1��/~x�����\�??;��?��>��F?��3�z������z��I >� �<�>�>e��Mc���f�>䈘��Ff����6�?I��?e��?ȫA?�'���*ٿ��������Д��kZ�<�}|=��G>Cݼ\>�-V=� ��>j�m>.�n>��W>�$�>d8>ɺp>w<x>���c,��ҏ�.�����9���M���I��p�_1j�����3q�����4 ���D���̽'�)������v: � ����=���>�=�>��>�e>|�&>���fؾ�4���?���8�θ�/վ� ʾVSξ�+��z&�w#x��.��Nپ�>���=S����>�m���%>Cq�>i�Q�s�>==��=�>A�M>
�W>�Ո>q>��=�9�=VÌ>�.i=�䐿Q�S��M��qVɾ����r�?�D��%2��f侓v	���4�~��2;?�K�>�~A�Q���0��]D�>�g��7|i=6�2>�����`�>��?�罾t٤<A2�>�������^h>.!?��u>�=��y�'�T�,>-�?\Y6��)>��=E=8?�w�?��A?)��62�>��>�=�=�!�=��>E��=��4�h�?:tW?�?S�3?��=�����5�f��a��iT�	-B�!s�=g��b�I*@���4�#�{��۹�L�t>E�=��%��K�;��>3|g?h��>ͯ>�L��a$���6��d���	^����p5�>��>�w?�@?@%?ݪ�=�N9�^��������>R�0> jE��\�@��=�R�>���>�6?��3?\{��]�n��~N>sz����>|?#?�y?���>_�|>?�û�����"ο>�⾉��~B�����?̽n��=�������p��Y𽽜푽Yx��ז>)a�>��	��v>�>�9�>�(>z���eJ�=B�=�����Ѷ��E>U7n�*=�Ma=���m��k�&��&�='wϽU�)�Y���\�V=S�$?�X	?J�=6Vh�	�<䛾�`x��7>�Q�>
?Z��>pu���*�&(X���4�r���ފ�>�;?�R?Sm	�� -=V_�����<{�>���>��>
���[��E�3�6=Z�>�?�2P>���F�X�'P�����pӇ>ؖ{=L����W?�?~��J��Sa.�MS��+Ӿc�=�52�l�꽞�Q�z���Z:������)�+��YA=��>���?Z�K�!Ƶ<�N���������`&���L����=��?.Y>
�)��w�̿��XҾ�v����;��<>d�h>��>\p?��>��a?:S#?�"?\k.�/��>	��>4Л>���>Ρ?��>�G�>qZt>��>�١=���<hZ��]��?T��J�"��<'>%:n>�S���+>n�>���=�`ν}h?=M�=`����7>�!=���=�%f>���>�"8?�0�=��>����W��v=нw����>h�5�/;��כ��'��>Ʒ*?�J?^r�>��<+")�B��E�Ⱦn�=��&?��D?��"?H��>��<	��É<
�e>NB>g��>�#��a���
�����>���>(.q>Q�b>�X�?.62?+�7?5��0�,�L��~fM�8>#�	g���?�*�>5 2>�FZ�� �N�^��z�k�5��j ���:��Gi>[j}>((�;�5>)���,<�l�<"�c�h	���>���^ѯ>l�?�+?���>���Uj��
�-�I?b/��%@�]���̾t+��l>��A>�	����>��w�x��R��m�>��l�>�B�?�i�?��`?�B��/����Y>$V>��>�<��7�;��qW{�5>X�=Q�w�y�����w�@>�7v>ͧ޽��Ҿ0!�T�d���Ŀ���`l���㾤w�Ձ�2���a�>߯����:����Lp��+f����g!p���뾬��Y�{�uf��	R?�>l?�5�=?iC�� �����#{�a2p>O$�G���S��-����3�Dv���E��)ӾB��;���g���>�2*�P���y l��d�t<�B>�1?u�ؾ-��-澙N%>��=lE�=-��E*���a��G��J+?v�:?1m�H/9�c��=��>N�?և�>�Xa>˂��j���>�\?o�?C��=^���̪��5ѯ��?J_�?�<?�=J���C�M��]���sm?�E?{a�>/s�����1������>��?���>c�������Y��>��Z?Z�N���0>���>�P�>u0!��@�� ʻ�|�������=����w��,5�!���=3�>� �>Mi��[���>9�5R���U�C���f��M�:F?>���=�=�)!>���=�&@�<����D������kI?(Z�?9�:?y"B?Ծ��	��)'�IϮ�ǿ�><�>V�>[��Z�>W��>�پ��_�5����?҆�?s��?�`D?�[���f���䑿����f�Y��v�>y]>�q8>���m�F��;�c!��_=|>}��>�&�>9�>9z_>�"i>�K%>;ƃ�$�����>��� �L)�Q%���XM=���ݾW�3�Yڦ��t�������;'��� �p����|�zz�#�*�Zͧ>�+�>i�<'�>��F>ħl�������5��޷��7<�&��z�ʾ��
��^���p�4qc�B ��-򽦡���(?��>�>�?�>�Q�֌�>v��ߴ�=2o>���<�b=�%=�=�Q>��>�2�>�Ǎ=^�w�Sq������M������=�����?"����?���?���&�X<	���X�_�>�?�$)�[-��>N��d �>����v �<�ri>�me��6>�z�>���dź<�s>�+,�l������>}�?F�Y>�o��'�о�L��x��:�=C?�p��2����%/?3l?�,I?g�ռ~��>oM�>��B>h�m>�
�>a>ؤi>5ê>}�]?�Sd?�C?<yV>�V/�Xx޾)�<wWW��E	> �Vߝ=t3�=��s�����B>��8>"S��ƌ=�"����<\��Q�� ,�>v�e?/�?��>!���PC��Qz�99���{1>C�{=��C?\'�>�}�>�$?���>�k�>��Z��hӾ����0-�> =G>�VQ��~9=�]�=#�>�>?��?̪b:��9�3v���۽GUM>OF�>�?�1?��>3 �=���.jӿ'$���!�pՂ�:���;2�<���M���^8G�-�1���lf�<��\>��>n�p>�E>��>�73>2M�>�6G>��=��=SF�;t�;OF�`�M=!����F<��P�ջ����Ƽ6y������J��>�d����ؼ�?��?��<������;���籈����>=��>���>U?�>�=����>M�T�H���-��O?�-o?1��>��#��L=Z�7�JZK���>XR�>C�X>�W-=U�	�t���w�k��S�>��?��>rp�E L��d���Z*�>�4g�^M~��{�?��?�d��I�7���R�F�ᾶσ="���`�o倾s���W����$1���,�=��>z��?WLO���5��"����FU��	�Ѿ����O>�4?��m>�fD�>т����-*������ˋ��Oi�!�N>�o�>��?�?!PP?.�	?��?z�r�#	?�>�A�>  ?��!?�?3�+?�p���Ԓ>��=J�>���2�n�
I�<�i�=s>R��=�R�=M>罒P4=">3]=W-2�����}�<ԻѼW�|�>[<���=S�*>L}?�A(?�S:����j���=�>E�����=R�U>nw仨]���q<�}i>�!?+7?�>��=i�߾�߾X�ﾤ�=��?�?z'�>�AX=?�/>h���1���>R@>�t�<�[h�)�������C̩>�m�>��O>��/>���?8=U?��*?��*&�#3����A�������<��?54�>�&~>�a9�Q�!��UB��p�!�.�聒������=���=c7>On8> ��=���=1�=�;�h�׽b�=l��< 2�>5��>߬?���>@�I������p�I?tn��[U�/���<Zо|����>��<>`��s�?>��,�}�����<=� r�>��?���?'9d?'�C�����\>0V>,�>0n.<�>��P�������3>��=�py����j�;��\>��x>cɽ��ʾV��J+H�Qmҿ���&Ha�@�پ�X,�r��iپ���=9�뾾"��&5��6�Y��.Ծ�U�K�8��Y��Zf��
��0?z?P��?��&<Fj���Y�Pf7���ξ�9�>Z��iV�����C���Ɉ��=�5��L��a���]��3C1��U�>��_�sE��2ct��X0���I��'>.?/wǾ5u��0��:�<>$r�<�
���x���js,��^I?x#2?P|��ܾY���%>f%?1��>���=K*���b��|��>U:9?4D/?�=��^��y{��Q���X�?(��?�eA?��N��3C�����Q�,/?~?���>����t�ʾ0q｀l?�:?��>����U���,����>tr\?w�K��`>ƞ�>�Ӕ>�i���c���}!�堐�����>06>���F��bg_�a?��̠=Ф�>D�{>�]�u�����>}j���Y�V7[���i�F��Z��[_?*����=}�=��=�c�� ���Wս� d?u
�?�/?�E?�?;�~�b���Ό����> =|>��#>c���U�7>�'�>@�ھH�J�iC�~��>�h�?g�?O.#?����4ƿ┿�w��ip�����>��G=9�>݂�h�=�Yqv=���=9]E=��9��)>�ְ>NO�>���=Ù=>��b>Z~�s��u���Om�����:����+�0����?þ�%Ծl����)�ӏ'���	����N���N�K��dP�������>*�>$�>���>��/>I!>���®��Z�m���� �;����ݾW����o���X������N������׫ܾyN?�#�Փk>E��>�AW��&�=�,�>8]�=jT>Xә>�*>��=dL8>��>`�8>�QO>�$>\��>�,��E��[ay���t� I��`f��V{?a���t�=�d�I��b�������;��>��%>7�B˙�n���C��>�C����n�^\�>l6e�
�=(�?8e@���T�&��好Ml��>_��
k?�I�>{����
�"�ɾ���I��>��ƾ+&�=y�D>.3)?(=�?O�a?[�����>�4�>�m�=��<�->>�c>��>�>�RD?�PM?�+?�
>�{�6�>%T>�b��x=������;ՃŽ1I��Q�O=���;&ϖ=�½�:��c>Y�����=��`>֬�>�d?�q?�%?k`�d2�x�T��\ʾ�G>��=��?K�?^�L?�?�>w��>����ꕾ�ƾy2�>	S*>s�D�Pqp�z~�=ϻ_>�\�>��,?c�6?�.>�n���M>��<C�e>�?s/?���>Rہ>
o":[��m�п%G�@2%�z�=���ZӐ��$���LG��,�֡���q���^5���=�}>"�>�=�I>m�>�\�>�^q>�}<���߽�����<�
I>\�E=`�S���P���<�@��"�p�+��P����=ki�=�D�>?9\?�m)�4��*e����������>�7�>6�>��>;#�=bm��U�v:A�ZmG����>׍h?���>�7�½=Ğ0��ȁ:�³>$ܡ>\A>0_�$��ٔ���d�<%h�>��?]�>���".[�Z�o�\�
�P��>k�<=@�����?��|?�A�3�<����sO�K\(�{͂=�c�=�1w������:���Q��Ⱦ���TPL��_>G�>��?gۅ=�_=>��]��%풿� ۾O�d��ap=��?:�>h[A��j���m��0��s����5��� >�À==��>��>V"�> T?C�?��/?�]F�� ?���>Զ�>:}�>N<�>��>�?E�=��>��ʝQ=|�ս��Y]�<{��=��=!�>��>�c���J>��=�����`�����#>��V=�U��{�K>ț�>�b�>�
?@�?�齠����;�\�)�>L�<K�=o��=�c�@e��0����nY>��?\�)?��>��ü����Y1����+)>��?z;?�+?�́=$�=�p�@w��>C-v>�P�=�<E��f��O����K��8�>ru�>g�9>7�r>�҃?�Z?3�9?p��q�2��ir��&<�h���ź�Y�>��>��>B��K�?��Q��'l��x'���̼t�a��=�f�=�C�=
2!>��]=�D�:q�;=�C�<�1�* 3<�+=Ʀ�>�T�> �?�>N�m=s���%�AoG?����x��4����Ծ�"���>!�S>��>]X �� z�\j��OOB�`��>���?�_�?dM`?,sW���� �Y>��F>�>�H���8��v�L�R��r">Ӓ�=��j��"����G���[>���>�e��o(Ծ��Ì��ҽ�i�P�݆b�����@�k���rǾy�=��.�P'�EY߾��n���k��P�-��:K����!2�eG���?t�~?�è����NI;��� �Q���K�]>e��� {�����:M���m�뾳[���M�i[�u���J.�w��>}e�<m��cq�#K4��VE���9>��*?��ξ66�����wӼ>&^=]�2���������3�>�D?�_0?�ྶ�Ѿq���$k.>�j?�E�>�U�=ӯ����b���>m�4?�55?*F��T�����b�v���?�l�?o�??�pQ��S@��x���#�S?p�
?���>;a���I˾���h�?�8?�<�>������ P��u�>�V?9R�ԍf>y5�>5j�>�ǽy������j��@ѥ��3F>irλ���W�AGF�TŠ=?��>�nx>�X�W��l�>v����M�xG�Dw��b%��S<�Z?�����>��f>X�>�'�/o��ò��R~��^L?V�?sR?�8?6�����yƴ��w=�Ǫ>� �>)�=����a�>�E�>R��]r���_@?��? ��?�iY?��i�h�ܿ[֏��ᚾV4��FΝ<��=�3>��=H5>uW#�,�(�*��
�=�e�>[�h>��@>��=�|�<�
*>ច�%�!�;楿K��$�,�Ӿ��,��gʽk�ǾL��JP�D�ӾQ����<6<7���@��['8����Q�콃�۾�S��I�>/�>��?����t�=�8����O��'`�������־����@��h*��s�V�cs��'���-x=D����>ZtK>FΈ:EA
>nX�>xo1�D�P>�0����>��5=`�߼��q>!d>��o>�z>P�>/Q>��>x��=�fp���{S�d�*���,��4N?;q���x�xy1�75Ծ9"���0L>z�?M"�=h-�R���y�x�ެ>�T��?e-��~#��*���u�>���>�q�=��;��½<M��'���P>�,�>�v�>6�=`�����ͽ)Gm��ޓ>�j�W�@���h>i?@"~?v��?ȫY���_=�T>/�T?�@1?���>��ӽ��
<}?�F?`�%?r�>���=������<>���fȒ��(/�����Zt=�Xk=j#U>+�ӽ�Oe���T; �1<�:�����<l6=�]�=��-�>+T?�B�>_�>�Az��M�3D�W ^��u=?FǽZ$�>��>�U�>ŉ�>l)�>� �>�"=�tľ�����>G�?>�uS�?f~�U�&�$�>�r>s4F?ub?.wA��ި��=/s�<���>�A?8�9?�:�>Cx�=���B�
�Y;Ϳnq1�P�8�e��<E~0�t�-������u�;(A>?#8� n�r��<�	�>��Y>5KN>ID,>�>�6�i=� ?�Z�=����\�>��G>��7=<�K���7�x����p>���t�<���0��0ܽ�Z�L =^�׽�ڽ��?��/?����(>� ���ؾ	y��N�?���>a��>�>�Y�=�����u�4)p�{�l���>��e?���>kge��T�>χ�=]`���Z�=��$>g<>�<����$��Kq�u�*=w?�nJ?%�>�@;�sv��!��1�Y��6?��=�\�觘?@�j?�3�=��� �'3������(�Ύ�u&���(;���g ����
qԾ�~��l�>��>��?��V�B`��R��C����������~i=І���>�>_žj�ʾk�Ծ{�����=;��_/]>簉��`�>�f?k~f?�3?-16?S�#?�Rľ=�4?�1�>P�J?�?eG?��>[&>�����)��h���n>X� ���依����hѽB���L:���=�r��,�I�M���S>�=�z
=�s=*�=�\!=��﹢�i��P=?(C>��>��\?�u>(���u����J=�����	 ?�g�>�<�>��Z��3����>J�
>L��>G�~>'  �ߣ���eO�P�	>`�1?��]?�v$?�>�=�0*>�5�|�;>��Y>���>�I"=� ��g���{����=޳�>z��>��n>��>�@�?JS ?�j�>|,��ο ��;��� �K��=��>Wy�>�x	?ã�<������g�:V��o�s�9�:��:=!`�<��3>�:�`�*=�K>���=���>���2�͖�����׋�>{�>I�&?�a�=��]<Jv�֠C�-L?:�ݽzȊ���d��l���V���׾�'�곈:�M2��T������I���D���~B?z��?���?�	?u
��x*�=���=EK���= 4=��>G*�=B��`�>C>K�<��нg�����=NW>������M�:���̻�+���q���ܾ�4��֩x>���\�yb=���>US>�E׾*os�链��w����{���~2��ܾ<�?��V?�t>��ݼkﾝ��=۾mĶ=�����1�}��KQ��ϖ�A�پ�l��;Q��"¹�\���蟾ߤ�>�?�����'���-�2���^>>��0?�o=��羶�K���J�a��>6�?���=0�X�m$��0q�<`�?�x"?x�+��R���w
�;�?13?#��>�E>mo�+T����>�1G?��?��>ҟ��Bz��-C|���?�ՙ?�~Z?�v�P>�J�"�� ���>]�>֡?|��m��7�P˸>�ȅ?|Q^?���'Co�Z�2���r?�/�?h����>?(�?��?����`ľ�!B�2愾��w�:5�=�j>��O����v�
��@���Vk>&�0>�\�����{>�>��׾��&���_�f�A3��``���;5?�m���M�>��T=C�=T�$�p��Г~�DЁ��dA?KN�?e�j?��j?φ쾟R˾ ��I^�"��>P�>؉=<��=E�L>�`�>8�(�
�{�o��I�'?<��?�H�?�WM?��E��Կ�����Z���=�J�=�qB>�#�评=�=
S�;Uc�Fz�=NeW>�B>�b:>�$'>��@>���=X!��$��:������8P8�i���v� }�����w���v�9�߾׽�@��@'ݽ?`��n�2��e$�	�f��A����>��?��>�0>x�>�hU>�n�����:����w�?���鰾=��e���eU��Ԓ�⮾���������>[?�=���=Bn? �=��w>t��>$��;���>� >���=XS>Á�=�'�=V�>Oi~>��%>�K>W��<`���r�~�����we�X ���O??�LH�vX���p;��*�����؇>u��>�2W>]I�Jȓ��,m��"�>~ˉ�BW������<�;	/g>5��>�> ]+=��������s2��Q�=;��>p�>u
���ň�b6��y�=+��>�k̾���=�6�>��$?�Sx?q�8?I��=7��>�f>�_�>��=F;I>fwP>�>�?�2?��,?r*�>���=}�l��E�<A�A=�;�d�S��۴��/ܼ+�4��P�;��ϼP�r=(�s=�<��P=�g8=������;ݍ=���>b�7?�>���>�pa��8�X�N���E�ݑ�=4�E�NK�>B1�>Ź�>�O�>Rp�>`3z>U0�{S;�V�-}�>��8>C\\��Yj��Y��,�b>�.�>�WH?�:?�O�<��c�)V�<�'�=/+�>϶ ?J%?���>�->��I-��;��#F۾R4��[ =��E����Ծ~y�L��>݈&��5���#ƽ���� �ܽ5�=���=�6*�5��3�>��Q=1�<�=�)>�͖�O��	ڝ�j����ZM>G9���>����������x���Z����p�����?�$,?��<)��� �����i'=��>��>"��>#�����)�ʫm���c���\�~?
�c?o?�Ⱦ�b}>yS���n>`�=�>� �>t;��懾7^��]��>�+�>��)?�">�DC��r�����p�^���?��=>)�=~�?��F?��+�mv��*���*��'�R�/�8�
�ƺ��ҫ�w��i:�Ѹ�M�Ҿ*%�z�t>�y�>U0�?��&��>U��ٝ�������۾-q(=)��<I~�>�Y�=Zz��f��;�׾�wϽ:�ݼ���;�	�>�Y>==�>4�>m<?�2?'�k?C�N?sq>�=?�u>P��?���>*�>���>���>�=�=j���j/�=
��G���F�$����=�\:>P�X=�Q�=�)����Խ�� ;jف<���=P�<a�{<�4[=��c=Ъ>&?>��<�#?�*?b`�����~d��>-�L��=���==*��Q���LI:V�O>[?�M)?']�>S��=@���rH������E>"?n�?W��>ˇ�=&<�=$�ľ&'A�d�6=�>FX�ok��H7�Ⱦ#1��f>��|>�_�=be�=���?�!(?T}\?�|��X_��}���)�'�y</����<>v��>u��=[E���2�Z*<�����'7��/�;=E�����=���>�����1�=3��>�@�w�>x�3>��p��aнMv��v�>~�?$�?���=P�
�������@]?��B���������Oѯ��h�V����񑽕2>r+�~}�a}���y��?P��?Z�?zJ?2u����=��=0ɰ��Mּ1�^>��νS D>������>��>�3�=8Z��� ���=��W>�{��Fs�|�@��+��=��9B��+þZ���L�>����W������	J�zG>y �wȽ=�Q��������C�����V߾�x��8�?��M?'�:=��;�Jv�����־��>�(�x�M��_��H�1�d����w8a�b���լ��ľ%D�NF�>����ି"������f^�=�{>ev??o�{�zJ���#�Q'�M{>79�>�����uq��v��+ùv�V?��?��"��	���/� �>&�>�"�>E>��⾸,�����>�\?c�?�i>@����੿�v����?o?tjT?�$�yX&�q��������8>�?�?�9�1~J���N�ށ%?���?0>P?6G������+Hf�]vM?��>_p���J?�:?�>Nѷ�:'[�i60=����y־�>?�z�5F(�Cg¾_U��Ϧ ����>Շ�>�(�6=�.�>g5��0:H��P�$r˾�
-�e�����>�:����i>vZ="׍=�.�me��9zx�֯8=��f?
Ф?��=?	*d?���h
�N5����[�;
�>�~�>�Ų=�}^��\>ZZ�>1a־��|�o#޾Ĝ+?�T�?4��?�\?��h�'�̿d���`���"����_�=3�	<	>���R��<�\k=f�	>uC�=��a>Z��>O/>`�v>��4>譣=~!z=�7��d��Ң�AS��<�.� ?��z5�^����i������:���.��0������.������b{����O8.������7�=��>�3�>��>��=��*=��V�g�پ��~� ������-���8���b�־��d��ؚ���Ѿ�nվ�ۆ;��ž�?�n��*VE>8E�>2�7���t>�̵>.�>l7>1�$�C�k=+�=굮=��o>��%>~"�>E��=�>��Ҽd5��'Ew�:<�#BA��M����0?l�5�Gɛ�D�,��^��"J��8�>
M�>ѹ�>�=��f��L&e�#
�>�a�����k��o�>�z�>�  >�4���_����{�_*�4>ە�>Dj�=�ٽ\����9�c>2C�>7�Ӿ�H�=1w>�o)?]vy?�:?I�t=(/�>�Tn>�&�>��=��L>tnW>}؊>�?�j6?��/?���>QF�=�~e�8�M<��*=�!6��37��5�7��g�X)�<2�>��dV=��=�x<
�=^�E=��伸��;�=���>u�4?@�>h6�>�J��=��Q��>�F{%>�ȡ�r�>�8�>��>�x�>�G�>�+>Y�μ�
����վI�>�2d>�a��}��&��Jq>@z>�{H?2*?݃��X���{�==��=~Й>���>��2?�8�>�Y?>������������j��s{=@�n��=b^@�ѣ�<���rh���ã��D>@>�m~>Pn�=��5=K=��>�>�<�>nd�=�90=	�z���U=�Jl�ݜ=�^���ռ����8y���4�
��E]�'�=�;H=�0?Q�?oĭ=R/�cᲾ��@�<w����>�e�>;v�>U�:?�g;>�>��I^���D�P���X�?kw}?��>?�2L�(Y>��Z��y=���=�]�=}���昼�m=0�"=ZÃ>g3?9��>���>�Ľ�r��w;z���8����>�=���P�?_fj?�F�́��l&5���n�w|����1��c ��ƾ3��a�#� e�˺����	��B>���>53�?Ͻ0��d
>���5����ǁ�|����ڇ>���?�>m�>!�|��R���� (_����=�̕=��>_�佣�?ZR?]ES?L�C?��G?4Tl?v!\<��4?�^?��1?]d�>Y�?��>���>�>�k>�d�SK�����񊮾�	��O�W6c>L/�>4�>����>�v=�z�Ug�=N߂��% >��=��$=X�=�:>v��>��?���>�Ľs�
�d�����8�� =�n>d��6���¯��ʿ��t|(>�N?V'6?�g�>���,���G����ysj>��)?�i&?��>~��7st�#����K��=�$�>�d4��.��2�.�
���;�׮(>��{>>�;�c>�ޔ?%�!?�|Q?�
7���&�&P��j��W>G�;���>�
?��e>�����6��J��f�Z�;_Q�Gn���Ͼ�*~>���>�ٞ>W>�dY>�sg>�]��.;z�}Y�F�C�����?�Y�>8B�>⇹>Vג<��ƾ��:��uV?�þ��"�Pr��`m���U>7�u���B=0Ď<"(�>q�3�z��[����*�5��>
��?���?��S?�����\=��[��l�(N�=w�=X�q���/>>>	��;���=��B=E���U�w<��?�?��$�Em�X�n�:>����]5��^�	H�����>����m徠v��p,'����<˾�>	_5�E�m���@�d��?��Q��K�$��Uf?�I.?=iW��3��n׾��ƾ���"�N=�u@��k��b�Ѿ��M�Y�%ܭy�:S��N̾>'C��Һ�>Ǝ�埿CU��j����=��3>�5? u��X����#�f�ٽ�g>(@�>:K���T����̽�K`?��(?��ʾ���i�W��q8��s�>��>}KP=�̾��X���={�'?A�m?]-;>T��_��!lt����?깥?�HQ?�꾀0/�ٛ/�o�1��I?��J?�?�>)����2���W>��q?%*W?5�=��b�����	?Ѻ`?Gn�Z��>s?��?�猾��ƾ\�<�wP�p0<�i}E=Fs_=C� ��q���{��S�N>b�4>�5�Ν�k��>��ӾF��i2!����Ҿ�Y���?�Ͼ�P=��V<�\�<*F�������t��M�<��K?a��?)T??f?�羰3��[�+s����>��>��=2�N=�O�=�>x�'aN�MHѾ"4?���?.��?Yw?�É����❃�Dl���Ӟ���W>, ^>�>�5�P><��=D���d���#�=�>�`.>%�>wz*>�K�=#
>�x��P8�'&��aΝ�"��Odݾ�I��F�����6н�<�r��������B������3�hBz�B�C��Ֆ�_�_>��?<!�>��>�H>� >�;���cľ��A�TI��������׾]	ƾ������p�s*���;��"mͽ�����>�i3>nm!>�w�>�t��G�>>
rS>i_h>��6>z��=�1>�J�=n�O>JRw>�,�>��`>_:�>c������ڃ���:�-K���;;�B?%�U��]��}7���龱O���K�>P�?���>��"�H����hb���>��~�b�O��*齕�����>���>��=���)�Ž��7�Ei���0O>�-�>W[$>^�8q��"Խ���=��>�zϾ8l�=���>��*?��u?H�9?W�_=�F�>yO[>�ɠ>>��=�6P>=Z>�8�>��?��0?�l%?H��>Cz�=&r�6�;���<�lP�K�a�)ʰ�κ���q�ƕ<lK����=y��=�/?<���=��q=�q�cU&:?�*=6�?M)?s��>q��>�t4��=:�,mQ��dq��>l����>��>�V�>j��>�]�>�-�>�.�=�����6���j�>;}+>�ft��v�ӴL9��z>q4l>yU.?kM4?�
�v_�����<�݁=ɷ�>�9?��7?JS�>��L>�%����￮&��+����m=��$>��Խ�4ܾ�����Q���>hQ��Fb�:�&����4>�����=�m��w����nF����>,I�=�&�<H	#>r)��&:|��q軶��<G+P=7e=h�����>�XF=��`��!����I=t�V�\�Q��7>�51?��?�8/�g{D>�T��5�b��� �>
2?�^?�S$?c�>�Q�8i���Q�-(���|?'Aw?	2?+���f��>�3>4̓=���>� �>��m�H+��ʛ*=1׿��>���>� "?�>�Q��,�t�y����.D�k@r>�Ό=�$� ��?�d?�7�r�&�'�(�"�G���}O��{/��ϣ���ľ��a�9�A��/?�MF��&y>7��>��?��R�Q�/>����e/��En~��э�-�<#��^��>%�J>N,���P����j����<� >qE7>�#e��7?Yg?C9@?n�i?ۘ{?%}?arN��W�>��>8�b?=?�)?b�>��G>��=7�Ľ��{�V-�=����:�̾��6=�>)��<Y|>�S>��<�Jս��7��,[=���=�%�<f9P=ӂ?=u��=�~�;E��=k7`>��?'H?����m�ؽ�签Q�F���=�+ >��=�,�ҫ������4>��>��?�=�>�˻��l�-��d��*��>��/?�P9?qF?H��=�S���*��Wо/�Y>]�>"��^���rN����U���U�y>��>\6>�td>ٌ�?Pk?�Z?�*�<+V4���%�V���
?>3٨�$ƪ>���>��>�� ���;�M�� �[��)<�q�龏����_>\V�>�F�=>�� >r �>aW��G�#�[Z���c罛w|��]�>���>��?!s[>�̼|2�*�&�e�l?�wž%)M���|�±�w7P�5G@���=|G�=��$>�C��f�N�L���0��/�>���?{'�?��|?.+�����=���<�ܓ�X�:;5�̺�e�?�>	�<>UG�=��%>�c3>�_̽f��=�M8>��>�*�n����mS�3zY>妶���D��[6����~�=��z��2�нʠ�u�>|�����c�����ˈ�9|�TR��t���Ǔ�H�u?�DJ?�%�<��k���	�^KA�ԛ�>3�>�Y���Ͻ�F�֟��ɾ�1ľ4ے����>`ɾx徙QѾ�M�>��ܾD��lT���(�n�V�BY>(�@?j*�KG���h�����>o1�>���O�V��X��zm�<!}_?K�%?뜡����6ཿ�9>��?
v�>}�>>c� ���n��5�>�?�4p?��>�僿|��q�.���?S'�?�Z?� �CN<��2�M���>i�1?*�Q?��ξ�K�=�p���=vψ?��\?��H>��a�u#5��6G?1/^?3vd�[�>�.�>Q��>��澏S��uX>��:���>�w>�p��v��qa��t@�+с���>��>IV��߈����>cپ�x>�F~.�tv��þ�7���>{���Q�=���=�\9=A�Z����s�AG:�N?�˙?�y2?�:c?|����2����Ԥ=��.�>e:�>�,/�����J�>�8�>�
��b��,��$?�?�?6�?h�J?��H��B���Ӄ�C/̾����}�=�ш>ƟM>�q����>�>G�b=��5�b; >p>�-�=�\H>LE>�>�=��>��<w���������Q�6�EǾ#��'�仝-��*�ؽ��:�SE�,*��,���k�m�K)j��L4�D�z|=56��%�y=Z=?�)<F�>k) >t�<��r�o�-�ӭ��0P��EL�?�׾�������֨�������(�O�����,�����:�>��f>�����>��<���>Y+�>�&���>�Pt>�mx>M��=7,>^$=G�
<��=���=%2�>�� �����l��� �Q���]5�=V?%½����8T:�c@������ލ>�A?��>+s8��8����-���>Uw�\���p0=jEQ=�5�>.��>a92>@�;�N�Wo��H>m5{>q�>�e>�4�*�뾗�O�V�=���>� ��E�V=��y>-&?��s?�+?^O��t�>}b%>�/�>p�=��=k�<>�o�>��?��N?�<?���>E��=k:���<���<��
&i��8_�%�d=��
<
�p<�<�&�=�0=^[���ˤ<�=�d�I�=��$=h-�>��H?���>N �>��,!��k�y�/�kN>c�4=Ms?!?�>n�#?�A�>�Ӯ>y�>�d��A��\q�>�1>�M���c�/��=z�>�
�>ʌ:?�=?��*>��a���$�D��=k��>_w�>��?�z�>by�>7���"_��Ĕ�p�'�7P�`�>�^��q�Yٻ���>�Z�>nS۾�m��9B��! ��/�4�D>��=�9���s�����>��>Z��=�"�>.P5>J⯾��g����}�Ὀ�m���/��}=��2<�H�=:;�4��k������B��>$?Q'?�ލ�сq��a��3A�-���4ˁ���)>5�
?I?� |=&"���M��^�����9�?C�?�?�p���W>�@>-��=~�<�(>��~<�ܽӠ��|彡��<�>>"&?
߸>w�w�cg��9�����U��Z?F��=w)�}��?�4D?L�Y�H��ܻ&�\�,�����k�ᮙ�"=����oY���N��@����=��?f��?�x�� >��z������E}�F\$�zX�jY>���>0�A>HԨ�sΠ���0�]�{�I��=��>J�>b6�b�?u4n?v�^?�g?~o!?$
?���( ?J?�pJ?ܩ�>��K?Z�?��'>L��<U)'>0Ľ%����Y���ľ�C>���=M��= m9>��>�i������qԽ]�1>�Ķ=�Vν���= _u=m����/�">���>VD?���>C�.����^E�� ����=t��=ws?�16�=��BrW�Y�	>?uoC?�a	?���=A��� F��Lz��T�>�C?u*�>�?��E�vӕ��U�<r�̰l>�6�>%�K�u����,�f��A]�q�>(��>��,��>�w�?)?k�X?M��e�=�'�w��<��93�>���>P�b?��>��-�z,�����֗\�WFs���:�;Q��,�=�3b>\�\>#�>%i�=��)���Z>���>�渽�`;:��>1�?�6�>�� ?���>�{=��@7���b?	�M��0(��vj�C@��ql>;�;=�Q	�Br���.>y��=h�=�	C����+�;��>3(�?�h�?=�y?Z����?H=r�=�A=�p=N�9>Z�u=�V�=��.>̿>�O�=Bͽ#=�9�:/	�=�r�>��>m$ܾj{���=cp��R*/�P���J����A���7������=���� �=�����U��������a�UG@��6��3���3����~�?ߚC?�,���l�WbK�e����T'>�+��d_�R7�������5�NKþ?�����4����׾h����g�>Q���B]����d�O����
�	k>k�B?�*���sƾ�(��&>�S>��>JՑ��n�bf��.��5U?4�6?���-�޾ψŽb�P<1��>���>�8Q>jy��t�K�C�>��?�+?�@�=��= ��gm<ꋽ?�M�?�I]?$���6��M�6���Z?�{�?�uU?���"2X��O��>Jv]?��o?,Ep>i7&��3:�D=?_L|?�	3����>�b�>��=P��C�P���^=7�׾i{�;�<>�ͽ�M޾)�8�7�G��P��ẁ>��>�9�Ж�x��>|s2�/�A���\�M\ʾF�ľ(ʹ=_a?zD��)�>g��>��)>��=��������*���?��?iG?�3@?ˡ˾���w-ӽz�=�y�>0��>"H�B�]�|[~>� �>�s.�Bv��N��h�>�G�?���?.V?�ֈ�/1ο�����넾�Ǿf#�=�_n=�%>�A�������=�='�M=�2�=�%r>�h*>%<B>ߓ>t/>&��=����CU��5�������V�t�+��}'�yX��V��7(J��O������Pھ ����'�
2��σ��ӎ���e�=D�����>�>���>I��>V|�>��=K�ξ^��<��	q�[7������� d���M�����晾��I����M-��5*?[\�>�s�=	.?ʢb=T)���>�ܽ��>9Y�>��w>q">�w)��>>�?@>ܟ�>�20>
��>?�2=e����y���$�����ī=e�C? C���#���}?�{����N�I�>vD?J�M>�&��a��hAz����>����Dn�U'��Y�O�lQ�>���>;��=oQ�=;@.�����Uƽ��R=T>�>�gB>֩�=�3x��zB�&��=ڠ?���s��%��>��4?���?� ?R�.��
R>e&�>*�=LH���>q�?���>�%+?:s%?�?�k�>e>����I����=���ݩD�m�=�>56>W���B�?Ă=��n="n<",�ڡ7=�`=�:;���<��
?s�#?�6�>%I�>�S4��w��6@��B4>���>|@}���>��>�	O?U�>���>�OC��%��?+D�+(	���>���=>���<z�t��r>5�1?�TX?�D?�cp���F�:t�Z=m��>�3\?Z�S?qr�>��3���V��5�H���G�)�Z��Y��h7�Z��]�S<7U��N
�U��<�)x>�Z>��=�OI>s�л�]@��z�>���
C�=�c>1aн�Z�Y��=8�=�>=��=@���H�;f��<*}�8��z��<0������J�=��0?��>&��!r���Ѿ��G�=���?�*%?�Y>��D?jú>��sƋ�=p���{�>(s?�>?������ӽH덾XQ�>t�>��H�E�=ڼ׼�K���h�=�VN?a�N?���=Lj�ra��������?�;�>�=~�G���?`)�?�k��?;���	��mT�[v��?���H#�-�������$ ���&�7զ��[Ⱦ�O��EB>�?v3�?Odv���>#4�=���V�����B��=V�@�[?�>}4���d��R��W�6a�=��5>#�{>򖓾$�I?���?��?��?�1?�AV?&���3&�>�h����><o�>�+	?�}�>O�>�ң<#P�=Q$�:���
��i���役\/�c3�=��=���<�W߼3Q��˒p>,az=f��=��1><���\=�2C��M�=���>u�x>��?.?l�/�Kl�=±d����=Y�w>�X�>t!�>��侴�޾p߇�|�>W��>��1? ?~-�%�-�#�wu-�@�>�?X�6?_��>m�e<�=;����툌=b��>����$��bgԾTf	��f2��3>�������;�F�>Ϧc?v�2? �?�V��I�n)����׾q�=�� ���>�b�>�
�>���nR�L=���t��vξ|=+�$�^�9��=}�z>�'>C�}>H6�=%�>�V�=��B�i3a�E�ս��h��>���>��?��]>X
�=P.D�z��[6W?����~V�eAX�!5��
#
>��=J�����v$?�ɾRƌ�����i����?Y�?F��?L�G?N �=�Ľ?U��=Vz?�>�<�̵L�㫻�7���^/>���=��þh��c���I>V�9>�A���澦���$>��ο�t��։=�Q����&��������mo1<Y�6������8]�Gn7��9���������x��?�Ƴn?�V�>�U*����gվ���!��/�>H��D����N���^��K���ㄾ����n۾������M�ʙ<>˾@���W�i�~
�d��:>��9?�޾��z�T���]>v@>��O���񾳒����y�W��k?!�h?�0��,�����>Lr�>k�>��>�WT�=0=�>
�9?��?nյ�x��s,��n�H=�S�?���?�E?�a1�p�8���o1T��D�>�>h ?�w�-��=;�O�(?�eR?g>'��J����R7���>��N?�pg��z�>>H�>�ʡ>vO��}�Ὥ랽xd��j����,8>���D��ޫ^��}U�pB�=й}>�J9>��JD �#��>+���2�]��W.�������">�r�> @"�ϝ�>�c|>>��>�\8��h{���!�S��t?
�?��f?47Z?��
�����Y����:�>�l�>/%�>���<U�$����>� �>�׾�Qo�� ���?��?\��?��M?��d�<ſ����և��[>V��=�Ϊ>h�K��'��sE��ڽ�E� T�=v��>!e>�x >���=C�*>ᗓ>��}�b����:c��@ <�����3�ݜ9�[�+���Ⱦ'p,��+�z�Ⱦ�z3=�����5�Ad������[=֖�29�>q&"?�Z�>�U�>s>�>��>*�߾���qҷ��!ʾ�C#�<?�V ������B�����^8������8󐼬��$�?/,j>�>��>�>0_=�>�%�=���=�l�=��=��2>�u�;�;>{�T>է4>�k�>��>'{�=̂�C�{�,�-!��O.=?�I?�V ��j���~5�B¾�N��v~�>��?�%Y>S�*��Փ��}����>�����9f�uѽ=v�[��>c��>叅=�l=_C��~�3R���=�X>��.>�_�<2����o��%�=�>U�پ*��=�w>̗)?cEw?&�6?+D�=��>HRg>�)�>瞮=O)A>� Y>���>�?Ӆ9?�T.?�~�>;m�=f�Y���=$&<=�NM�.D]��꨽�Ƽ��j֒<��Y�!�9=^��=��<�Ev=ɠL=J�P$<�5$=o;?�!4?���>Ga�>tmb�� 0�'G/�i��>E��=1f��>�>q2?ۜV?[~'?L��>���1��h���̾y_�>O�a>Z�$d��i�w��>�>��Q?0�Y?��ؾ/ݾ1�>��(>�
?ެ#?�I[?G�>p�=���j���F��U$C�չ�s
3�)`%��!�a���P��;r���p��F=����=2�v>Y�>���;(���T�v|8>u��>���=<��=����"T��S�<q=;Nvw=���=��>�]�=�8>J{�������^|��Gy<�I�Hw��T3?��>�-i>q������O8��+����>;�F?��E?�`n?���>�Ⱦ�]��zV��m�|�#?8�?��?���|���-�<.c/=�ц>�v׼�.>څ��ĉ�+a����=MO�>70<?��>�Ƚ�jX��3���׾]>6>86�3�?�[�?����㳽2 ���M�6ʾ7{=U�N�J�Hؾz
���!�'�Ľ�*������Ȍ�>���>��?XR��� 	=�C���c:��1j�=A��>��s>Ͻ-?X��=86�|q��n�V�h���(=���>R<�>|>.��?��Y?Ύ'?&�{?K&>?��9?����#�?.Pлp��>u�>y!?2��>aS�>2�=�u�=��O���u����ϐ�ӫ̼�,=��=�>���=f=&:���=�%U=�7��:��չ<=�������N=�M >�N>sA�>�Pf?�f7��v �V8ӽ�Z6>�V=0$b>Z�>�M�����k<�ޣ>�6�>&7J?�w?��9�2����Y�'�p[�>Z�?�H�>>��>D��=�Hֽ���%���3�2�Ov>Эo�ԍ��ξP{��������=��Q>�􁼓��>CZ\?ߊ_?Hf?������_�ȵs�K�־SJ���:�=�O�>`�>��>2�;������dM��r���}=Lb8�4jT>� >]ώ=&J>[�>�^=�H�=��9�r߇���KӺ���>5�>�w?wJ�=�`;��۾>qþ�XZ?=a3�Mt6��/=���0>��K>�Y�>| G���Y�9#?��=�Dv��C���Si���(?���?Jĵ?R��>
/��;<U�x@�>��z>6S>�\վ�����m=4�&�>�}ռ*%��<���� ><��>��>�I=9 �x�Ѿ�/�;����4H����5޾�֮��[о@�⾲BR�m���]C���۾բ߽^LX���8����X��כ��0ľ'!�����?,N??<�={�<�
�]5��S��2�+=3@��s�<�el���%=�r�<о�AӾ4�O"�6��\�㾑�z>@������2�z�S���˼ݑ>=�?�پ�b����(W>�O�=x$��6������F���!��UX?�K?�Rܾ-6˾�bg�?s+>/��>3h�>^�U>�ޢ���}=��>L�=?�$
?��ۼ�p��0{��nk�=t��?l��?4A?���~<��=�AV�/�?Oc?/?T9����x�A�Ki?�"L?��>Z�޾2f}�l�)�/�>�:7?_"O��e�>�ʸ>��>�ꗽq�e�ظr�,!��;�|=�9>d��~�	�+�������H{>=�>ٟV>�4y�Ů�'G�>T� ��6<���m�ྻF���H�a�!?�Q˾i|�>\<>�Ě><$�8w��c���Vj�+�e?ܥ�?��?��n?�����þ�����>[8�>�ނ>���=wu
�tV�>_g>+c����K�ݷþq�?�h�?h>�?��^?;��#п�⇿�������� J=��`<���=��0�!����b=I�!=/N��#�=2$�>ˏ6>�w;>H*(>:$e=9�=�o���j���E����8���C�a),��Hm�����܆�u��޾�Cľ�V��J��&������Ͱ�w��0o��1B�>�2?��>�>T�>+��> =��5nھ�%���{H�>d�)��������L�l:��t톾�훾1���d��o����>�۽�%�>��>	(��Cg��ip>�U:>���=E�y>���=��=Mh�=qX>F�>xA>_[>?q>�e�=0��%^�/~/��/����
C?��Q�l����2-���ƾ�!���K�>`�?�E>D*��|���hw�@�>|�"�Ud��_���佒�>�7�>�D>S�;��ƽ&t��
� X�=5�>HjM>N(���u���>��=X��>'�˾���=:��>�3?9�j?Hl$?�Y�<
��>a��=�|L>Ș;�O>z�r>�q�>�?~y#?3�3?pO?2��=�QL�0�;9�w=O,E�A��6�}�ǽ����f=0f��v��=t�=��l<R��=�8�=�67��&�<�
�=���>��?���>�"?�����41�[6�����rl�����t��:���>2��>?7?D�?��>�-�=|q��1����>���=�@_��7S���C�(j)��m�nB�?�a�?	�=���+=ZK7<y�U=ڻ?y�Z?�{?x�[��k�&������c��0#�7�Z����b��VA��򽻺;��o־�/y����������=D����E
��t
��1���>
&}={�-����=���=6D.=m��bZ�=�Q����=P�E���\� F6<�׽���:���=G�<��!>��(?�?̉�=^Ay>b%�D�D���ƾJ��>z�>!̶>Mh_?it�>��@���f� 	Q��,6�,_�>o<r?�G�>ݸǽ�`m>�8���:�_�?���>����>�:���y{�����>0T?G%�>JN�� T�����	.)�r�>>�	=��ɖ?�qY?�/����\�����F��
�)=HHս��N��ۦ��l�SZ1������{�l���=M	�>���?�F��w�W=F����y����Q��r1�=O��=���>ig>�-�:P��ߕ�����S;��޹:˪�>�M��|�-??�J�>���?�`?��A?bZھ7�t>P)>�t?�w�>��`>{#>�o�>�����RP�OpL��|-��ސ���==��<��6=���=���<�N�<3~�<���=3Y�;�Eټ��PM�<�e;��X��c�=�)6>u�>��?=@1?��O�V��>���z_>s�>��N>��ɽJ���� <��>GS(?��3?c��>��/��������u'�,��>�tK?@=?���>R1f=U�>k3� >�s���R=	��<!�`���q��А*��G>?�u>*&�>��>�ez?�O.?��>qW���~��N��V0��[=�|�>�J�>hDF>1��vD�Ãm�6�d��F*�����I�S\�=��w=���=�2>��Z>��!>B;�<�	���-��7b��d���l�>���>~V?��t>��=2߾�sA�ZcS?݃&�e(�,Hľ�'Ǿϭs�8�5�i�?B�8?��a?<��˄`�:T���3�[ؕ<���?A��?�4$?����:�=>½���aDk>����.��B>�yr��V$>\>��>�F���p%�G�>x�>T�����+�=� ,�;.�Կ�.�l6�r��ʚj��������3򇾂Į���[�-��x���G�ƾ�j��F�y�����Q,ξ��)�'���e?1�1?Y����%��������*���'�=�|�nAI��Iž�A��y%��Sù��ǫ���Ӿ���꾱�f���x>�羍M��p{h���پ�\��Wڞ���>f��,�S���!�|�:�6D>w}>W���7is�{ˈ�AVu�Rۄ?s�??�Q���엾j @�	h�m�e>�ٞ>�_>S����z��T~>{�6?�u\?b�9>٩h�
���V��=j�?[��?�aS?N�ƾ�dL�:j��2<�d7�>��>ܧb>�_�	ڛ��<��w5/?���?|Y?P��w�T�?$�,�?��?��d�_�!?�[�>,�>Ʋ���Ƹ��V>rz��a�|'Q�)�>�]i�����ގԽ���:���>G�|>�&����Ҭ>E��.�\��v��L7�h�W<���=h�%?��+�Y�>^�b>�۟>5�-��rp�Sy���2�K?'W�?2_?��c?����$��sǪ>C��>C9>����R���?�R�>����p�kB!��~?%��?���?�V?���>Gӿ����������=%�=��>>��޽�ɭ=x�K=tɘ��Y=�s�>|��>o>>;x>o�T>ś<>��.>p�����#��ʤ�3ْ��[B�� ���wg��{	��y�����ȴ���?�������;Г�v�G�X���T>�
g���?R�N?7{�>DNx>�s�>��>�����@ξ�R澋�������M���^���ѽ���N�� ��c0��a�G��	�oV�>K1=	pa>�Tu>��,�@>�>|�>�@>F�i>�!�>�	>`9<̼�=�4>�M'>��N>�&R>r}=,ł��w{���9��q���4<�>?a3n�
���,�N�ھ ���L'�>��?rF>1�'���h�z���>��e���\�Z�ŽS�����>���>b��=���;�7�4]{���ӽ���=��{>�>���݋��C���=ξ ?�\"�>�H��+[��mD?C�z?O2?)��%%?��>,�>��ν0\�>�*>f�=}?�C?�?�T�>�[�=P���3Ɵ=�N>\ڲ��| �z�v=��<�<3��޵=Ď�=\'L>���(��%v=�׼���`+�=���=+:?`?	n�>qE9?�� �JQ.�W�ٱ�=��>�tL�o<>8D�>�d�>��>ϑ?z�|>la�=�o�LѾL�>߫>�
\�R���i3>���h>E�{?�Mv?�����:��'��=�������>�_�>�F?���>�EN>*?���

��ɿJ���Q��&�ڥ��.�/�7�3�� S:��+�E���;M�V�C>���>YhM>>X>N��=t��=�>���=�{?=ԭ>R<Ӳ;�C����%=�����<&/>�?���89O�Sʺ�^����=(�xc���n(;�+?pq�>��>g��7S��066��D��Q?��>���>�`?{g�>�u��|�v~��N�����>#+�?�Y�>:�{���>�4��F}�=���=�^>S�8���#> ����2��>���>D�?1��>���:�{��˔��@����>��:=,��h?C�i?u
���i�M����E�"1��m�<��(q��ɥ�
����/��S�{WﾛEc�4o�=���>�W�?갑�,�>�	���H��/n��z����x=�W_=���>M�Y>��B�Si���;
�����������=�>�鲽���>�=?P4
? �}?)�+?^'?ծ����>�'I��3?3�>�5*?���>���>�ۙ=�J�<#�4��W�;�*½5���R��=�I<�9">ْ�=�˰=VY½�5/=��:>��>8ù=��y���@����<m�q=�c�<��I>�T>�q�>��/?w���:>����Ϻ%�
>ؓN��L�=9-��-�)����`>	v?5S?k>�>y���v�/{��l]�:��>� ?�?)V�>˔>Nw�=���2,]�p?��e�>=������Ⱦ�.��ȾV�6�6~>��=au� �>h;z?��?�}!?��'�ҟ��^����˾(՞�ݹ#�2��>��>�E�>�ñ�g�+�'V��0z���+�S�>�,P��">y��<*��=�Tl>n�(>�>Up=�ʣ<�{�$_Y�苶��8�>,�?�$?p��>{�?=]���l!��F?�X��[L�<���=�-j��Z=�k�=���=4�E?߳��ۢU�e���w���1m�>d�?��?��??esD�����'��w:>�xP=�ּ�ڎ����L���ݡ>V��=�?���Cо[�1>�m>@�>�Q�<nČ�os��%�#=.׿'�.����^�������;�B7�������J���;4�u��.k'�3I���1��ؚ�F)�������|b�?t%?I���s���1�%*�n��4�>�����պ��6�������ȽJ,G����z	⾀���
��� �=�'���zu��ˀ���8�7��ER>N`??��*�i�����n�=�%�=�t�=�k���Ǜ������D���?�{?�𾵑��.��\Ob=B�?S�>���>@���(\=�~>)D?���>�#=Q���qX���<L��?UJ�?��@?�ҽ`�9��$�����4�>p�?.y?%P9�;(��ї�G|?��R?�P�>�ھL	��*��>a�??ۗv�z�z>Z��>C=n>��b���T��=m<*�Z�=���=OD%����%���-��(>���>e��>*����	۾%��>Ė���P��Ɉ�?���V����wf?�Ҿ�V�>�U�>&�>�|�������Y����ǽ=�j?v��?�� ?pkH?qľ5<.��J��H��>=)�>�J�>閮�3凾\?�>#��>��~k������a?5��?y��?w a?��R�>Gӿ�� ������
��=%�=��>>��޽�ɭ=��K=�ɘ�%Z=�m�>���>o>C;x>v�T>Λ<>��.>r�����#��ʤ�4ْ��[B�� ���wg��{	��y�����ȴ���K�������=Г�y�G�]���T>���ʾ���>8:�>vZ�>+ i>��>f<9>�˟��v꾽O	�\		����".���-��G㤾���������%ƾ�[׾�U��<��"&?F:�=g��>��>�fT=0HZ���>\2>��&>��d>��>-?>N
�=RP8=��0>뛄>]�J>_%�>&K&>���b
����3������`��Z0?x��O껾��;�ǎ��u�@���>З�>��=6�*�aU��)��~��>�ߢ<8�����ɬ���s>�� ?O�>
�<���������&��.�=�d>��>�^A=���翽"�T�^�>A}�Y�i>�	#?z�m?~C?���;���>L'�>�{>f½�n>���><��>�?�i?dQ'?�?�k=�L��jP�=�fC>�i��6m��==�j�H��;]�m�:�l���=��>U�a='y'=_��������8X >�5?:�>fr#>x!�>]I��9�6���
�س�(w��<�K�=� �=Em�>�Ef?�/?s��>�=�uξ� ��s�>��h>8Ʉ��z��(>Aտ>�2>$@_?pƇ?�������H>'O��%�#>`��>g|N?wV>�)���u������ѿ��=.�Ճ�4Y���11��t�2Ol�zb�m.� C��f�=�xt>���>��k>�qB>��>�S�>��?�8�>1A�=��=��=�\E��r��o=�g���d:�����~�;|2P��oE�M�VH�dϭ�<�����#?s��>�h�<"�> 
���X@�J�*ǜ>���=�>�:a?Ic�>�fU�I�t�� \��%�� �?��O?���>Ч��q��>S����/�=�Wg>��R�7xU�ߋb���P��?<���>'{?��>�e:�`�g�4ٌ�yVI�!��>�I=$l	�oC�?�_?����~��!��]F�!���m=�C�cg���`(�rt4��E��� ���f�6��=���>�Ԡ?���ѫ=�=���ۛ�Y肿a籾Q�R=ڑ�=Rp�>K�M>��(�d�L��9о�1I��4g;ۏ>�Z���P6?�c�?�j8?l��?��?_�j?���?�kg�gzh>m�?r�>��F>
��=�.{���b���k�F>�&�d澪[ƽ��m;��=Ug�=�*=#R�;���Ӻ2>�Nc=߼= s��+��6<=EM�<��> R1>�]>�X?���>����p���]��q���=�1&>��=us6��1�궃���> ��>�{<?�$?�kD<�������[sJ�t�Q>@t#?��>��>��=>hv��ߙ��Yű�

M�IU>F'�2;v��?	�����i��<im�>�Ѵ>�"J>��>Re~?��>r��>�jA��������u"��<ghl���>R�>�K>�闾�S�O2��l�h��<L�O���"��n:[>L�n��F��:��=~Hp>�t�>�8<A���_-ȾD��)��;��>4�?�!?��K>���=r�ľ760�]?rN��>N�?D���v�K�0=~<����>�WC>W�A?ğ7���%�%w��x�-����>��?>�?4%U?8+a���@=���ސ^>�?�F�=�,���BC=�-t���&>OM�>E����a����=�˴>�U�>Tw����I���!н��ʿ.%A���ռs(���>��1�.��l���|�_I��'9�s����ӽr'�h"W���J�Z���R���/
��,�£?�,?�,h=JjR<�E����p���O>�͒�~=��Խ1�K ]�뉾ʖ��y� � ���0��>���x�o>�,�������2n�ڄ/������=��[?��ܾI[��;��k�b=t>E�.����\����8��M��CpP?Қb?�(߾�%�~����"�=,?�7�>T"�>Q+R�����2�>X�G?��2?S��E��S|��p=��?�3�?*�I?�վ�Q��HO�Z'��g�>�=?9�>)���HQ��Vn�K�!<kʆ?a�? ��b3��f.��l>Z�W?����H�>�B	?�{>���#���r>Ƈ��T=��~����ܻ��[�R�C���.�	gq=r4�>-;�>��t�y׾� ?
����z��8x�E'�_�	�s2>�T?�i=�4
,�����>�F,��[���[��m"�s�N?F��?"x�?ug"?�����n�XQ�>��ľ2
�
i�>:M�=�ac���?nX^?��,��k`�CI�#h�>w�?�E�?M[?Ѡ����ٿ���ٟξtL�����=y��=��=�<��~�<�X�=�6ν*���,��=�-�>�ł>���>��w>�>EZ�>L��[�$��.�����7� �8d��T���쾆߈�\��+�ھj)����;XY�=�鼟S�!0^�RY!=9n�pr>��>L��>� �>UjI>�*T>4H��+��u���蔾�y�\���Qt���_��A�m���;��g��ߖ�n9̽ې��,�?nb�=��=.��>�=���=��>ɛ�=QT�=_VK>h��=X>�>�(e>�>�	>V��>���=jMi>��=:~�yZ��+�4������p%�ʓA?6���\��78���K�۾�NG>2�>�55>��-�S��8�x�8[�>$ŝ<�{2�:�6��F]�Uȗ>�s�>���=Ȱ�� (<�L]�IY��T?>-�Q>��=V��oI��f�$��>���> ���P> ��>�B"?U�o?��2?��u��>?�j? �=�2"�ZȆ>裨>�?Ϊ'?>w?>�>?�j�>s͚=%9[�$�=��+�v�۽'ڽ�����殾U��M�=.gG>��A>:��=!w)>��=.!>�־<��}=}�=a�>��6?AU�>W1�>���#G��"K���4=����龷	?��>$��>���>ZS�>�W�=�PX9�ʀ7� }�>�`>��b�.h�����=0��>�X�>Y�B?>�����#/��>>�� >s��>@�E?�T�>����\L��ۈ
�վܿ��.�x5��n�mE*�(���s�7���z;Q�%<!Z(����<C�>�Ŝ>Ϩ�>V��>�3�>��6>ٹ ?@|'>�f?��b,=q��=9�ѽϮ|�=&M>c��Ϗս�\=Lq�=���<L�U��Ԁ�>>�������x�������?G$?�!��iE����w�XT!�/?�b="ނ>��?Lc�<֧)�Lz�Z�t�>W����?\i?��
?��ؾ)�b>�&>�R�=�K?w<?�C,>'j���5>2C�*!���>/�??�<�=�i(�����:*���>�>gI�g|�?�va?�?2�� ﾰ)�����\%��>NV$=B�ٽV���D� g���#�!,Ѿ�S��/�<ȇ�>Eպ?󫽼n�y>�l���뢿0/��[�A���(=B�8����>Qm�>�	��ɾ�1���/M��v�νk$>۝�>�`�>��??1�?#WO?�3\?��V?�ߞ=S�u?uZ�>�G>Y>�?b�?�.?uO?jQ>��=Ag��z�X�q�.�5�u��<�h>�a>^3>OK�=������$���Ƽ��=�铽��w�	�;�ZU=��=�b>��??C?���=r7�_S>F
������_��={�C�ǈ��w�=�w�@Gf>�.E>� ?H�?	��=1��GF�����|>�?��?�_?�2>��p>�<���,>PT�>���=�,��(Ӿ'9��ߕ.��|���>k��>�>��>��s?�I^?�Y?�ZD�;Ą��%����m�|�*�.�ܾ��? T�>V�(>��e��!���R��Á�/1��Jо��0��{S�^�	<�=���=�,>;�Y>���=��께4��tG=� ߽r/>($�>Ɔ^?�v�>��>�:�ľ�Ͼ[�I?\6�����䟾�Mо;�$��>��@>z�N�? 
��N}�b����=�Q��>��?f�?Yd?aD��t��?Y>��[>W>���;��C�NX�XT�� �1>A>�=��x��ו�9&:;�7\>x�x>"ȽZ�˾@��V�B���ff��Ǿ����L���� ���ھ���=��������6�����к+�(�N����?3�O�J��'̾�䜾V��?i܋?��>�K_����8:(�#:�L?>��9N)����Μ���"�%������F���A��E��
���>.�z<�'����C��K<����(�>?��0�����_����օ=	+�*8�<N���bYÿ�AǾi�?,|Q?z����C��ா���"�:?^��>��\>���;������a?��_?��󑆿�܍�y�����?9��?4@%?DD��&`=�!6�^#�=Mf?�?���>��]���t��q#-?�F6?�X<>I�`T|������>4�W?�`t����=��?��>x�����w�M=����=5�9>2wC=��m���F������d*>Y��>r4�><�|�pn��F?m~�� |��Z�j�l/�O6ڽ�z>ά?s��+�S>�=��^>���n��|�����Ӿ�z1?�ù?��?7t5?s���ؾ�u:�F����>��?���=����|c�>�?�@��B&=��{�����>�K�?=�@�At?Z@��7�׿�5���J��s���L�=i&>
��=�~J�M3=��<�W <E����Z>��>f`r>���>�>6�G>��'>Y��?~ �\$���2��['D����&�=|����s��[��{�׾q;˾�K<�u����e�=4A2��r�A\�B�d���N>N��>U��>�}�>���>� n>���˾�'K�߶���mӾ��ƾ����]vþ������ڽB\���4�Zq�jeK���2?a4F=�t̼�/�> w2���9>&G>w�=չ%=�`�>�e�=���>�>x��>:�^>�O >X�=���>��>�um���j���4��$L�3�:>j�2?�d�����K<T��#��Y�ǿ=n�?��>���ʝ�G���eU�>��0�:�O����<�+H>\2�>Y��>��=�B�9������M|��M3�>&jq>�Z��H��B��5B=��>�4־�:E>��0>wO?~Zi?l=	?K�">��>���>�^>�s�>2ڕ>�Cr>¶�>;� ?�2?h�,?���>Á)>쪹���`>��3=�������]�WO｡J���WS���μ�I>��l>�R>�1�;J1=g`@�wiD����=Ճ?Y�=?�>E�?���lL��>�|���
��f>~��>���=5Q�>��>M��>c�H>�?>K��G�.���>T�>}�/���l�>���1�?�2?�lN?W?�?t��X�!�[�>�c>�C�>y?�< ?���8F�A����ٿF98�'�~��_9�ʐZ���;�H>�U� �M��`��V݌� ��=�O�>b��>TY�>篑>RK�>ۨ>H�>�
>1������=&{�=~c�J�h�v�=��m<ܯ���a�j\�<�d ����Ʊ.�Vc��@��9
�=���<�D?ؒ?��B�-�2��^������$�>�z�>��>���>��=j��2�D��OY�v�����>��q?�?���'�K>6�<�μ�J?�v�>J�=�]E<�$ϽP��q�����>��?�}5<zX����'�pZ~�al0�邛>�!4>&?�T��?��w?�*������?��D�Y�V�>��>zz<sB��~���l&�����������-i =�>_�?�
���)�>o��X�������9<��9L���H>��?R���ɜ�j�ݾ�@�~�������<w]0<��\>�>��C? ��>�g?n?e͎=�
���e? i�>��>�P�>X� ?�m�><;?lT?W�=�1j���3��o����s������L)�6�=������p��� > >�0W=�3)O;��;b<༨0�;�e�=��A>��
?�$0?�>Bzq>��>����� =���>���>�3U�- 	�w"��NN>F�>�K?�? �>1�%��_)��kྫ�O=e;?=�-?M?Q��=� ���Ʒ�Z�,>=M'>F�r>�G�=���=�̙�D50�H��<��.��>농>FX�>)�w?�@?1G?�����N�3����,h���A���@=_k�>p��>C��=鞾ݧ>��gU�u�P��g$��n8�#3��	'>h옽���<F��>�%^=�>=�U��I < w�;Սu<f�P�%�>�"�>9;?z��>�>-����#�~�G?{�G�������	о�	�=� �>�!w>$U� g�>�����?��T��q	G����>�k�?��?�!?�[���	�+E>{�>s>|K�=}Ŏ�/����,>�~�>��	��2��?�8�9َ<��>���>�g��k➾0�оu�V�m��o�ת���s�� ���%�<�f
f��ѽ�﷾�@��ƨ��J۫����}�x�1>��yТ�l9�0� ��+����?��x?+�>ͬ�>�"ھ��%�Y����f<Zr
�r���:�ʒ���M���&(�mDR��0��k>��J�?�>�����kO�I�$���̾2G>}�*?.���w���S!���	�$�������8�'~��)�ſ1(��o��?8f_?J�\��P�G�ھ��
=?�ٷ>\}�>e�.���z���˼>�W?��m?��=4y�� ��Z4�<�V�?���?�;3?�"�=0�w�';�ⅾ��?�zk?�'?���UK ��B�=-T�>~�
?�h�+�R��I���Ͼ�=?cg?����z>��2?J��>��H> �F������@�>��>��=�M������g���{>���>!3�=~���p��/�?�6������3`�"/.�
ղ=�;:>�R?��2�)�d<V��>e��>�q�3Ԓ��ˋ�v���u?�?�$�?�B'?��4�O�$�8�D�葾�!?�B�>�f�<³����?Q��>��=U�7�[�,=4��>$��?��?�{W?��X���ؿI��������B��U>T�л��>&  ���=�|�As޽�'����=��>T��>f�|>�M�=^��=_/�>m��+�#����b����?��6$��a����C2辁�����:U㾣;���r�e�7�@�_���?���V�J�Iϧ�л�=B��>&�>`��>�^�=���=�u����a��ӃH�������Ϫ��~���􌾲Ǌ��6���e��G��<��ᾁ��>M�H=Nk�='.f>4j�;��=?�?>�y=�tr>�v�=���=�+w>Za
>B>�=:O9>�;>ü=���>�=I>��i�*,t�sc �8M,�t9�;?��s������RU�#q��%kھ�Ԁ>��?��I>�$�u���a��UJ�><��E!��?�ce��9>7��>���>;�=��k���L%�DEZ>���>���>aŷ��fZ�z�B��yS=.�>��g�7>�`r���0?�n?j ?��>�?�??��">���{k?���>�s?��W?��2?c�?�P?�w�=�k�_�J������?��kJ!����H㽤H$=���=�_d>@<b>�2=�<�=�=�����-ދ���<�a�>j�9?*�>�:�>��8�t �e�Z�U#���g�=n���£�>�ռ>"�>Ҿ�>*O�>��A>XQ��<��2)��T�>D�]>�_E��e����=?�>�W>sQ:?�?�bd�줼��O���=��=}��>�?���>�*�<���E7�&/ſG���3K�W�i齾]P���R����;�A>x��7O�gl-����=��l>W�h>S�:>��1>O->/��>��?>�^�2�N=Z��=H�j=%􇼆��<�-�n3�=MV�=m�=8谾(��������u�κ�H��6�F?>m*?sE��.~���þu�	�(�=8�?Q�=�Ո>@?��>�Ͼ�b����e��j����?|?�w?��ӾvI�>"Uy>�O��n-?S�Z>���<2e�D�)=t��^�y�D>腼>GO
��$.�̬U��,����8�;��>_3S>�،���?�?l�W�7@���E�5�O���D%սY~?=�
=�.��Z&��6R���VS$�3z�d������>���?�ᇾ�k�>�f�/���=�����\"C�Jf�Co?���<ؖ�sV���	-���Ͼ9!۾��V���3�<5U>�`�>��8?���>!`X?��@?@?��= �H?���>�>z�$>JQ?��?o+;?2?�>R���I����ν��+�?������s��=�#�<��-���H�>�U>@�=i�X��7j:`B�=���l��=�U�=@]>���<�?�`A?�H>\�>�'M>����,>��>[�?D"F�nF0�����ky>��	?�X^?���>] �9�B�?N$����z�_=�%?�T?��?���=X�`>���<��B>����@>kӁ���߽����4�(��=���>��>���>��>�o?�?QN=?N����C �͝��VL��F戾�7���h�>W�>�z������)<���W�abt�J�:�ȾD��G >���~I�+5M>��1>!��>�P�=�}�	���N�,�$��)�>��>��:?�m�>�U|>٤��`	�^J?&����������wѾj�!��J>��>>%���?W<	��}�����n0=��H�>#�?���?��d?�B��Y���]>6X>��>o:<ĝ@����ć�R4>�6�=��y�����~N�;
SZ>%xx>��ɽ��˾��,�I�7"��zN�(���\��K�	�@"�Q����ν�y��9������d�7��zb!��!���v�`�s�OoE���X�Xf�?^�U?6,>-�K=��<��H�Ҿ�Q=B�1�<,����ܾr�V��?ڽ����a��7�)�����u���ܾ��>*,���5
e�����ʍ�=��?��Ҿ�g���"�`$��!a=��O���;��1��(����b��,]?�WW?�猾�'E���I��e��g8?GN�>���>$#׾�_�>��4?�H?��<G���m��,>���?R]�?w�3?#>w<_c�ڍ���=
�>�f3?��-?�P־����AF":�.�>j�?�����!�h����վ��$?�т?����f< >�|?���>�^��ľ���H��9����>D��>�O`=PK	�.jd�/��\�d>#.?/^ >�cw�k�m�t�>&���Yb� w�}N2���P��!�<��n?_w�ľ�> �>U��>��}����u����}���Ŋ?i��?�{?�x<?X�R�?	�������?�;[U�>��=n�1>�H�����>��?�?ɽ�P�������>�~�?��?��E? �,��ۿ-��%O�����V��=���=Q�S�1lz�-_�=^�=�|1���۽��=�w�=�!>�ߊ>tF�=ǚ=�\>&��`���ߖ�XϞ��D�M�V��5o��t��;���B|�=���>徎a�PI:��n�6�z��yx����@/�Z��>�7?i�?�:h>��>/��>~�K���o�!ԝ����8�%�Qa����վ
�x�6�_�2սi:���6����,���?�򄽙y�>5()?駊��F>�x?@:>��(=�>>�=��^>�J{> �>ܿ>��p>PZ>K�{>�ʐ=���� �}���7��]�p�;�>?k]������3�J�վU���o��> q?#�J>�&����x8y�vl�>�&�>�\�f�ڽ��C�>xz�>��=��X�m�޼tW��� �ċ�=��>J�>�D�拾�(�苾=��?�ҽ���5�03�:�O2?��?j#U?��=?�"?%J�>�/�����毯>9�E>7�"?
T?�?��?8_�>cuQ=,��;��eI/���̽<=���!�<JA�bh�=n�>=w<�S�=x�"�����_�X=�,����>}H7>�?m)?�U�>p�I?PpG��N�
�6��Z���Q��r���O?;c(?Oi�>��?)@�>|:=��:�gH'���B� �>�-'>4�6�Xp�"/�	H�>�
?(0?�G3?���9�Ӿq�|>ְ(�?��<S�?�2�>�ش>Q��=������
�.,ۿ$X�W����>`ۼqß��қ�f�ͽ*B���-#��3�<X=�u�>�r�=���=���=��5>�A��<�>�f=�vH��4>� ���+�,�X=�>����z����O<��<jD]��5>^�=R/
����#I�=O��=| ?=�>����w�u�x־B�gG�{oM?�8��B*?!;?�A���J��
����o�A%��i??�߆?WC ?|�;�_t>W�>1��>�K�>��=78>Ύ��u�>�_���"�mн=�1?�a�z��=T�"�і��}O%�Z�>�K�=�I[��^�?��m?.�9�E�$���:��,�O��u5>姽�F��[^����,�sԭ��%�����r��=�]�>L�?���1?�s&��ç�o�>�'�o�͸���۳=��>
����)>��4<�T�`���G���;���-9�w�H>��?*(?���>� e?O@?�� ?���.�Y?@��>�O�>��>��Y?̜?�[.?���>厮�.[�퇼N�Ͻ�m����-����h�<�2&�����<}m	��w>���=�+�=\�O=��R>��>��;�TH��.F=
u�=�?BS.??Y(��]=�S >�����=�>v��=Iո>�-���|ɾ2��I&�>��>��J?��>	w������ؾ7ӾPl�=�?�?�)?�x>Lد>��5�ӿ&=��	>J|�s̭�����`����P�����V�>$+�>�|�=8�g>Cd?��,?K�I?��ʾ/*���p�y�����u1���6?��>�\>��Y���K���3��#n��u1��E�� �<��Kf=�@Q=un�>Ұ[>����/i=�>iH�,Eӽ��4>��=��>��>K|9?��S>,�B>#�侏?�C6H?����?��˱��3޾��G�
>���>2)�� ?�Խ^=i�������?�׶�>ʤ�?Xs�?�cj?�����ݽe >�>�O>�2���4���j��緽�3'>QR�=Zm�𹔾5��<�a> p>��ؽ��پ��k7b��-���jK��5�+�ؾ&�A���Y�|����轧ľ�뀾����L_��l����F����-��;�������ƾ>�?���?��>�'-��5:��.����ž6�<�I���T���X	���+��2������P�Tp ���&�=��h�>�`�Bz��U����F�Ǭ��o�g=ԃ&?(�Ѿ����4S�"NA=��f�O�-�cc:��眿�ꉿ�3齞�Z?qnO?Ĥ����!�$w���K?���>ΰ�>�K�� �]�R��>�68?i��>� ۼzN��4��L��=�T�?b��?U5>?kx8��&A�Pi
�3���?�A?q�>�'�����3�����?��7?�)�>V�����d+�K`�>�x\?�SU��`>%,�>+��>��ڽ���N�������$��O&>XkL�$����O���.�mq�=��>}|>��K����ˆ�>�l˾�Ԑ���U���e���6���_=S?��#�Z�c���>���=ߝ
��v�_���;����n2?q�?��z?�x?�y��ӛ��Ƴ��!�n���P>���>��>�rk��?�
?����"�/�2S��32�>k�?�c@�"?������ܿK��� ���&�̾�g�='Ͼ=�>�a�����=�ޝ��^�yH�>?�>R �>W�x>�R�>��d>/">��C>�;����#���������4�gD��-�^�� �r�t�5����� ���Vv�;��6T����a����pꬽ��eF>d$@>��w>��>Ҁ>b�2>X-�������2��B�=��70�y�(�Q$�!�U�]B��(>��L+��ܼ�нc�0��,?��~<G�>֗&?��4���>G��>	c�>,I>ׅ>�J>���>BC&?<�.?�o�E�>;���ڄ>�,;�H����~� a-�)Е�u�<z�*?݄���ǳ�
���w�T�о|>R>��>EK�=��0��;���}���>�����E@�cu�?<��m>�ı>��=� %;�Y�j(U���5@[���N>�^>�F&������F����=
��>'j?=� U>ă��To7?�a\?�(?���>� ?��*>겼=�kq>��&?
��>�?�8H?��h?�U?c�>3�>Y����2Z�# 6��Yk������y�kc<`�{<�x�=�|D<)��=��>H�>�0ܼ��c;녶��1�=�D�=�r�>[F?m?ρ?٭c�}�ݾm;2�J���y�!>WQ���tx>��>k�?؟?~�>K�=�3�<���i4�EӔ>�)R=[:�7�w�KH�<�z�>�|�>Z}5?�Z?
������u�A=X#���{�>�"?��?SA�>dH=C���������,�0��E8�%�ֽ��
��\𼧡��!�/�����"�}�<&k=�0�>C�>��P>o>f�->М�=���> ��>[?��{½�t��W=� Q=T��=]����=`���M�{��T.�=}I=E����BS��)����=�������>s?�L�~@^�]���&����#��>�(>���>I[?g`�= �bq�Uo� ����;%?X-Y?��?�ƞ��p�>t=�c���<?S��>�	��N�L�i�>����]㐾b�>R�>&%�M�*d�'d���3P���>e�.>{���ҍ?�;v?+��Y�p�;��o��l�9*v>�������鵾�����U4��K���� �r*����?��? \���u�>�N���q��Y%���!�G���=��4?��6>*PD�Rᾪd�b����ƾ9���l>A��>N��>�]�>�@�>�q?K2?�?ݓ�>rMW?Baj>T�v>i"�>o+?3g�>�ME?�^$?}��>�>��)=�Oh�طs�E&�=	7V�g��=d��=
g�>���<����Ae�������ζ�|^Ὀ����Ie�$�̼6$5>��>��A>DM?2�?`����<)�'>:��=ql=�	V>Ǚ>VZ���3���X9�s&v>In�>�+C?e�?���=N��ƾ���8��=�o?�L*?Ev�>��=]�>t_žG
���4�=��>Ii�<֬�G�ƾ�����[��>'�>g�����>4�x?h%??�K?�{׾n�S�Ll���������=_d?1�>�
0�u����*�Q+e���Z�v m��澾6����<��uF%>X7�>���>�)�>D�=S`<����U]5�km���R->*A�=^'?M��=��5>�����C��D�D?�2�����������0����?>q_V>�+�H?į���y�Ƴ��A�7����>8F�?!��?��h?��7����u�o>s>ؽ	>�F<=�=h��x�[Ӑ�<�=>��>��g��
�����6>��t>���s�ž���1�
�־�M���!���xQ)��ˢ�P���սrG<��"����E�L~�z�{,���v������/�|�v������?AB?wo>~��>��#Q%�4����#��7���Q��X�����ˏ��ǖ
�xU��!�g41�kG���=E�p��	��BT�^�$��Ǿ��:>�\?����'������-�c���w��4-�n������ tm��
�?1�U?F�8��?��-������-?��[>��>ʓȽ�/���W=y�D?ח]?ϭ�=n�����n�)�Pd�?�t�?:�=?:�J��bB�������[?�T?��>԰��f�̾����mz?�
7?� �>���c8��1��6��>��[?4�R��b>��>PO�>h�ҽ��� �!��^����׻�W>>� 8�4J�\�j�v=���=w١>?-u>c>e�������>J���L�H�z0��`�^[���	�?h���Z=�њ>U�=5�ㄿ/����s���5?Y��?�Q??a7�中������=H
�>f�9>/ұ<Y�B���>"W�>�vξ�j��!׾�E<?K��?�W�?Ed:?��f��9ؿ�e���W޾q�ݾbX�=|�K>A�3>��K�>T>^s��&
`�z�¼��T>��>@��>:!>mz>�0V>S:��'��Ϧ����Λ1����7���7�,�%���ǾW4��dپ����\h�s����A��R3y��u�vډ�������=>��>:y�>���>�0>c:=AH2��'ξ$�<�����l2	�Q^��)�ԾWؔ�0w�y�J��2�7�!�B���$�9,?�����LN>k�?w!��#��=�V|>%�J>Xա=X
�>M�(��ȓ>u�>(�X>��M>�W1>@=��n>sc>�P���������;������?�[�6�y�_Pd���M�U�����>R �>^��=n�2�����~�i4?�BD>���E�|䊾Ww�>S�>v
�>�	C�����h:�o���ȭ�=nt>gL�=���ڄ��#l�>�2?R|���&p>���>��>��=?��?��k>�?�Y�>B��> �G�vxf>/�=L��>�o?�	*?��F?<�/>���=���.>M��ZM+�7�X=�a�=���=��5�s�}l��/[b=�()�Y�D>b��=�%;n�M�F.���(<0�>�L=?�X�>�/?�S��5�TU�qȶ��c>�L%����>~�|>A�*?�؏>��>P�?>���=�������>�1>Ve����.�s��A6 >-�?�Y?�r2?��A�����s���K�=�v�=Z��>IRW?6b�>��n>[cC<i����ϿG��A@$�L��x�=8�=W˽rͺޛ�3�Z��U��0^���	���>jҰ>�.�><�>b�7>�a�>`p>���=��==�R"<���Faؽ�Б=ϐ���n=��R�>���;�l����n�y�{�e=作�<��?��?.�4�Ї�wS����2��z��>�w�>��>2u�>�=�վ�Z��<P����0��>�kl?���>�k���=��e�vq]���>��>[��=ۗI�y���[���ۋL=��>:$?[��>���"dJ��oC�V�����>t|]=����ə?�T?��;�͜�f�6��X��p�ԥ��Qv��J+J�+�ӾV�޾~���j�m���R�����NM�>���?����=3���
ᒿ"א�(�nی:��H��>��=��n�QbA��+����b�F���Q>� >Ώ�>�w*?a�9?�t&?�*?N��>�va���>���-	?�W4>|�>��H>�;�>��>V%�>�ds>5���(����.���<��=��=��+>��>.�=�I�=��t=}�'<<{��l|��δ=�2��z1=@�,>��=���=i?%'�>����O�=�o�����ҚS>�X>��>S����/�_�.��J�>��>�S?.1?fp >�1{����uо�]�2d?�?�/�>�'>P =_�޾�B��6>�G>�x�<PC̾xq$����>�s��0>�ȭ>'>�E>ւn?I�^?'?[U#��1����S�������8�>�:�>�˔>�]�1,��I{��9���2�ڏQ��?E�ƈ�=�%=S�>=-Y>-���"��=�B6���=̓r���@>侇= r?�^>z�?��>J�4>�\���Nؾ��J?�H��Sl�&���a�ξ>K/���!>��@>�A׽�?(��dL��j��aZ<����>�k�?���?W�a?'�S�B=��NAZ>F>;�>6�٦C�R�⼶S?�(s:>2�=�:s�9虾�'e<�\k>��w>u��� �ɾ�z׾*�<��ƣ��j�?p缣-8�%�>�����
��S=�NS���ׯ>T�P�7y�>=����<�PƽR���AC�	��k�=�e<�?x�^?�j<�����Ǿ٩۾!�Ծ��t��=����Q�= uZ��r�;�&Ѿ�|	��[@��P�����^�>5�=�����!Rh�qʹ=���>�9G?9r�����͜*��'�=F�ͽ�#5>�t!�4���$����x���W�?��&?@��\���sl�>e@�+�z>>F?���>��&�jx�>��?DX?q=�ڨ���ꖿ�萾*�?��?�R/?��=m�K�y(ƾ�[��D�~=��?�?����������>�/?/*�>K_�{	��xO���?�2�?����'>��?�f�>�}!�lBѾ̆���J��G�=�/7>��6>6��s�v;�{��~�=�"�>Z�?�-�h@���>���;�D�Ϫ?�r���˖�nF<��?�y��>�>p>(E/��j��\G��N�i���'?!5�?�h?��?��ok��)�;�$*>&u�>�X>�U��jA<F�;>�a�>/mӾP�@�������>,v�?"�?#�H?�|���տEr��Z�W�*������;o��<o>�o���=i�V=�I�<�ս��<z� >ܤ>9�>>��.>��$>X�A>M݅�	a����Έ��s +�v� �����`����ΰ��&�:�R�׾^ؽ��ԍ��q叾�Y��a�V<��Q��OG="�>���>��u>��>E�f>�����������i�]���%���Ǿ��ƾ_gǾ�tb��������=ƚX�4�#?K����e>ڜ?j���葽6�>,H=�`�=��>���\f�>� �>(A>�Y>h�ռ��N=�2>W����x�n뢿	�ݾ�0���E� �>�«�ͼ�=�2��#�'�Ԗ���
?���>�->�b��k���s�B�?t� >�d�eCt�)�q�W(;<1�>�R>�����';������=�˫<�B[>̋Z�W�=������.H�+�?��x�
�=Q��>�-?U ?W<9?�;�>m�C?��>M?�:���=�>Ă�L)�>,�E?�n?yH�?QA�>��c<�L��~B=���`�#��k+��+�ݞ��9J���P�=���=��L=	D=å�&�)>��>���<�9>��=��>έ*?�?}�?��7�E��o�N��"����>kM�;��>AN?�D?��>~�>b|�>���R�;PI��ĕ>A�=�'[��A?�f�= ��>ET?�*{?@�
?�zu�&z���d�G��=��#>��>��)?�g�>&D>�Gn=̶ �S�ǿ��K����+q�=�N¼d�/��<��M�߽��Ͼ,�����f.r���=��>r�t>��g>:�=D��=��>x�&>��=T�U����;H(m>z{�<e|������4�=�TV�`=�&��Tw �jr������= 9�= �>��?rB?mT�����O�}�ƅ�L���4��>�U�>�C�>���>1I�=�M�y�X�=NK���m�3��>�`?�>?ntZ�m��=xf�����<HN�>0�>c�>E����w���#ĻJG�>�z#?���>=��~wS�i�X��9���>��=o���J�?
E?M� �<���C���Q������D����J���E���`�5�)� 5��
������0=�>�X�?�]�uV
>�2��������������	[��>/��>�A>�>$����1�1�ʾ�ʞ�������0>�#�>L�>�R?��3?��"?4^?FA-?�:�=��>1gW=�o?2g�=�&)?���>�-�>� �>�>PGp>Ɋ������O�hݽ�q=X�>X:=���=��=���=k.�6]��h��z%V��C=�k����ٽ�h >���=�8�=��
?h?�sŽѾN�����`�Zm�<���=�;>�-��]�Gv�<߸d>+�?�*?<j�>�b�=��վ�Q��-��>�=��?Y�'?���>��<���=����{��l�=1�M>��������
��~J���>��f�>�~�>���=�A�>��?�H?j�?@�����B����cI��� �f涾y��>"$�>���>�-��[/v�����	M�oE-�_	��+��M}��]I�=
0�>L4U>��^>��=����9#�>}i�]q�<��>J+?G�>�$?�g?��>`�:,���I?2����Y�,q����Ͼ ��S>�=>ſ�ٶ?N�8�}�b奿C�=����>�w�?p��?�bd?��C�@ ���\>MpV>��>)�4<_�=��?�����3>���=��y�Q����ئ;�^[>z�w>�ʽ�˾� ��G�Oi����U�K��M:7�/7O�N{۾m���*��Ԛ���Tr>��G��X�<ŀپ�>n������i�P�ؾ	�׾܂?��Z?󈘾����F�ݶǾ���6>���O�S�������x�;��p���&ھ���'�D�2I#���?�Ȋ>T��~���Y��bg��-
�>o�p?�@J�N����;��<:��پ��=`�*��P����ſ�{þ8>�?�M?,趾[>����?qso=��,���>KL�>\��x����_?�@�>~�?�[K��Q��젿hl��*�?��?=�??tjI�B�@�a��r�m� ?��
?D,�>&%��"wʾ�'��
?_6?�`�>���υ����cb�>��\?��Q�l�b>^#�>ˌ�>�޽�ۓ�BQ�(4���3��4>	s�( �Uc]�D����=8�>x�>Q^]��f�����>19� �N���H����{���U�<�?h��$>i>A>�(�����ω��:��L?w��?_�S?�g8?�_��u��4���;��=���>4ά>���=����>1��>i^�}qr�W���?�H�?+��?(ZZ?N�m��_ܿ�A��ߠ���8����,>��'>ϝ=F������!)�(x:�_��9�9<~�=<s>�m�>T� >�Ӌ> yb>�f��#��|��
u�����Πپ!]�x���d�-��1�0 ��l�l���'|c=`�����Ͼ�\�@����|�d�d>���>�d�>[�>�p�=�E>��K�uپڲ��� ���;���ˈ��ؾ�*¾�þ���~N�����"�u�,���?ڈ2�f�P�t�?��=�|�<��>�ܳ>6Px=���>6�+=��q>�I�>hr>��&>�9#>kG�=~�c>Hp�=x܄�~w����/���0�M�E�C/?�>��)��	�M�*�
ľ�ȁ>��>�b>�-�jᘿl	~�W�>m*]=g(��<��9���nV�>��>	��=r3��E!B���;��E�<\�=��>
�/=����z���X�~�aR)>R�?���Ý�>J]%?6>�0f?P�?�l�#�<?3�>N[?Dn
>�L>�Ș��3�>�	/?��d?�E?mu�>�k=�D�R�Ǽ�~�=w�o�S��_a������{�����f;=_�= ;��^t=���W�> �=�B5��M�=`"�>�)L?�q?',�>��Ǿ��Y�U�������!�7>��\���>�W�>\B?�\A?\�>Ʒ >Ȍ�<	r���3�Ә�>��=��=�]�-�����rB>�>ׯY?b�g?����J����H>���>��=�?A?���>�?�V�=�)��2���}���H0�y�>)�߽�o>���=06�bM�>����W����	��I.>�m>�"i>{�S>o�>Q�����>��Q>5/�>�������<I�
"P�բ]:�!���Vɼ� `���A>��<�b�=�U��|d��t��Žr@�=�?߅?.$�FP��@g��6��蘪����>c��>���>�G�>�^�="T�q.U�/HA���H�g��>��g?5F�>��9�N��=�w(�қ�:j��>R��>'>�d��~�[7���h�<'��>G'?���>����'Z��n���	��>)��=Mս��?��P?��"C��� )��+-�q_��<3��������쓾��b#��O����J���g�.=���>(�?�ǆ���A>B¾+��n���G��\��<�D����>��¼�/Q��ǿ��S�9����M��e ��E>�e|>��>!?z�0?�2?qu?dt?�Aɾ۷
?���>��?$C>sG?U�<v ?p!�>���>�@�>�,�ip��c���	�<H��T>ӪY>�>���=.�%=���=��An��c�1Ԇ<)B���qý_�=�K>�a�=��>��*?e�=�I�=���l��<1��=5��>�-����нpye���>��>�w4?~��>)�=d���,(���ƾuº=���>iH-?�n?A!>O�=e	߾�8��OyE>�E_>�dA�4پ���󤾁�3��� >a8&>2��=[�]>D��?i(?�X?=�X���<�W�������R���@k���>��=@D�>��q�pE-�6�m�>L��~[��=�%䅾-7�=/)>���=0ۯ>�n�=�"����I���=/�b=w�s>�;�x?�%�>ĥ?}�>��>�i:�!���I?�k��Ȉ��E����Ѿ!)�4�>(�8>v��9?�,�|�������<����>�f�?���?�cd?�B���+]>RU>��>��X<�?��6�-х�W0>��=o�v�[��jOn;;�]>��x>s�ǽ�ʾ�B�>I�h#���QI�9���B����>�h��Ofƾ�Y�a��*j>-lZ���=�2	��	�>ſ<������?Ǿ�g�����z�?���?�퍾E�������P�>O���_�=��#��n��`9�O�����{�gr������t~�A��W �7��>��n>mb��ܓ���I^�#->|O�>I�6?���6�8��	6��ꚾL韾�l`��b�S!������^ ��|?�&?B����=���>���`�p>s�?��>5��Z����?��?� ?s�1=$gg�z���1�mM�?���?ŷ7?(l��u$����M������=�?�E?���zb����	|?	��>��>�9����,�H���}>��}?�z���.>C,?�'
?I��"�P����^���쑽�3>m�=I�)=N�N�2�=�<ހ�>u��>�������ko�> (��H�5@�3 ���&�_�"<���>� �����=�J�>��0>gn"�W����މ����G?��?zL?w�4?xc��
��Q��{��=���>���>U>���M��>���>?3�V9u����?4Q�?�g�?++]?�~j����b����������9YA>��:�<>�	ݼ��=�۬=�ws�檣=���=�2�>�6>�+�>�MO>α->�/$>���K�"��$��Ǡ��P2��eH�:D��A��s��WR��K3�픤��s��T��:���ӽe�Ѿk�������/Z��K>V�?̋�=���=vGڽ���<��\�,%������i��K꾐��ܰ��_���谾M��_���?�7"�ň7�S?[_>���=�;!?�d-�{��=�J�>�>>RZ<D�+=]�;>o�>�>0'>��>8\�>�r�=��</��>��w�L����8g�y��
���e?b��F��3�l��aԾe�ƺ�>Xf>�6��$�S��ٯ�C}����>��=�if���O�<^,��i�>ܚ�>�9V>��<|N�������;L��m�<}v>�8>b%j=G���d�i>b;?�d������2x ?���>b~U?�V!?�'�>'B#?��>>2c>gvξ}�>�����>T�.?�xP?�,9?ԩJ?�z>y���h%���(�J�����XW=���=���=�y=�&���?����=ɶ<u\�=yS�=X��4��<
�<*��>��?���>���>�ѽ1�7<g�h��C�L��K�I�?��*?��'?�?���>?��=� �,ľ���ܰ�>�K>ݺm��>6�f^�=*y�>K^?��y?���>(WK�PkG�iiȼe���6^���>ZE?T�>�;�>D�Y;ľ�|?ӿT�#�@�!�Um��§����;�<��RS��䢹��-����ʮ�<"�\>e��>!�q>~�D>S�>�x1>"A�>�(G>Q2�=P��=#��;���:G�H��NG=�����Y<��O��S��VEż�̖�P��J�jB�-*��~ܼ��?��?]��������V��C��~���m�>أ�>-��>i� ?�>U��snU���B�� N�v?Rh?6�?*46�1G�='s��L�	���>+�>.��=������B���F��=5
�>�c?@"�>4�*��G���[��O�`�>��� ����?�OH?mV���E��2�g�DY�%���*�:�Ž5�Q-���+��8�	B��$� �S�g��s�K��>��?���#_d>1��������i���D#�]0+=�Q�=<�,?7ݹ>�\�=�D��|Z�e�(��P۽��a>�=�p ?�g?L��>]P?��?�V�>��~��ү>���=w?k�>�v�>��ڼ?��>��>��>°>�?F�'k���j��m|Q=�æ��7>vK>t�->4��;�u<�<�=�d�<'���:|�<:p=����Z�=Ol4=�N=��?�-?}	c��X�;���e��J��<�Y9>�y�>�q>�tz:�d���Յ>O�>��4?���>�e�=�𰾑оPm�.��=��?%~?d�>��r��ٞ=�A��Uݒ���$<z:c>�,��i��L�߾�z��?�<���>w�>y*>`��=��_?F$W??�?�\=�HA�? ��-]��\罏.7=�D�><1�>�k>�Y���c�,�r�6�`��7�s�:����P�=J��<�:�=�*>�>äX>zV�����I@����= q��ǡ�>���>�?j��=�K=(毾����6L?�_��
Q����Vcؾf� �X:'>M*]>}�����	?������y�<ꢿ/.=�f�>��?�k�?ْc?��	��b>q�e>�� >2X<�a8��!�����QG>P��=��}�fɛ��=�7h>��>JýPGƾ�׾�9��dr������� =P�.�<y��z.����%���¾��]>�G�o�-�Ϳ���]S>��r�U�����
����ʎ���3?�Jc?l���e��x��zw�_�����`���<)��>׾�Y���Ϳ��:��s���v˾��I��iK�j�pn>�<>
2��N}����z�fS���p>��?���k9�qSK��A>ؽ��L)�>��!ß�?a��9���(?��"?��þ�|�H>�ͭ=wV�=LT�>{��>��ݾ����̪>&�-?�?�옼��V�w`k��F�ˇ�?�ɥ?��\?�[�Qvt��q���ֽ��>`�?j��>!GO���v��^K=�2
?�^>?��N>���1*w�) ���?��c?��,�AVO>���>�]�>"�*���f��Y����}�=|�`� >�oi>#l�<�Y���/��ٛ��l�f>e�>��)�Ǿ?�>��پD�H��_B�͛��7�@��+J<�j
?���Ʒ�=|*�>�>ok+��鏿�����
���8?w�?�&X?��.?� ��.������=A�>x��>��w=�@ܽ�V�>S�>U_���]��4���?kb�?�8�?YH]?�q���Ͽcl������!̾��u��ǫ=ĺ�>&�ֽbk�=��#=:��u�� ���9�>O�>�P�>Fc�>���>�$>h���(��0����h��qL��-�������,�R[���8��+�7��?�g=xt��{)=9P �vc���M�������Hn���>�۾>#)�>��>o��=<b=.��0%��@Ih��:�������(���� װ�~꙾ׁ߽�����q=�8��?�;���'<�	?�y2�w��O)�>���>f�g�x>T��>���>V�k�g�=;?��>%�
��0>�N>�����*��	�Z����!o<�<?g�;A=־�0Q��I����۾���>_M�>��=��,��E���Da�;��>E(=�8X�#-?�z�ͽ�
6>���>f��>�鑽l������L�=��I��ȗ>[{>�ͻ1��������">�m�>Y���^ >���>�/?QVW??�2?�}>"��>{�>�v�>	>��>��=6�>c�-?\�9?[Q4?��>Q7�=���3�=H,,��N�7��i^!��=��=��0<��.���ڽB�a���=>�h>׬�=K�żkז>�R�>�\4?�w�>a��>�0�'�;��JH��g�0�>K�>��'�>>,�>�?.K�>.��>d =>ۓ�������̦>�>>^vY�� O����<��^>��>�T?�?Ҿ����6�y � ��=5t�>���>P*I?I>�>�5><���J���ؿ��J��FF�F��=�\�����~�u��|���>6Aܾ��޾A����?ͣl>a�>M�>D��>[M�>���>e�>z�=x�=1J�=��v���L�f���f�=x�[���>C1�<��o�}���	�����yd���� >��?�?�$��\���g�D���.��D��>7	�>׵�>(�>�9�=>�/ V���@�T�H���>CLg?�b�>��:��$�=&X+���;��>s?�>�>��e�;m�􉘾v�<���>�?���>h��<�Z��_n�D�	�ܳ�>��=_�]�Mڗ?f�E?(B�����5�1�c�1�p��_�=Z\E���ㄾzg5���_����վE��?vӼ���>3�?��c�Oʓ>��������4珿<O��AZ<�~/���>�+�=&G��f�۾a,�
{�N�,�I�~�+�0>��>���>���>f)8?^H?�C?�d7?p	�E��>�JN=m�&?'>r�'?Z�>�?�?���>1[�>^�v�%!�8�*�~Ҙ�y"�b�>�ZJ>��~> 90<u������=�ԡ=��I�3�|����<gGa=lA��c>��>�W��^
?��&?İ��Ao��n�`�S�ޮ�<�>*�>2˥��`N���4=?�3>��>�t)?M��>�u����ᾫ�پ��ݫ�=��?�;9?�2�>��I�v��=TB޾!Y�� D=)��>�F���}�����D��U��S|>��>w�>MȞ>�2e?�Qq?|�?ϝ̾��$������=���=.����>{T�>��=��tR:�r����<G�ȇ5�6/��N�9��oo=3��=��d>��>�">�Z>�v����=�G���*>�tZ?2�?�?�P�>�fD= $W��m��d�I?\����i�U렾pо�C���>c�<>V	�<�?F����}�)
���G=�|��>��?���?�>d?i�C�'�	�\>MV>/�>�./<Z�>������o�3>��=�~y�#���;V]>Hy>+�ɽ��ʾ�1��rH�@綿��Q�~�H��9��o���E���g���, ��G�=ڕ"�Y���l���l�<�N���р���x�� ��Կ�	��?hؘ?t��E���\�ݯ�%ϟ�n�*>I���d辥��&�	>u���̾�bؾa2�O��w�^���bT>��'��>��a��)?�m^��u=>�w\?�M�����a��O�>�|��
�=xŞ��z�y'��+���*�k?��?�־��]&>���>�:>�TS>zrW>-��'YE;�S?�t?	k?�����P�g�[�v�I�u��?{�?��??�L��4A�x��s%���?FA?���> ��μ;����2?��7?�j�>L���O��SI�T��>��[?)_N�oPa>m��>���>�x��͕���-������V��8K:>JK=�}3�#%h�1RB���=Ț�>�Cu>�2Z����
�   �   *�;?���ƪ���1�ѱK�	�ƾ��}�v�>�O���D�=�)�<㟾�jO�=!��l��ڡ�=r�4>=\�>ϐq>��>V�>Kb7��ޭ=����_P��M�=鋠>�&������F�=��0>�h��C�%�OjW��O{<&�@=���=`�=��>n�J?R۶>�=?D��w5���@��$�������-��^�=ҝ�>4}]=�ꗽ!����%�V ��?����������u>�ێ=���=��u>���<�+ܼ솩���Ͻ&���0V�z�[����=!M�=���>/hּ�����
��Gb�@�Ϳs2���dp����b�����>ra��w+��N>��3��(�����>B��>�t> o>�a�>���=�`z⻫�J�3��o=!��u�������A���"����Z��=�I}�HJ�8)@�����L��� ��/<��"`�ש�v �}��>�VI>�2%��\?L
?Ro5?�"��>߿�
x�=e�o�]Q�>&�>�>�k>��>kq�=s�=3����h=�
�r=ƺb��<>��>>�=E]<�hm>��1=Ƭ=;j�<F^=s�=�K�;�O�=���=��>H�>��"?Q�o9ᾈ�例7A��ʊ�K�>J�>��;�n�B>�u^� S�d,��������T�>�>V�?x�>K�>��r>ωh�����K�ýE� <X^<���=�k���s?=f��=Mj��<JN˽66Q�ޟ];�y�=@��=&�"=SSE�|�r?��?O|+?/0>cgξ��\��������;mؾ������>\��><��=�­Y���H�D*��w�5�W��_>��D>�]x<�E�=�_<{�ʽ>`<��=�e��� �<�	X>�>+Z�>h:s>N���ͽ�s������ΰп�a���ǻ����'�a����WX��j���������R��]�=j~>�QN>���=����/�$��X��COq:�ˠ�-D4��Ng=}HH���о҉�Y'پ�%ϻ�R�����g���L�@�}����^�C'���a߽�e��K�J�\��>Z̟=�>�8-?]0?�X�>%(�����>Y�=;�9>h�Z>�'�>
 ?���>��>��=����۽�s�����=U�>*:>J�w=B�L>�｝�<�r(=�/��N=2��	��<��f�^t�=�uJ�S��=W|R>��?n���F���� ���S�l����Wr>>8#?�*�=�D�>�>&饾(V���^��~�>�vw>+��>�S�>��>�÷��0о��R���HD������<%�p��]�=�L�2�==���=���ȹ��6�]��W�=�!=���=8�+=d�f?�g�>u'?�(>�Ͼ��J��U>��;.����������J>
�>^3A=���5s��0Y�a�b�b$�*k��şh>��>/�>?Y>&M�<����gW�g]�=��Ƚ����Tg���=ϝ=>�>��>/��w+��ž���z֭��1����M>�<h�=~ۈ�e�;Ě���<,��E���"�j��=웧>��Q>>2=
����Q��|m3>���=��U>�a!>��=>Ւ����'���[ J�\+����o�!$���3��Ȋ�9{������%��H1 ��#9�jO��`��<	8�>�=+6�>rH%?��?�<�>\�3��>[Ca�@)�<�
}>�#>R�>_��>F	<>Eګ>��>��g��P��Ljk���i>
�;=���<� �<�}>�0#<��<�v=&�>e�M=����=�m�U	��f����=�;#>�� ?J����¾w�	�]�G���h�M�>�>�>���k��>��Z�ɫ׾`C-��7�Ͳ�=���>�X�>��?ƭ�>�T�>��$<z����X�ln۽ڤX���=��>�JJ��:�Z>��>3 3�{�������xɻ�9�=���=Y�>�F�=EdU?���>�&?`�<�Lξ�s�	�̾�����ƍ��r�=�9�>��>��=��ƾ_!6��D�;�-��i��h���*>�?�=7�>yz_>8�1�1꽻MV�h2>!nU��kJ�ID�c��=d#>f�E>��=��p�3��+߾�X῟5���mZ<,�~��p>jcy=��q���6����>Pí=�L�=8n>�IF>8�>LO�=�C~�)Z��t�G��1!>����;���=���n���")������꽇�p��}�W!����
�����')� ���-���Ľ��5�
��lS5�>?�r�=��>��G?C�?	ʩ>�J=�a�=�и�w�ѽ#�J=Н>���>�u>Y(=�1>���Z����L��n"��7>Y^d=,y�=�*>/ >ںq��ƈ>���=�ֺ<H�<�`�<���=G��<�%n=��'����&>��?Z�2�w$������v=�0�o(�ŭ�=�/Ⱦa�=��� �	K%��{޾#��>���>���>$7�>�->��>���8ȹ����d����H���4|;<d
O=\'ѽ���=_.s=}��=�$k<�_��g۽D�����=���=��X>Z��=<W9? �?���>�r��� ��ξ�Ӿ�P��MU�<NC�$��>�?�>eR�:ޟ
���=�45S�9L9��I��e��Δ>�b>Ow7>N��>(��=˽��=��(�q�޽�˵�i5��a��La>�{�>c�>3aĽ/F���Z���iw����=P����;���侴L��쬝���>
�B�̏���V��j=�o�=`�F<o���.4��x�� ���KS�G׽^Os<K^d����>a���d&���N=���꨽C[�t���]��,���������Ys�V�w���|�Լ�J{?�6���>�Q?c2�>���>q�s>���>���<�2>��>�p�>���>��<`�2���O>��	=ҏ�=9�l������<>�=��c�(���}=M�ĽR�E>�ʰ�k�a=9V�J�-<��.�ӯo���=�Y<�=��>H�8?��4��@�.k�$�G�|p �֦���>�Z�=.İ>;�=Hg>��˾:�Պ	�v�Ǿ�Î�y�\�茿>��>j�>����O#�L.�b'�<K�>��>>����;>>����=��P����<�f�<�f�=�2W=%7K�#=M?�z/?�.A?]<�=ʶ���j���>'�w�<�>X>�9��;�*�z��.�ϾE��QJ�s���,��=]��=pMx>���=�=O,�<�T���Ϩ�u�>U?Y��H>�6o=L�=%�->Fl9=��=I�%=�54��\x��Zʿ���� z>a�r>��<��=�j=�t���i�L���
�*��C��	��U�>3Ͳ={�9=?�I�C�=�?���VB��߽�ϋ�qր��0��\�����bʻ�z��d����������S�v�5���-��y�&��,��_���>��<?ｔ>�Ĉ<=?�$?��9?���=7�=��E�_ل�����a?Q��>r�'?�=?�"?�:>�ߔ�+�P�D���e@�>�h!>r^�=.?=U�d>ІH���6>3<�����<��_<��4�d�=��=T��)Bٻ��=��=H�8?��4��@�.k�$�G�|p �֦���>�Z�=.İ>;�=Hg>��˾:�Պ	�v�Ǿ�Î�y�\�茿>��>j�>����O#�L.�b'�<K�>��>>����;>>����=��P����<�f�<�f�=�2W=%7K�#=M?�z/?�.A?]<�=ʶ���j���>'�w�<�>X>�9��;�*�z��.�ϾE��QJ�s���,��=]��=pMx>���=�=O,�<�T���Ϩ�u�>U?Y��H>�6o=L�=%�->Fl9=��=I�%=�54��\x��Zʿ���� z>a�r>��<��=�j=�t���i�L���
�*��C��	��U�>3Ͳ={�9=?�I�C�=�?���VB��߽�ϋ�qր��0��\�����bʻ�z��d����������S�v�5���-��y�&��,��_���>��<?ｔ>�Ĉ<=?�$?��9?���=7�=��E�_ل�����a?Q��>r�'?�=?�"?�:>�ߔ�+�P�D���e@�>�h!>r^�=.?=U�d>ІH���6>3<�����<��_<��4�d�=��=T��)Bٻ��=��=H�8?��4��@�.k�$�G�|p �֦���>�Z�=.İ>;�=Hg>��˾:�Պ	�v�Ǿ�Î�y�\�茿>��>j�>����O#�L.�b'�<K�>��>>����;>>����=��P����<�f�<�f�=�2W=%7K�#=M?�z/?�.A?]<�=ʶ���j���>'�w�<�>X>�9��;�*�z��.�ϾE��QJ�s���,��=]��=pMx>���=�=O,�<�T���Ϩ�u�>U?Y��H>�6o=L�=%�->Fl9=��=I�%=�54��\x��Zʿ���� z>a�r>��<��=�j=�t���i�L���
�*��C��	��U�>3Ͳ={�9=?�I�C�=�?���VB��߽�ϋ�qր��0��\�����bʻ�z��d����������S�v�5���-��y�&��,��_���>��<?ｔ>�Ĉ<=?�$?��9?���=7�=��E�_ل�����a?Q��>r�'?�=?�"?�:>�ߔ�+�P�D���e@�>�h!>r^�=.?=U�d>ІH���6>3<�����<��_<��4�d�=��=T��)Bٻ��=��=J�5?5B���:�C5��5���Ǿ�=2��?�����=��>^�,>̩޾�h��L;�ש�������w>"�zP�>ԥ~>�V��'����������<�o�>|U�\Jl��f��<�ż�3Q�H���j�klo�x�={A	�3�K���=�v?��?��2?ыQ�8��/($����Oн^Ԉ<�e>.	�>V��=�� ��,�YT$�Z���[Ӿ�
�ɖY�AX>��Q>��U=0>��=[޺o��;��Y>e��=���=%�>�I�>e�$>ȓ�>k�5>x��=��9���^ҿ[����- �X,����O��Lo�=!r���q�=@���=�5��L�<�̄W��U���=z6>2��=e{>�Î�t���	�d=�
�<n�"�ԡ��i�Ѿ�`���Sؾ�1l�K!/���!�C,�"�P��_3��T���*����Q������=��?� �>�@�>#:(?�m?90?4*���>[=�ԅ�r`�=���>Sr�>$k?1�>��?��>c=~Y�==˽�� >�Z�=�I�=y<�$>�<g��'>�-=�i0<C��;�*�=�= =�̠� X�< ��=�P>�?X,��M���8�ߦ$�n�H��`�?��<�ʽ�m�>��>�|��,ҳ��I+�l��������=�>އ�>� L>zľ�U����E��ɔ=��9�,B=�T�v�����<�>>��A=�P	>a��=3ƽ�^=B��q�<��>>���>[?��?L�ʽ�%�� �b��������)�fQ>4T">�<�=΅��@ʹ�����"������>�)�A<F>D>1Ј>���k�2>�J=c���y�����=�=Ͽ��F�P����>�c>�|!>�ƃ>� �:
罣=˾�οK���[t�<��=�e�2NC��t%=��߾��9 ����Ӿ��E���I���gw>ͶY>j�a3��t>�<׾� ���h���,�wqs�(EV�Hhv�IȞ=)ӽ���	���;1��+d�0���|���9�i����r�5;�Q�/>k�?X�0>�QS��~A?��2?m!0?����Ǐ>$x�>����I���>�)�>��?`�?hm9?R>���y�ҽ��l�5�t>�%>]Q�=�X�:KWW>%B|�u<=�!��>7�F�����"A=7�=���=�ߛ<��=��U>>��>�\6��o�����
�
�2����g��>�Aо���_�վ������;��6>�A�>9��=ҹ�>��r> ��>�Z�>2P��E��;:�=\�2�6�@>��=�Uj=od�dh�=�-��4�ݽ'�=���D<d>��=sm�=%[->�x'>:Y?ܒ?6�#?t���������;Ҿ����=���>?*>"��<|@�����7�*��農�־FT뽸�l���ļ6��>DX�=��>�� =0#ý�P�g�ͽ!��=��J>B�5>I�E>LT�<iĆ=��Q<���=�F���ː�ҿ�b�~�w�!�vv>+&�>�"d>�F�=�!�>�{>A)�{瀾�1���V�=P�@>S��<������(C�;y����课b�"<ER��ݽܾ������1:��	zj��C=��������j���ƽߗ��'��YU�u_!�q���t>8�|>)A�<��=��?���>M��>����s?>-�`:$��>�}>z��>�Q�=s/�<r;>���>jM�����s����$�h��<!}�!�B=G�Q>�K>>�,;:}N>������ƽ���W�=�#>�?=�	=aw���2�>�з=y5�>�A�<�h����q���3����������>�Mоܜg��D�9j�iA��=ƍ>��;>m>ci�>6�?�Vs>'��>.MؾN ��OU=��������������=O6>��=�%j=��˼�%�}Yw���1=f�=-7J<���>	?���>xy9?�S�k����ټ��̾׍�� >���>�t>���<��ݾ/�,��2�+}�J�=�1-u��^�=$�>+KO>܄_>��=��1>8��=���>4��<D���D�8<Lq�=Nk�=A\>T{>���pH���ŵ�u�ۿ g���>���!*�=�{�>6�6<ɂ����=��A�`ڷ�F���0b�^�7����E�L��O��]�w��rt�0��Sc���>
�_��q˾�g��-�����=z�h< A�@���i��A+�e�ὑA¼3��=�k`��˽A1R=Ɔ>T"s>yՓ���=�(?p�>�@(?�J?q�?�}�>N2+?�'�>��>�6y=��=���>^�
?x�f�hzþ9"0��s���Y�=�E=�=�T=P��=�]/�.`��|����<ה�7�9.B=��<R��Y�"<��>ȍ>6�?�J�=d�陗�G�N�羛�>�+�v�0������'�b�6��2�)��>pq�>���>�H
?{T�>.�>��>TN�x�<�0'�^3��Ө^>w���"�SE>J������I�?��=��;�>��=�?�o�=R��>�\8?�!H?��=?��'��V���<���ؽ��$�X��=�J>>FM>.�>����*�I��
�A�08�L価�o�-i>S��=! G>Mj}>���=E"����=)�'>�M>���>��]>v��>�xq>$�'>���<}�8%��Y�Z��O��Й��b)N�V�c�A�W>ܓ�>��Ͼ�X�%�?R�5=Ɬ<��g>��<KL>8�>`~<���=ڏ5��?�<��!�E!���]����7썾��<�#U�D�>���}����W%|��z/�j��L!.���Hj�N��2KD�዗>ᝏ>�p>^�>_c:?���>��>�^>��>&��=",�><�>�P�>r�?�ǒ>]�=��>�G>�������Q���.<=q�齂X0>/�K>Z��=����T�=�z.�&́<�$G>37T�g�rл;�'@����=W|�>���>m��>1zu����������(֚�!��q��=��:��p?>�_k<m��=��z���C�|DS>`�>t��=z=�ѹ>�)�>44�>fGO��`�=� n=h󜾰 +>�6<��Y;��>sv>��һ��E��.s���g�qd�=Ž����q���m>�.>�(?h��>��?���b�&ݾ�;�������ط=��6=N?ѼnhE�M2ݾ��.V⾚��R&���;��r�>J~>��>%;z>�;>��c��JJ�M��=����ܽ����qU>�@�>�:
>ڌ��J�<IxQ=��6`ʿk��� t�v@���U'>�1?�>f�g�*锻چ��v¯��tW�:���<�=� �	p���	>�[>���^﮾���lR�=�`������v���g	
���Ѿ���ш�����暽N���������y���������='
�>�]y=3F>�-�>*�>K��>�'�=_;�>ܳ-�4>g���W�=���>�YA>��=ѩ�=\�=��X�}�?�2��=��݀<Ƥn>f_�>8�>�]>�^��x�N���,=���=>�=�x�<{�E=g.>�<r>�V_=m��>1zu����������(֚�!��q��=��:��p?>�_k<m��=��z���C�|DS>`�>t��=z=�ѹ>�)�>44�>fGO��`�=� n=h󜾰 +>�6<��Y;��>sv>��һ��E��.s���g�qd�=Ž����q���m>�.>�(?h��>��?���b�&ݾ�;�������ط=��6=N?ѼnhE�M2ݾ��.V⾚��R&���;��r�>J~>��>%;z>�;>��c��JJ�M��=����ܽ����qU>�@�>�:
>ڌ��J�<IxQ=��6`ʿk��� t�v@���U'>�1?�>f�g�*锻چ��v¯��tW�:���<�=� �	p���	>�[>���^﮾���lR�=�`������v���g	
���Ѿ���ш�����暽N���������y���������='
�>�]y=3F>�-�>*�>K��>�'�=_;�>ܳ-�4>g���W�=���>�YA>��=ѩ�=\�=��X�}�?�2��=��݀<Ƥn>f_�>8�>�]>�^��x�N���,=���=>�=�x�<{�E=g.>�<r>�V_=�\?�>@��Ȝ��;l?ž���=d}�>���=F!��ws>�N>[O��~+���@���W��[���H%>�t�>�=�>�4����4�U�=�ܻi��<�~�=��
>]�=1�=x��bi�d�='��/��=�N>7h�={̢�ݺ#>G�5?u�?��?�@��vȾ���5lؾĩʾ�����=�Y=�0@>Q*�<�Z��ɺ�R���q�!�ϣƾ�y�IB>�Q>�ʨ=\��=�;��<ϴ��:�g]�=�1z�:��=�%>.�>&u�=�w =���<�2�����<�Pƿ�����!>W,��Z��<$��>�J����*��k�>�u��F����D>�\;p���k��=��i�ڽWh&��%�>� �Z�>��>���������l��wܽ�T���Ƀ=�8��h%�<"�R��1��ۘ��Ʈ6��Q7�����YJ��!t>aw]>���=�E�>I�?��>�a:>!>���=��G���=+��A�^�&�P> �>[��>�S�>�g�>O�=��c�hWv�a��=n��<��}=�ߋ>g>�>�����=�-=Z$�=H�G= >Z��=�q�=���n�ݼϵ�=�Xw>�k;?5�#�����2��`V��¾�G�V&?0��l
>I�D>�]�7����㽾1�=U̾�Ȉ����>s��>��>��n>�c{��ֺ<�}4�{�9>~	x>���MSV��``=�yR�U&>S�>�t0<��,=�f=�+���.��X�>��&?�!?��A�.�I�r
�����ξض���3��k>�B,>��
=Uw��*پ^���4�W���I���[>F�>Qsc=��A=�S!>��9��T� ���������<�c@>��>�',>��*>W�<�%<֙>�0<a�п����U�b�Ѿ}^�^o>��K�0��(�d>�ؑ��g��Hr>暮�͛�=��>>i9>�y*�%����A��6���톦��h��#p��v��zm2�d�����#��}��]�l�j]��S��<�9���q��l�u������ᱎ�J>��eO�M�>�7h>� �>�V�>/|�>7�t>�&D��W>h[�<�X�<_�����i>j��>�#�>$s�>A�>2�1>*7�m7�_c!��Ը=a�=\K�=8�>ݥt=K�N�3\�>��>"xL= 宽������}���<��=O�=�1*>�>]">?a���� 
�#���Ė��ϩ�%m�\>$?<2�>���>:�p<\��H֨�(���EX��4Gd=wl�>r�>�И>�Ȋ>|pξ�����=��->J>e^�>O�=��v�B}�=u�D�	��=5��=�P$= �=O=B�=?�<�(x�5��>��/?�2K?厥���Y�h>��� �񯿾����Mb�h&>P�r>.s�s��=����d��$�/�+F�:���6 <K®>�!>ᢜ=��8>>��W���:��3��vȽ���> #�>N��=Na=�>�c�<Okk��A���ȿ�ĝ�y��;O�C�� P��1M�� �̬پԥ��稅> J˾̠��^��u��D�<>���=IUc��S�hw�K½�ᶽ> >���=�������yž#�5��4��a�B<;���v��������ڡ�g�k�
a��i硾E�]�����>;>�=jN/>v�?��>���>���C>d̐�Q5ݽ�}����>6��>\A�>�I�>���>I��\u����a��~f�q��=jƂ��	�=�;}��`=�����WG>��I>�#�=;x��U
��Pսcʼ^n����=l�=ޜ�=TW)?#�����"f-�K
׾����[}�=\y�>n��>j����>���o���_/�_���(���� �S�>b��>�^�>��>pI�H;`�Dw>�S.�u��=� �=���ʒ�������=B%Ľr�;>���<r*�a0[���Z��4����?N�?�I6?��@��rԾU�'��,�N�Ծ-5%>#�ݽ�'�I�2>8x�=�:=�Aþ�Ҿ�Q�����h.��m>A��>s�\>��E�V��=�;�xI�=!S�=�{�=Q�>���>�R>U�`>̡.>��B�=+��%<�wƹ�C���x��>`)=&���x�>�"ɽ��׾q����=���F��Og�=B�>��=�G���G����|�eG�:ܾ�-4>H�>����	v��M߾�:��������<B����/�?��$��%��X��IOU�+��M[���>D�?��63b>�b?Y5�>jm�>� �=(a�=׷x�̅�>�܌>�K�=B�>���>il ?1�>�>�=����=|j���I>����=���=��\>��<�\>��(���*<T�ǽ����Ҩ=Q�?����<Bp�=p!>��=Sy/?����a	�����}󾀸��'�Y'?��>P&�=�	�>:���RɾܟȾ��پ�`A����=�_�> º>an>j�>��;����Tx��_���>���=n��p�˼PtR�V�<9w�=�e:=�V��S_�=~Ƕ<������>JI�-�?��5?�T?$�l���d����<��Užcb�<� X���^>��><�����^;�R�JY��a���{¼$Mz=Oڥ>V�=���=F�&>�ܽ<�"<c{|���X� ���I>�">`ʈ>�.>��=�=���=zH*���ſ����!�=un����M�T�*����ǾF�]�C�>7����Wܽ�Qb��o,>�O�>������I�  f��Á��j|=#�< ��=ۄ%>�Ͼ�r��뾁����������<b h�M�ݽ}�5��"����%��u�<���j��|�Z���<Ӆ�>��=<�=��?���>�z�>��C=�:�<0RT���(�=��>�ٟ>�գ>Vh�>L�I>@G��[S=�9��d���E.>
l��Q8V>��=y�>���=HB>���<�F>�ʌ���ͽ�����}�<%Q~����=O��=��<��?_@�>I(���:�>u�#�>�� =5��M}C�����Ƀ��=TN���j�ȳ��'>B!??Dԃ>3R�=K,�>��>��d.��z;=�����Lr�6p&�?�2�=1�>��&���,�9�VtϽ��o����=U�<:��>iD?��?T�m>9����(�-�۾LSվ�7���=t��>�>&��=�쒾����A$���N���^��F�b�����<ڮA>�:˽A7ͽ�O�=쵓=a>.
r>rH��>6>cV�>��>��>"�e>�45>��=�x��T�w���Կ�S��%��?p�����=��������=�E�<�5>uJ4�}��]b�=��>A�b;�Y�(�˽k�0>@#>@4������U=��������#"�Ygν�!��ڽ��~0k���Q���E:��սSF�7ф��z���8�>��ν�
�>� ?�w?<�>��p>�m?�3?B��=�1R>׎#?��?��>��=P�ɽ���;}j�= f'>+h��sD����^ B>�7>�a�>N�%>���=U�=��6=5��.��<�tE�c˘��D�<��<�wS=��F>��>�]?~�,>�n��('��=�=~�ɾp������Ծ^M ��pC�����I�=���>oA�>B�]>e��<B�U>E�>� ��2�$�L	>��B��?'�մC�+}��ݖx<��A>;����ӽX^��n8��<�֒=�s>ؚ�=P��>uv8?T��>F��>Գr��\%���ݾ1���n��.�6>r��>�Gf>���=�����3߾��f�8�r�@�w+��P�_C<�<V>�
a������<./�=�p�=�i">�H�=�>�\`>D߬>��>��d>@� >�vf������Ϸ�}ؿp@��a���G�I����=�>I6R>��=�Az>?�k;��ľ��(���=�tW>�K������Ai}���<��.>���=�fW�e>-5Ȼ�J׾����%�7����)>>��HC�FQ��~�{8d�.;��������D�o`[�ǡ9�C�>���=G1�>�>��0?�F�<)F�>>�?�
?W_�>��>�_?i�?��?GW>�\��������^>�(>�^?�s�q�#��=�q>>i�&>X�>�_$>�U�=ޮ>"GO=GA��%E��D	=mC0=��k�����=��I>�$Y>�J?To�>
�>�ÚW���`�9ܛ>�~��⏾� <�xA���<�K�K�F�[����t�=�H%?g?� ?5p�>���>q��>�����a���L�]_�����*wY�֍&��{e>+�<����e�;����������k�μ�w�����;�>�$C?�.?��>�d��!6�]B����=˾.kH>%K�>o��=33g=8R[�aP����^C6��[X�kM��j
�(�}<��s>���.ln>�ʫ����^>�׍>ۭ�Ǝ>��>�$F>;�>>�>W>�>�[-���Ѿ�dۿB���=�0���=m}�=�d=C8�;�f߽V�P�7�оn�~�+��=�R�=���5��:��|���/����E�L݃���=F�X����^��<��w@.�lA�xK"���.�SFl��Ⓘɸ4��,����J��U�1�����>�w!�|��>��
?��:?*�<�&?�V?�1?��>@�>� ?��?<�?�1I>�o������l=p�C>%Y�qA��;� X>�&>��== �=%q�=��=�����5���1�Œ=*�=���<:&<=�&=�]>�n�>��?_@�>I(���:�>u�#�>�� =5��M}C�����Ƀ��=TN���j�ȳ��'>B!??Dԃ>3R�=K,�>��>��d.��z;=�����Lr�6p&�?�2�=1�>��&���,�9�VtϽ��o����=U�<:��>iD?��?T�m>9����(�-�۾LSվ�7���=t��>�>&��=�쒾����A$���N���^��F�b�����<ڮA>�:˽A7ͽ�O�=쵓=a>.
r>rH��>6>cV�>��>��>"�e>�45>��=�x��T�w���Կ�S��%��?p�����=��������=�E�<�5>uJ4�}��]b�=��>A�b;�Y�(�˽k�0>@#>@4������U=��������#"�Ygν�!��ڽ��~0k���Q���E:��սSF�7ф��z���8�>��ν�
�>� ?�w?<�>��p>�m?�3?B��=�1R>׎#?��?��>��=P�ɽ���;}j�= f'>+h��sD����^ B>�7>�a�>N�%>���=U�=��6=5��.��<�tE�c˘��D�<��<�wS=��F>��>�]?~�,>�n��('��=�=~�ɾp������Ծ^M ��pC�����I�=���>oA�>B�]>e��<B�U>E�>� ��2�$�L	>��B��?'�մC�+}��ݖx<��A>;����ӽX^��n8��<�֒=�s>ؚ�=P��>uv8?T��>F��>Գr��\%���ݾ1���n��.�6>r��>�Gf>���=�����3߾��f�8�r�@�w+��P�_C<�<V>�
a������<./�=�p�=�i">�H�=�>�\`>D߬>��>��d>@� >�vf������Ϸ�}ؿp@��a���G�I����=�>I6R>��=�Az>?�k;��ľ��(���=�tW>�K������Ai}���<��.>���=�fW�e>-5Ȼ�J׾����%�7����)>>��HC�FQ��~�{8d�.;��������D�o`[�ǡ9�C�>���=G1�>�>��0?�F�<)F�>>�?�
?W_�>��>�_?i�?��?GW>�\��������^>�(>�^?�s�q�#��=�q>>i�&>X�>�_$>�U�=ޮ>"GO=GA��%E��D	=mC0=��k�����=��I>�$Y>n�?�\���*�
�>B�M��7���Y����<r�v���?j�=�	��U���)�E*9�����bPh>4?�ų>`?�>��s� :2>UE>���=���=R�*=�2�+�z�1��=�6j>:�.=���<�Q�ۡ<��G�A�}>t5?ց?�A.?�V����$�Z���F�#�H=ƸM>2LE��p=�݅���߾(�����Ⱦ�ǝ�Gh��k)(>��s=+G�<�#9>��6�=��QJ=�=@^��t8Q>&�M>�G�=?2�>ύ�>{��=��ֺz�;��j]������͗=����N��\�>:ѽ��H�^����b�6���͘�=�����=��Β=1p�=j��=���<�X=��u�����.d,>�d�"2+��&�=����6�<st�����=�qP���0�O
��9;��Rk��<f:ǘ��b����μ����>nϽqZ���l?�Z�>��#?�>Y�>����М=M�>�>*M?k�#?�
?��?Wѧ��E־�u�����s�>�	|>�K=�]=�A<>���\�=z��;|�=��=�<��8	���Wr[����=�A)>I>3+?����{�=���Y�7�6�M�.���޽�r�猫>n�� K���1��w�.�=~n�>�3�>R���1e����>"4i>HZ��R��?�Փѽڇa�{��=���=�������=���=%lR=5���DT<�2�<� ѽFY���;�!f>�T4?�� ?��>7���k �	�λ��"���:z�z�>��?>/>�S�n���:��c �*�b}�����Z�>v>�>>]=>��Z�a�!=�˪=��Z<'��v[�=�q�<Ca�=T�6>���>�z>q��=�˙���L�p�F狿���������>��=Y������m�f�щ�6j��t��0>��?s��=RN��`�"�>cR>�,ƾ󄩾s����G!�����x�����׵��땙�Z��"?���B���l�_e���b�"�N�H1]��e!���4�k���Y?�B{���=C�>�>">�?�,�>��>��<�w��>��>E�>(�/<�a =1ޭ�ު�<�(>?#G>���F�˽�0�=�2>7nH>��3>=|F>�ٯ�}<�Y�=�Sl����i�<y	�=���Nߟ����=���=(�=�)+?��������;�=�(d�M �>��Ծ�� ?��@*>�/�}Cf��c�`S$��	c���?��?�(>�e����>�<>$龘��=;��qcؽ��W���=�{�O.=�I[>����Մ��߇�߉�:Z5��q>=)Pz>!�>��>�AW?FH�>"?�"��oW���-��RY��&��c�N�p��>iJ�>�ҝ=`xڽ\�����"���J�X��H��E��|G=0��>Xr[>W:�=�=<L>���=�/I���]��_>K;c>8�>�=���>�4�=-w�����ԃ���\ѿD�����v�FIp�:��<���=�Y>���J�=�����@��>	>#��>��>xQ>ta�<�'�˻J=�c=:~�w�;��N�=�^��?�T��NQ������c�0��&�%�M
���[#��=���f!��.�c�ܽȵ ��r ���I��J>��?��=z+>b$=?m��a�?�|�A�C>C�= �>���>2��>8�>��=2��AǄ�&�>�t>���H����=d�$��k�=B91>�iQ>�᩽[�U>�:�=�^ �M]Լ�m�=.f�=�����y�<G�=Y��<C��=�I/?������Ѿd>�{��F���9�8��>9��Ƀ�=���#.L�*+��r[���!�T�;�l�>�#�>,	��*�>h:�>z1�.௾�����0;Y�Ž	�>�9=����C�=�y�=�X�>g}>'p�>Yd]=�Gu:�Ks<����P���,?�~4?��3?�x=�l"�7�A���Ob���Z:�!ڢ=<ֿ���3�`�����������Fʾ�U�</TG>sL>�ج=:��;��Y=a���s-���=|⍽���λܽV�<U1�(V���=�#�wpǽ��X���޿�lT�:��6�=��~��->����˾��q����� ��=2��>�S�>��޺�-��7�
>�}�=�L���yB�-C�=?�=�$>I�V���ľ[{���� �qw����=�%�kj��r�����[���}&�E ��nQ���T��vK>2T�>���=���3�? 5D>��?Ge>�?S�=��>Zg�>;��>@��>�|?�\;>���9)�y�>�B��UR��z:�>�[�=m�=
>�3=>}�Ž�8�6��5ѫ=Rz=��뼯�r<�ཋ��<v�=�ȼ=Q>' ?ZSо�=#�7��>�V��Z�>KI���+?X ���{�>U(��!W�{�e�.�־/���R?��?���>�䆾�5�>>>f,������HM����E�ڽ��1>
�,='�	>�fu>CH>YQY=�ܗ=�<�+��o�<B�?>P�>�7]=�9?�b?��$>B�ýT���-^	�K�򾱳n�t����>�x[>�->3=S����aG�,�6�+
?���������{*>��H>ue�>�R'>�ez>2��=�`6>q��lD_�ɷv�d���	ξ��m�=�٘>��8>1}�47���^��\ݿ�Ъ�!����N��&=OC�wŚ>R����e��2>�㉽�>��0>��S>-NA=OU>��=)Q����=����9@�s�=�87�����P��`����"�ΘJ�e���Mܽ@v�=��c�����dU��;SV��Z[��H*��,B���K>4?��
��z`<=?����@��>]�O"9>pX�����>V��> �>��>۷A>��m�;_��/>|�>4�"��'�TS>�D��=p�=ў9>Ap�P!�=�|�=����cX���3���k<o���82=��>�&�=PU�=�? �F���M�e�[�������
]�>2y��T
��'.>�=g!���!�� '�c!��Υ>>9��>�t�>�0�>E�#>��;��l|�@&��Ҙ,�P��6�p=Kܣ���=����cP�=!�=�|����f�����4-Q��~F�uv	=�^x<�!5?6�:?u��>�d��I��s�� �3SѾ����pM�������ѭ=A4�<�U�<��jK���H�ي.��A�<t=>E��>���>Y�g>�|8>	H=���=����s����=��=D	<=ܴ�>�p�>��t>�5�=��|;����ܿ�Ⱦ�da
�Z+	��:>>(>�O�=4#Ӿ��3��??o�=�)�
:�=���>�C,>���>Qm=bv?<��B��S󾐜��^g���5�f���w�0�֋�0�U����^
���*C�7TW��gG������%�bTƽ�mQ�4������;d=%(?q��>R��>a�D?d]*?�e0?��Z�/�>c�������^6>��?`��>�?t��>�7>��ȼ���=�!7�����q�=��a�{= �>>�D>v�ҽ��=��=���=���ݹ��ȵ��$(�x� �yԲ=q��=�B�>$?U����gѾ��N�"� ���߾�,�w�	?�����d�=��>�}F>(��P�1�V��(v��
>�?�5�>u��>�Y(>��\�����:�G�<�s<�ZN�=*C�=���9
���5�)>Y�>yy�=#+;�O	�*�M�ڽ��*�;�K=
�"?���>ϣ>vJ�{��@��i���O��s
!��^�H�޽��y=:ة=�����"��:U�]�M�C�6���	�hGR>�-b>vy�>=D>I4��$�>��>�����=�H�'=l�>�Q�=��B>��>�K>���=�C��._Ⱦ�ԿOP��Dw���+��}T�w��f�����B��'<��$���̾j&�6ǘ>�ܩ>�j>Z�C>Nڼ_� >��j�w�s��c�P�݁�b������	����~�e�De�u3����{�aN>����aҽ���p^��$�Z���9}(?fǝ>=#aV?��C?��S?=�=��>��E�$3ѽ�(�=�_
?l?�?��p>-q�=rO���߽�y9��'����=��9�I�=h7�= ~<>��ƽy�o=�>$6�=ಽj��#?�<_a�|�=ng>�>p�f>?�?̈́ؾ�K�P�Ͼ��43پ>�5�ل�>G�N����=�<�>��=~辙5#�e�)�B���b�>��>��>���>�>%ԃ��z���%a��g1;l���p��=wy�Lj���=0�]>��=�IF���<�_��i���=ly�=P0>-N"?}�?0D�>�n�=d�ܽ����K��������?��hI����=��Q>݄�:�^���? �K�q�����}���ֆ>4�>�7c>h>�vJ�+꺽�J�=c&���(�{F><,�=�/b>:)�>�]>T�P>�Ϊ=-��9���ӿWІ�)�.�������y�ս읏>79�M��>���>p-����ڀ�v�=LZ >b|�>V�}=�� >���Í��M��,�0�?��Cf��1��a$��j׽H���x���ʾ�ξ�q���\��Eb��K@�`�δ�Us���N>�7?�H�>Ƙ�>x�K?��?��a>��>���;����������>� ?(+?��,?+ �>�>�ʉ��zV�d�Z���� !�={>\�=	�<�OI>���ھh>�-)=WL >�cz�?}V�2���I#;�"�==]>c�=o!�=�(?�����ξ}���)%�P����=&V�>0ܵ�Q�>*`0>���������z�r�C>�ر>|��>ܚ�>��h>��>��O�7���_�g>v<��Ž�c>�S=��������%>ݶn=d=`} >��ƽGo���˥��2���R>;�*?�L	?)��>��=�ꍽ���y�վ.����ɾO��W�b�b
�<h���+�o>4�7r�rY;���vo�@Y�=�a3>�'A>�պ>��Z=�m>m>7�=h�=�nY=4P�=b�=����1�=nˊ>�>�S��d�5"Ϳ�O���P��֙>;����o��S���L/��J�>�V9�㲷�|EW>�a��	0�>ϙ.>.�Q>S:����=D*�>�̱����>=.}��ɾ6�O��̿��u�:�?������]���sy�=�G�(�7�'�:�B�/�\^�+�н��5>	;�=�K?��o>:;�Op[?J8?\�>��0>�}�>&lĽW���1�>L��>�0?Ƌ?��ϼᲘ�7h�E��,���L��*B>��!>�/�=�db=�P�>����/Z/>ϝB=8�=�����"۽�&�=�ݽH�ɼ���=�>�hW>"/?����{	��Bꃽ��C���XHk�)S?M��=ʚ>9+�>�h�>³ɾ�V!���,��c��~����A�> �>�0�>�h�==����J����ͽ<�(=&7=F�=-Ȩ=����.=@+�=�2>Q�>������%��FE�\�R�;��=!mZ>�"?!��>+��>8D*=��Z��3 �K���a�=k�>��� ��}g=���<<.;�h\��[�m�
�<[2�Q>�=⛽�>��V>]x>�Ę>w��=
<��Ԧ=+
C= ���"v����=����^ >�c�>���>q=>h���ƾ�Vۿ~���D�n�5�.>&;>�p�>��ྖ�ؾNhh�{@����3�����>�/�>�Tw>�*W<���=zw�<�k5>X���~�>�s8>؍��-���b4��ގ�=�6��*�����z�'��պ���~��aT�z����Z�b>ܽQ)�OT->K�<?ǂ�>�>(7?p+?�h>qtl�{��=�����:��8>�?��?��%?l�>�W�>�{O�����C������N=�,>�>�t=�Mt>l�$��=wgV=DA>�>=��垽�r�W�e����<\�7=�+s>4dH>"?�fa=����9=B�2��zܾ�T���
?�*�be[�G:��ˁо"�2��#���=9��>���>&?��=��}>�>R��u&T�8J#�&�g��&^���T>� P�m(�:|"�<��u>�8<��F;o(=�d�;�bV��m���=�b��З?�*/?$n�>|=q%��c�f�8�žFo���|3�cȬ��0>�r0�����k�(�� )�P�/����fm�=������>2i�>`��=�]>�<��a���=}��=�Xs>�G=u�1=M6�<4W=N:�<��=I�%=z���ܿ����)�����iܠ<�%V>�7]>�<���:Z�<�L�5���ѽ��@>'�X>ǎ����ɽ?��#��w��=�ֽ�|:8�0p]���z��N �U��t���GwR�pQ�i��������9S=�7��g���+{��p�L!d��Ѡ���R>��>��+;?���e5?��>�?��½5 ? ?j�$?�� ?�?�	?4��>�B>�ָ=�y����>[.��lg�z*�=�`>Z�>3��>=�>_�F�S�=`����ڽ]0��I�=�^=�?���E>#_�=s��=��=�%?��$>��v�N3&>��]���)�����o!?mܶ�8��7��gM��94���ޅ��1�>%i	?=?`>�y>���>}�4��ҽ7�H��W���Հ���s>��+<4B��`z�<�><R;���Γ��mH�g�C<��v�{��+�>O9?Z�?��>���,�۾�=�a���l׈��'�;9�`�$1�=0)>��T��"�O��'�&��ⷽ�]�=�b>Gĝ=���>�	
>���=QH�%E)>`>�>>%�>�>� >��(>f�>/�?�bL��o-�dĹ�p.��Z$'�N*���r>aO�>�ώ>�ܾw�۽Wt_>}�/�5j���a=��i>���>C�O��㓾9ļ�=�E1�rD��EX>֔�ƪ�!��uʍ�VN4�ӿ��)��R��������l��f8�S�+�+��5�o��B:��6׽�>[T�>�>�3�=�q?���>��?2C��X�> ?�>��>���>%�>Q��>N�u>D�=�[�<���=�+��i��U1ýpը=�X�=˪�>�u�>�����s=��<��=� ��"=��\=�n#=Q�>V>��9>���>�!�>�@��7�ƪW��������D����.>�⏾ǔ�=+�.�9��ξ�㮾nd�f�Ǐ�>ҭ�>�]><"�>O[M>��ܾ僣���C��AT��ƽ*S^>�X�=4ç=�
c>���=�W�<׌T=ڣ���>�2�<�>�<��A=ʾ��I?��&?`0$?nYT>�@U�þ�����p(r��ǎ���鼄|<,�=��ʜ�����
���(�P��޼�+F��>��'>�Y">��=��
=�%>�昽.�F�d�+�*V��5>W>D̥;�0=y����ֽB�Ϳ\]���Ü�8�Ⱦ�b> �+>O��>/�R?���F^>��}=cr?>M*n>������a%���9S��p����놔��<+��=j�I<z�dF)�iRW��:۽��I���~�����A���
{>�u�.�D@���h�_�J�P�*��5�>�JB>̴ѽ�����>��> ��u>�e?_`k�y�=m�=ď_>1�1?~�'?F
?�a�=L\�XP�>#x�S���wx>�'j>e�>x{>�c�>)�f���'���>�j>'O/>)#�=Oh���kI= �ؽ�=H��=�M�=��D?�i>���E-� �C�i~ݾ��Ҿ�q6>G�=�|��.�������b	)>C��>��>c��=��d>���>,�z>��>�7���0���T�=�&�)��U�^>[�">��8=/Z�b��=�'�<}��<�=k=әļ5S��缽xn	��!�=�#?�� ?��>Z>!w��l���5U���r=6`�<m�F>|��=�#@��z�����|�9�^*6�7���VX4�nҒ=���>��>z,�>R�B����=������>�󷼹̨=$�`>
��=���=�w,>���=��7<�W�<h~A��Xſ�	���D���]=�����>yE@�1���c�^>�>ŉ�=���M�l.�A񼞍_=�F=\nH>e���,V<�w�оlp*=��r>Mk����g�&�;\���z���(˽$����ڷQ�ѻ)��HT���O��A�݆�%�S������=���>[��>{�4?�I�>��(?���=���>U8>�Q�>0w�>~M">��/��#=�.�b�J
>�d����:��a��X����='?ڽ�햽�t�>�}�>l���	V����<���=��^<��<�.?<�f�"��=�)>�H�=.�O>��>(ݫ��C��nbW�p�ھ�x����r��=*٤��t�=mt̾֓���	�����9��==$�>_
�>h�Q>'�h>�6�>�AN>��߽�'�;�t�T���Zn�0��=m��<���=K��=M̪��*X�T&�<��i=�g=��M<ֻ�=�vO=�J1=�B?{Y?Wݘ>���;���:<�F#��="Ƽ��k>%#�>��>�Q;���������kq۾�0���[n��#�=)�>w�>�:�<8��=S����t� mG>tH��������=x��>yQZ>W�
>/�� d����y�8�þ�sʿ�ޜ�G��"K����y;��>1��=��0��NE�t3���IQ���¹*<a��=eV�<��<�T&�_
���wr<������ü�����.���x��ؚ���3�»���=�2���G������y��������C�@l��q��]��!B�>�X�=v+E>x
?H¦>R�?��ռ�v�>	����H�>a��>
 ?��>��=�ƅ;��<r�=�e潚۟�d�]�t=�vG�v�>&�=�5S>y���}��k*I���r=��|�̽�Ul�_��%A��*>(�
>�_\>|�?w�Q�}ľ�ʾ��N�-����>�U>�햾�_����`酾�&!�1�^=���>LZ>}�C>��z>W��=�_u>*?�>�����=�,����=
�=�t� ����>�=�ؐ>�+ ��D����L�N8�=$��=�M=��oL=K�+���>�$%?4��>
�[?� >t��q-�h2����W�'��$�>Ч%=�=�>����v�\Uվݕ(���/�8�#���l��e�>��=E���]��=��Z<L:��r�<�b>T��oB*��o�>D,�>-[O<�<�=�黕��<���:�0��(˿����j=�=A����^=[�>��]����?>?m�>�yg���9>0�!<��=�c��`}����&���D�>��m{�L��>�V�>9�-ͯ�B�����;9�8��q/�"���gx��J���L��
S��U������r[�A�l��=�-�>�%�=,<7>ҽ"?wz?�>{�o>u�%>8T�=dȣ>.^�=�g.�����d��<J�>�O�>!�,>��=T�'�G���Zd�<��U����<9�� T�=_<=�̝=G��=�ꪽ�L�=[u�=�>o�w;6�G�uM<�dh�[��=?��:��Ⱦ��t�CA�NP��ò`��[�>�E��g��Y�v�@q��bF뾶��YA��@��=@��=v��>)nb>�1>��>h��J׽�^��n���k���I��	� (��~��>���;�TA>�m>��� ��$�Ƚ�q�����\#>�kG?�k�>uV�>����}���5���9���<R90���>�=g>4$�>���=�R��Dӭ�cX	��+$�W"�	��݊�=�8�>n�`>/��>�V�</ �=i��d|�>2�=����z@�>�Br>�>��z>�ۼ=/�>�L�=cݤ�1˿�ԙ��=%��}�>�?�>�9%=R��*�H�=���;<�K佭@��bܽ�[��S�0=��>S�Z>2�$=�8��"D�>������,����{�������qȾ�,)�����wq���F>=�̎�9u��La���8�Y	�J>�`>�>�3>y��>���>ߣ�>&G���>mn>�~{���`>u�>��>[�?1�>�H>�7�Kw�<5���u��}��=��2��ݤ=��Q��>v,>f,�=���=GF׽��X��@�kV	��	=j�S>J�>��F>���>�92?�Y<:(%�_>I/�Q�̾5J����%
�:�Ͻw����w&���l�༇k<=I"S>��{>NA=="~>t��>�浾���=EL�׈����=�9�=�uf>e� �%��>q}ڽ�8=���<�pT�<��M=�z>(O=�f�=PM?�??�?�p1�-4ܾ�d�������/�Ji{=��3>��>��������ƾ�m.��N)���0��"�u�j�����>'� >
�>&�g>���4%�=�b}���-�'Pu�`�%>t;:>��z>���>���=ɠk=�=&< ����ҿ֡���ѾV�>��� =]�=�>M�&>H��=���>ߴ���>m)ͽ����l�)�;���`���Z�8�=�b���у��5�=��V7����饾.�D�9 ���bw�!����:�T;��+�k�E�E�y��3���#�]�^�,=>-�=)��A?�?��y>�E>%h?\L+��aY��<?4�.?�6>W�P>v->r��>��>w��>8���̊�g~={�� �=� >��=�<��+��O/>4=`�J>�w=�x��g<)#�=hjo=��1;W�>�e,?�C=�j���ʾ�'�o'��;J�=hR�>f'��^c�<^5齄����=���|=Τ�=��>L�_>���>F� >�I?>�N�>K#��v�;H]��j�'0>��>!~7>�����>�*|=Ŏ�=����IN̽��k<�qQ=!�=�>����=ɧ�>~.?�?�C>�����	8Ҿ�ᶾ��<�o6�<}v�<5O<�ޑ�������U���ܜ����2=�*> ��=��V<�>�xi=X.��u�������6�Ce��&~��M�=��>�[�>d�x>tR'>Y����O��οZ����t���6�$>~�ٽ�++�ŏ4�=zG�Ɯz>�f��Υ�>�?�;M�g�����<'D����K��A$>T�b��*�`D>��;�%�rɋ���]�h�s�j��א=b5����ͽ�o��W4I�+��az�S��N�w�bt8�e�m=4?!|�=��=$W?5w?}�>�=�q?K��p%>��>l ?�3>���=�P=ƴ>�w�=�L�vl�-k�V2l>��s��p5>��j>���<�>Z�Ř��d�=�!�3d>ӌ�<"F��p���߼e�<J�;�[Q>:�>j9<��~�������Ҿ�鈾�8��M8<K1Ծ�w
���J���������}����;�=s;���=w�E>�v>��F>����2,�����g5*��.	��A>�!��Q�=�>Џ�=t��=x��=�z����,aȽ;{��@�:\>�?��>�<?>�
�Ҿ}"������nh�em=�[�>�<>�Z>[CB�ٱ��]�Y0�� ��4����D����=��=�C=�p�>�:�=�0�=]8�����=�C���I��=�a1>L��>Z>JD>��=�䛽T +�ɒſ6֛�k���Ͼk+|>X��>�(��j��7��=)�=�QJ�;��>�`�U�
��n=½\��|t�<+���`=9x�Z�>΍R��۾����Y��#� ������<弾s���?~��3����3�z�@�������Y���ռ8>L�>���<ǐ7=��>ћ>��>��>(o�>_��<D7>ü��t>���>�[>~v>>+�=��;>�{�fR�@�k>D� >��S>(�:>��>�iǽ9>/>���=��=<)�<�^��X弐�O=��c>��>>Y�=
�$?��"��_���	�+��&ݽ�j���)?�J�=�r��-�O>������)�B�;��ݾ�>���>?m:�>��'>��q>�ϾlG��s 0�|����ҽ~�)>Q�>po�����\G�=LQ2�(�j�[$ �����W�U=>�Hc>P�S?wE?콏>���{sF�C�$�
|���:��E�>㳾�>���>/�>m�� Q��{7���#�J��.�ܾ7�=��S>аM>Ln�>�cz=h�A>89¾�Ᵹ��>ԏB�r��;G>���>}��>+'}>�Y�=�Q�����r�ǿf�����.�9ԧ��=�e�>0>/a��l���ڏc�{�ν{p�w9>Ӟ>�F={Ő=3���5X����=�b�>��:D>(�=aZݾ���j���z!y=���,i��(�ʒ�=A�ٽ�Y�G2�N3��5�}ՙ��94���;>{�>�з>\H%?�[W?5��>9M?�5���={Y>
|>Ã>M��>nM�>`��>���>��>ă��=�����і���n�=�/�=�d>ѣ>�9T>��=��j�Ϟ@��=>�.�F�|;@㊽fH��E
�=K��=�
>e�V>)�2?s�d��,M��w���,i��B��n���E?����Bn=w�?D���U�:Ig��W[�9�g�>�@=��?�-�>N�K>�0�>Hȭ�O�x���>I�⽈�ҽj�=��=�U1���ͽ��<�B\3��JW��S��v���>���^�= ��=J�>�PU?�(�> }�>�N�=�����L��C9�i!��sm>6ڀ�r�3>�b>�x	={`ʻt2���+�'s;������V��[=��>�M8>�� >��=U�<>L���L�D��>�a1<���`��>�Y�>R$?�p�>���=<���u궾@Կ"������h���5�O���%>�2>h���t���o���3��P�|�
	?=���>(˺=3FV�B�=Q^����=�0a>L�N�A��=��a>i����u������-'�(Β�F0>�/��3Ō��u�Oo�os��(����&��U,�"�w�K�=�A�>�:�>�,>��/?��?s�?�L���>���Ĵ�UN�>��>:~�>�
?�"?�;�>s�h<��`�z���VE�]e�<~����CQ����=˲�=��=��=��q��a�=�=L����żz[� \=�W�<�g�=�V>WiE?y吽 @�L��+ *����=F�����(?�X���f���]��P��G��<W��s� }>8??A?#1d>�Մ>���>�ǾG3潜V�=S�ٽ�@�<i=c��=\�	>g�T>��=������2�.��)��˝=�o6=�>�S?d��>�>�>�/��]�A����Л��;	>i�~<�R�>��>�>����O$�v�4��M?�͓��I*����=�0�>w�K>x�>V�>�KX<�5m�-���	(t>��]7=�>h)�>�0�>�A�>���=W�2��h���+ȿt`��&���<>e� d����`���Y={���;w�z��E������|y�g��<��>Ws�=���	�۽.}`>��-�HMv�gx=�~����ɾ��l��"��$3�=�%&�����z�!�ڽ���J��l2-�,5B���b�˅S��0����A=N�x>8��>���>$l?�|�>�3?/�'����>�=}>�[|;<�g>b� ?G?��>:��=��P<��7���=u!߽0N�&�=Gd<B�.����=��=Q�g=��=��G�$�>��*�ЕT<�C-�/o���5=6s�=�L>�>�E7?��/��F:���m�9�(|�;H����J>�4=���A�������|_�0��Uͽ��>���>π$?D*�>��s>��>+Ѿ�7��e�=e�*:l���D>�� >Qk4��k{�&�{<|�C�I�^���%���S�a=@��=�K�=�m>�=?R?�>%��>��Y���־/$&���]�x�Ǿ(�>Vb�>���>HSS>O #�R�ݾ8�6�J>5�\�5�\�Ѿө���g�=YW�>�`��"�i=Q�1=���=��	�9�,�'�>���=�G#>�g�>��>Z9J>5Z>1�1�yq�{��(�ſ������f�<�ݾ��C�-�޼fۼ�#�<�&<_xK�*ӥ�O�ؽԍ�=mc>�}>V'�=i���r F�+Ñ>�g�[~M�*唻j��<zx߾��C�����E���LI�BC=��'��νI��(���"��s:�ϐA�_)�쉽��W>~��>m?��?|	Y?�W�>]�S?�f��g^>��>Zf{>Xr�>>�?m?	�H>e�/=�^�>�#�=��^�����͐���>d )>��Q>�i>��L>L<�
7>.Z	�s =��5{�;��;k!�����=��>�4>"�>pN(?_>���wO��*F�^�
����^:?l2>�~�>���>u���_5�k;��������=O��>vZ?M>6и>(*��񠗾�	�=��׼ ��= ƽ����� >�Y,�H|D>2Ey���\����=���=LA :�}�;X	�S�>p�E?���>��|>l�&=\��`��>���� ��E�=D蔽�(�>�#<�\�[\<�5�	� ��f�O�#���n���H�8�>��)>�E>���Ǽ���=:E8=�[ʽ��(>y���	�>D�	?���<��;<0[=j��?0#��ݺ��ڗ��;��p��uq>���>��w>�!�)���M�����2�Ⱦ���>A��>��ݼ'�= ��=�]����4�4���ЦF�B^�=3��<G�� �׽�z���= �����Oc��¼r��I�E�?!�!s��2�u�нSJ���Q�>�7D>�{?7?�x,?�
?V �>@�
����>�<=VZE=�	C>���>:�?��?6�?k��>�Q������S��Z"���*>zJ>�5>B�e>�>�3=�� >쩢���=r�&�*Ղ���̼ş<�^�=z�=���=��O>�*?�+�;gv��)s���y��;�վN�������>��d�Ծ@c��H���0>x��>n��>���>\�=$[�>~)A>��>>C��.>z�=�-r��~�=��Q�� ��eǽb�~�d�=1�,�j�v=m�g;�3�<F�X=Z7b��|�=�B>f�M?�e�>\�8?����B,�U4��Q������J>�"�>���>����|�c��I ;�-5�t��^V���.��݀>fH>������=;L>�b?����h>-߰=�V�>�~�>"t�>.��=�,�<L? �޹�P�%=Ƚ���������=����vA`�(��>�K���?�dU<c>�d�ֶ;���1��!V��-�X ��R�(>�S�=-g��1�=K�*��Y{>�x��2���ܥp�K/���
>���|��x�齑�S������˽�n��B�:�ny�r�k�o�a>��>���=�L�<z]A?
�?�?d�۽�y�>u��>�>�>|�?E6�>a�c>��>�� =�MT<Ű�>�d�<�}H�Zо�$>mo�=x�;>�`�=���>�y>S|>���<�u2��
���8�<��|����=s�=�g.>�0�=�3C>�A�>�ZY�*pž��m��"*��n{�5+�����,�%����c��-9���]�O��>�>�[?TM�>H�a�<��֝>��>{Ҿ�=Nx&=��þ.�	>��a���<��Zn���=�H�=��=��X���4���M>��=60�=��>ٲ8?3Z�>��)?^�<�I�-���þ��Ӿ[������>��>=X�>��>��5��I�C�A��g�������Ͼ�׉�w�e>�u9�����U	>���>b���W�2Д> P�=�.>�L�=�/�>�\1>$�=�"=Ia�:��awB�-l翁a��*��>��.�}�2=]9�>�݅�	��>��ƾ&O�>�L��~�,��;Ͻ�f����8��h=`H���=��e�k�g�%�ӾL��>��ٽm��>�����:>>묾;��<�u�d[�����R����1���(�x봾�g��<C��c�>�~�>E+��?�K=���>IJ>�$?0�N>k*?�я=�->�j�>z�?|	?�^�;R ҽ���<S�G>-��>��y�h�#>(�=�W���\�<�>O�=:�8��d�$�=�9�M��F��<H}n=�H�<_�>���=o=�*?�+�;gv��)s���y��;�վN�������>��d�Ծ@c��H���0>x��>n��>���>\�=$[�>~)A>��>>C��.>z�=�-r��~�=��Q�� ��eǽb�~�d�=1�,�j�v=m�g;�3�<F�X=Z7b��|�=�B>f�M?�e�>\�8?����B,�U4��Q������J>�"�>���>����|�c��I ;�-5�t��^V���.��݀>fH>������=;L>�b?����h>-߰=�V�>�~�>"t�>.��=�,�<L? �޹�P�%=Ƚ���������=����vA`�(��>�K���?�dU<c>�d�ֶ;���1��!V��-�X ��R�(>�S�=-g��1�=K�*��Y{>�x��2���ܥp�K/���
>���|��x�齑�S������˽�n��B�:�ny�r�k�o�a>��>���=�L�<z]A?
�?�?d�۽�y�>u��>�>�>|�?E6�>a�c>��>�� =�MT<Ű�>�d�<�}H�Zо�$>mo�=x�;>�`�=���>�y>S|>���<�u2��
���8�<��|����=s�=�g.>�0�=�3C>�C)?ٷ>�C?�ѠH��(ƾ�"��X��w��S���s�>����oS>�V�>z?��/>T<�=�;~<,�q>� �>�ݬ�����#�<�g���=D�4��.��RȽ��|��|4>8�H���b�e㓼�Ae<Lx�=Ge= ��=w>�Q=?|�>Ъ ?痘=��QO��\��a-�N>r�>���>4�}�E��U%��:4�M�,�|�Q�xD�����#qX>��4=W60�S�,>��^>��n��=���>Kf޼�>f�=p��>
�3>Ռ?:��-��R�ÈٽV���aϿ8����\�Y�;�B�V����=6��B�>�>M�
�p>�{������M=�����h���H˼/A�>��g>��w2��4�>>ҕ�����p=?v��HCP<zȸ�]�=\$��k��c����Uؽ�2e���(����J���`>߮�>]и>���>/Yc?>�%?A�A?F'�>��J?�Ս�?�>i'?�4�>�@%��������U�>"�)>{ S>�ͽ�����>A'>�������&K>f��=%cF=p!"=������<#�;�<	��=cz>��@=H��=��>�A�>�ZY�*pž��m��"*��n{�5+�����,�%����c��-9���]�O��>�>�[?TM�>H�a�<��֝>��>{Ҿ�=Nx&=��þ.�	>��a���<��Zn���=�H�=��=��X���4���M>��=60�=��>ٲ8?3Z�>��)?^�<�I�-���þ��Ӿ[������>��>=X�>��>��5��I�C�A��g�������Ͼ�׉�w�e>�u9�����U	>���>b���W�2Д> P�=�.>�L�=�/�>�\1>$�=�"=Ia�:��awB�-l翁a��*��>��.�}�2=]9�>�݅�	��>��ƾ&O�>�L��~�,��;Ͻ�f����8��h=`H���=��e�k�g�%�ӾL��>��ٽm��>�����:>>묾;��<�u�d[�����R����1���(�x봾�g��<C��c�>�~�>E+��?�K=���>IJ>�$?0�N>k*?�я=�->�j�>z�?|	?�^�;R ҽ���<S�G>-��>��y�h�#>(�=�W���\�<�>O�=:�8��d�$�=�9�M��F��<H}n=�H�<_�>���=o=a�?������D��_�4�^���g�=�`�>�aS>�>o����	��� �>��� �Ƃ�>��>J��>��=3�u>0ZF>�iþ�����G�>�%*�ݺ�O�s=�Ľ)t�;��=��L=S��-/�˾��l�9�w��=� d>�_>�g�>�"%?�|�>*,_>*&>m�~�.�C��Z9��㗾��@�}�o��%�>���=�7�=2(��y�$���ݔ �.���_���t�>��L>$O=��7>i�=2����� 3>��=���<㙃=�^�>#ɓ>
nd>�>=������o�gb�fuѿ�ݠ����<t'�=jc�Ǡ�>���6�������\��/�w<D����>Gr(>~��>�W�=�A���>z>�"�>��j�)��>4Q�>�j �掉=8)��S�=�F��+⇽8�N��zk�jn���^��D��N2��"F�������i���N?EA�>�	>��]?��?n4?"�8�2��>����>-6�>�9�>Z9�>�v�>�t>��}= b����
>�'��a3¾h�<�!b�����ἡ�n>50	��𼂟U��{<��K=Ђ�=�o��c�5=� ��=�A�=o�a>�-?���l����������%	#���E>���>�j����>�A��3ľ����)�%���d>���>D�>��>Pڅ>�Ћ>Y����d����>{���:����P�=L�=(Z'<t�Ѽ9��=%�=�ۮ=$����$��w��<^��=^++=:%>΂?�-(?C�?%[�]��HP���&���g�c8���[����>C|�>yV>R6�������;��M����fr7=7+�>��>3�G>���=�T��_����1����������Y<���E�1=&>q�E>�tt>g.>�	�,z���dӿ���,X��k�d��O!��V>�4�vW��/~�����w}�=�D=�)`>�v�>��>�����]2�g5|�����u3n����� =�_T=u��ڭ)����*y�ӛ��yn;m��N��x���_9�V��#_��r�!L ��Wƽj�=J�?�/z>펗=�}A?���>;r�>��k>��>EXG��?�=	'>��>Z��>4Y?�>^X>_�=����B.��^���v�=��=�f�>�[�>1�<�gZ:�F�Zx�=���<r�ǼbS���Ы��7Լ�I�;.Lh=ӹ>>�&?������QE\��b�+㜾s#���I�>B<�{��~�Qӳ�e���ƿ���i�nE`��m>BS�>�>�>��>��>�6��멽|�'>�]A=To%�J�;>J�>#w��o�9P�<�\���=.������_6�<'>�=@꼷�&>�l?=EI?�4?�gm�����-�������
�����b���4�m�>���<O<A��	�����?$�(�Bv�<�X�>�S>�/>�o,>钻��\�|��u��c�j>�����-T>���<Q�=n�h>�}�="�����������ſq��5�x� �޾ⶴ��H$�b�콇s�@n���L�>��>���>ٱ�>�ԛ>gk�>!6 >�+ļߡҽO����y��p���ϲ�6��E��)���&*��}½Lc��/�E��]��\��A�q�a*���	=%["��Or�H��t<�=��,?���>�@�ȿX?��?)?�˩>6?�>w3L<�$	>F�Z>�>�>J*->�5?Ԍ�=ղ8=���=Nia>h�5������`9>$���T:����>�<�:�Jؽ�>=jZ>�� =��N=#����"*���G�=k��=��1>a96?4�<56@�mr����"���0M���?��>�<������= �5=3ƌ�J�����������=wD>:L�=�jQ>��>o����%���)�>��8��l�<a�>�P6�n��=���+�f=M.�.�=]��<ް=I�=,��=�~��8&>4A�>y ;?�.?�������?�lʾ��w=oux=�	U=�M\���>�pt��%o��9��'���	Ҿݕq�q�=�F�<��:>���<˔��n�=o�D���=Q{>Z2u����=ή�>�)>~��>f��>�1^=���ur�պk��]ſ%➿�7�>i�.�q>��g>w?/������{�Dؕ>:л��cE�� �a��<�_�>㵶>�N=��<� �=:�i��v��=3Q�<�^��"������[�м��ǵ�����I�~�ηýCG�NX��
�;�l��!��Ƚw9�=H?&A�>M.t:l�?:�?Ċ
?B{ݼ��4>$޻.����>�V�>C#�>d2?;��>��>�*>2�7�Q��𕾺��>�}�>���=M`n>�Z->�&�:�ս���=��&>���b����:�v���.��,>��=�n>M:?ώ��l����	�=*�/�R�N����>�켽��$=�%\<hݾ-����%�M-�&�=`��=r��>�)>Қ'>�N�>�����{��P�>�����8�;��>��;�0=�̗��_�=(j��e}�=�_g= �)=��-=��%=���<1�B>��
?�JP?�?�O1���]�B�>������Az��+�={�=��/=�2�>�׾���)�	����n4><3L>?�>r}>�	�=YF������͞<xAt=�{��wb�=�g�,Hc=��>[��=io=yNb=��E�z��98Ϳ���R������F<�Q>��D>��־e�P>��m�^�#p=���>�)>.V-��h>�Q��=ѝ=�2!�m���	���B>8k�=����B=Z��bm���F��A���)�?>�I��5��ky,��? ���K���%��M���r��G�#?R=V>��R�0�J?��?. ?N�=ֆ>�EL>>�>>{�>���=ۯ�>�YC?2��=�{�=oJ�����==�^��&����=vv�<)>����=3�?>�A��#�=]V�<�E�=�!��z٥=�cĽ�Jw��(���&�<\w>�>4*5?JAo�ϫپ��-�0&ԽZO=J���I�>\���ɾHA6��%轏�=�~�>c#v=
٭>e�>�}>`J�b�A>�\>#����=�?=�<��s�=�N&�Բ�Z&@���"��bܽ�|ۼ�x���I<���-�<e\>�s\=@��=%�l?�$N?�A?4ܾ �n��SҾ�8$�Ā���S���4[��n"�L@<�LY�ay0���L��C���T>�OQ����;�E.>�y��+�=���U6�~��=Q�r>J�q>8Y�=b�P>}�t>�qs>��!>���=G�5�ܾ�^��5˿�#��-m�r.h�O�}��έN���t��Z ?$?^j>��@<{C9��+n�*��>Ӭ����ܛ�>����=� =�\�=
r���*޾V��'-��\ƽ�v꽑L���9�����/,��h��.)%��񽾢*;���v[=���>�h�>{�>�pF?� 0>z�9?|�3>�|�>�A=�z�>�P�>�<r>ZKM> 4�=L�h>��=O,��Z ��$+��<���g���h�99V>^{F>Qg�>��=�/�<�L�<���=�4=9^��qS�*��;!�=�h�=Ϝ>x�>=�?���<��&�϶����V�2U-��S	>)�F���>>=Y;>7vI=�Xݽ�ȃ����=\n*>X�6�d+⻹jM>HU�=�(��np���ٻ$}=��"=NK6=~�>��=����ȣ�1�:>C��=A]����Y'=]>=�9<�O�>Du)?b�U?t�>�Y��L£������ �A	����>l;>^�������?��̾����	�k����K�=�1���ܡ�6g>�Z�~�"<�Խ�%Nc�C�=���=�_�=1��=Q>��=��>>n�B>5��=&`'<�c�����C¿����b��.��<���=�/����=�U�>tG�>�d��k�>��=�.�=�bD�~m�=2�P��>p�p�ͽ5Q<>tV�*[�*�ǽ?�	=4;�FA*��X�|��f ���	�ܽ�r�e�[~ؽc�<@G�<�4�0νۃ"��,�>ZE�>(�<>�>� ?g?Qh?鉓��Q���B��gq<bNW���<VJ?��?ِ>r"�>Ԍ�>�ֽYom��ʾ<(-6>�֘>p->kF>�z�>�Xp�.X�(⽧r�=���|��F]����</��=�_�=L�y>PB>���>���LXǾ~���/=T�{>@t�˘b>4V���6��⛾��̼�c<���=*�0>l/>�V>h�><����=u��=,-��I��Ze>D/h=�؏�p�@���)>8��Vʽ� ����p�ؼ�C�>q}|>؅>"9=�ņ>�)=�??m�C?�l?� �P�������n	�yO<�c_>W	4=23�������"x� k;�{���o�\>Fv&�/�$�W=���U�='ȥ=�ґ���Z>z>ح=�G>z�S>�G�>��>�|5=��\�}�v�5�m�+�m��޿�觿ߦ����Q>h���=�)$�>aN�>����r�>�>/����~�G<>�=��8>�؈�aG����6=m��>��8=�b�>�'>�����O�LB�pF��)�ƾ������>������U��a%��c���h���ŽI�2�� �с�>I�U>��.�����Dy�>�v�>�VS>���;��=</�t5D>��2>H�>4�J>��>�?�><3�>cc�> ;4��;��ǘ/��#>S��=��<�7v�2��>��l>3؞�b��<.=�<g�=4�ջݟk�Jv���T���p�=Z�:>�'3��?��׾^��*�޾�L�Z ���#滩Ok>*V��F�<�!�=�	>]c�=J��i`���>쮘>�p�=4s����f>�V>�󈾝��<TS�=%A;>�K<>��<v�8>a�T	�;:����e=!�;�Dt�iO�B��=-�7<�=�����\?�[?DI(?�����*����V?�>�X�����=����4����Z�j⾲�9��g9��)�.˼D`��p;��=�N��f�{>꤅�Pst=�g7=Na����=V��=��U>Vz>5�L>^�,>���=�3
����&o��ؿS�s�C~o�0S����$���!T����p<�������j�5�+�-b��~*�E@�(��N����;bU�=&�=~n
��=Ivt�_]�� 
���>��e���|=PӠ�����=�Ç=��=x��:D���,
>;��oǩ>Nq�=4�_��k�#�?A~�>;�>m
�=��>��`=�������+>t��>��>+�><�>bՍ>��3=���+�=�n�=��=��5�=��;�(�;V	�3�<x;yH?=�`ܽ�ë������=.�?=���<�*>��C>��?DM�d�t��6y���(� ��}��ِ>����0�J����K=K>P��=�zz=Qօ>{��>�^>nx0��Ks>�a=��<���ͼ���=�:���=We�=d�[>Q!%�z�-�����fq<�쯽
�Q=���=FQ�=�t'>�?��^"<x�`?�s?kdA?���>��71���F��>�ѷ>.�6>��ý��c��>�o� �(9��Z����K�>5<f;�L�`C#>}	6���=�9=��%N>-�*<��%>S�9>��>m�>���> ��=��;�gh��LA%�����<�ؿ�͋��F��þ�h:>(�l�@=�jI>��=�b�0>�>�='�s����N�=�]I>g*K��0���=�6���w�I�s�K����?=]�w�Y�h���q�^Y2�&��d	�9޽�Jr��F��Q���鶽���7+����&o���?a >��t��X�l3?4#$?'$?��_>�B�>�4����I�=>�x�>���>���>"p�>@��>��9>�������u=Ԧ�=��5>����=6A�=<B"�/�<����ʾ�I񍾐�v.Ľ���_=���=��A>}��>b$�>��νM¾������"��!���H��r��>�ls�b�n>�7���/���-ܾ���.��Su6>�߈>�3�>0q>�]q>O'�>��R솾��K=}�#�+��=� ]>��>�h7�<��>�Y�=�ի<jB�=�~
>#�\<����0�=���=;�">pPE?��>hl�>�B�=�L�gް�胖�����t�>�Y�>���>hf�>FY�<�嗾�D�Q�-� ��g�����{,��Tٰ>��>=>�4+=K6-�1�'����=V���9ؕ�=Uk =���=S+Y>�F�=#�Z='e��[��7�㿷c��xB|=��"�f=�>f"�>@��;�TϾ�B��\1�E�u��V=��>>�Y>-�H�ՙ��f�� #��{���]>� ���-y=C�=���I�����۾j<���D��������3J�M�������A�|��l���銽R�[��q>\g�>HZ(>��i> � ?J�>~�?_�=ܔ�>XV��5 =��=�o=>���>���> Tj>��'>BA<�3�=�������JB
>��+>�>	�1>�$@>��꽨��<��=<c���E��>ړ�<�`��ы�p��=���=4Qk>%�?��>�9��qx��o�M��}�������>)���t�<,�������V{�%y����>��p>��>Q��;�f�>(Y�>N^��% �$遽zmh� #�=�"j>�ҽ����g0�=�_7��QC<�:�=���L����ʽ_�~��7
=YW.?@%,?dr'?��=���
�������[�E�-������ ><��=
����2���_�z�$�@A0�[�r�\�ן�<��>���>d>�T>�	���@�[�>,��>
v�>�l�=��I>��>eN��W�=@m
>	��=�O����Կ��#P��'�$�us�=RU�=���M�ܾ = >��P����=Dm=��F=�7>��=��8>��3=�S>}���ghʾQZŽGJ\��w��������[!�+״��m��}��u���ǒ5�(��ꗂ��� ���	���=�ѱ꽳*>�>L��>���J8=?T�?-�?���\�<?$�>�q�>�e�>E1?��,?�d�>�&�=��V��(�X`�>�u��V�W���u=V��3'�=<HR>`3>7oN�O�>���=�R<u~=�hռ��`=�\<=#��=���=7|�=Fs�=�(?cڽ\9޾�{f�/�o ¼��վ�{>J�i��>�N��R�� ��a����H�=�U�>
�>_�>��/>S�>B��>�䡾�Ƅ���=amS��3�m��=��^��+�4�G�m�<q�=���=���<���S��x�<���=��>�
R?���>��>� �<�C���z��`���,�R
���'=>�Rj>M�Z>*V׽��}�Bg�7P��W�Z	����=��>�խ>e�'>YF�<2٣=/�̽�g�>����!?>����00=F����@=��;B5>�D�WÉ�%�ܿ㬿~3���ؘ��Qm=fu>L��=�f��/6��MHֽ��N�(0=߶D>m��=V��E��;���;/R:=�; �B��+=��W��I��Jǿ���;?ת�MN�� iE=�UJ��-����;�����8�����9r���H<�{؞��{>ħ�>�
>�+>? �N>/�?I�_:�1?H��L��>�>���>�8�=�VA=��2�KO=pH	��g->��<��ƾ#=��o=+��=d�7>]o>�U��^K>'ŷ=jhI��D=����l,�9ݒ��ڎ=).>�;�={�)>qS�>�y�M���߈�8��ו׽ϞV�;���|H��[��ྭ���Ŵ7<f-�=��m>��>L�<o��>	��>���>�w>v����T/�ɹ��½���4�<��C>�F�<[+��J�=�Z>���=(\���;r�y*ͽO�߽Y3x>�h���3>��?��?��?4�I=N������¤�qjn���.=���>�%L>���<�=�~t¾fﾲ1���~ﾮٌ�Om�a<>.9�>�>8+>K��=\�Ľ��I��$�AF�>��='�F���.�qE8>�j;>@I�>=0�=%��5���H��F���k�����׾�`�S�0<Y�<�VR���*��=�@=�=�U>;�D�=�qk=�1�;��&=?���ٹ;>���$�*寽C,������T�����ԑ��\�⃽r���P���\0��w�p>��V��T�<�p�&��q������?d){>�] >��=?���>M,�>®>�?RqY>4�>��?>�r��6��ҽ?��=�u�>�pM�^ǃ�R��w�Ͻ}�+>�!>���=;:=>v� >�C��Ɛ(>i������O��&uo���<����Z���>��=��8>�O?�9�����ԃ����d�������JW=��{����9E ��*ýF>�|�>���>�q�=[�W>lP�>B��>�Ś>��3>9᪾�k���^F���M�	m>ئ�=gk���ѹ=z=��t�}<d��E���e�X��=J�=A��=s��=sS/=��!?fP?P&?#��=�ʢ�V-����c�K������\>��=@�ν��� $����!
�����E���
���=�x�>�^�=�(>�+�>��/��aۻjHE>l��<K�ڼ6�=.#6>��#>[	�=�,����h�J�"<Ľ9�׿�;��8��G-+��>����J�=�G���6�=�8>�H7>��=H�{�� ɽ|�;��w>q7'>/ս=�Q���Ծ�,��E��=_i������R�V���e��Ͻ=iq��۽��g��'��I�$������r ߽�$�6�=�#�_�u��=uQ ?���>1��>`�#?M�>_�>p5�>i��>���=h��>O"�;�����ӽ5���]&�=������Z��z���$6��E1>�*>"��=i�>ve�<w_���>B~��D��=�4�=�g-=W��=	�J=��&�a==疾=�,�=Һ�=�Bk�7���6������� �>�
�r"\>�#Ӿ����n��Xؾt��B�+�U�n�6<�~>e�>c�?Ne>��W�agP<x��! ���= D�;�-ʽ�x�=��'�����C1ھ�]���1��6Ͼ�y�L�k=dB=s�N?�NY?$��>tRt�C�>��EZ���2��X�F`(�sz�-w0�')f>3ؾ_�3�2�O��'C���S��w$��x�<*RH=A�o��=�F�>��Q>(��=	�8>뉖>�G�;ݍ>�>��>��j>>|>p{�>b��>��>L.־,�ۿ0������!���鷽�N>8�Z>Ap�tj��{���6����;Df��)&+>�w�>:�3>n[\=�I�=�g>v\�.��P��=۸���<�\���6�����6�>�����"��ｌ�ؽLέ�T�M=M�A�V��k��=��?g�q=ޯS��v>�??�2?K*�>�*�>[X�>�O�3�?�k�>���=��>�U�>8��>Q ?*5?��>�/�;�ͽ����r��}�<��5>��,>��սNN��q=���<�2>:�����M�=�pQ=�=�
=`_=R7P>a��>��=>�:��o��D� ���J^�=�0>�s���:=�����Y,��_ƾ�"
�￤��>��<�ޱ:�->�ݺ>3��>��=�H���ն�9.��GI�;V'=���`�=�U�>@%8������<�@����� ���!=��ns<v%?
??��7?L,(?���<u�5��zT�4�&�*G�<���<��?���>�l�>�D���!��C0�o�*�����ݣ�����&Z�S��]��=��>p z>7j>��=���=�%��^hݼ�r=0�>��">�UE>��P>�#>�{=�*�����h���4 ���5�<�=��U>��
>�t�=>��g�e�z�l��Ճ�Bm���i>��>�v>u�=�3X>;�>�*��و���ٽI�-�Ǔ���D���!�>��<9ϭ�(�=k������������t�@a�!���G���<�j����<����.>��/=%��>Y/?��>�m�><r~><�=�f������!�=���>�Y�>9g>���>w>������d������=w�=���;��=��}<�Q�+�0=ƾE�H�ս�S>���`�j��>�k�=}6�< �>����X���:�1XR��9j��"����>u�?�eվ��.��zɾ^[M>u�;=Y;N>.?��V�k��`��>�"�>N�>n��>�g>u��=��m�:����`��D������7�w=��=H�@>'@�<�8��7~��p��*),�� � Cj>�*�\�"?�Z_?r&?�S��Hk��2��C�R�OU�E)=n�-?�؂>�E=����k&��p'��7W�3f����D��6}��f%>I�=o�6=%,�>��=ŲL<A�c>á�>�>H�-=�}�<"�=���=9X�>l	�>��>����������╿��Ѿ|C�C����<7�\=�����н2E���@�����y; �=t�=��=�=�g�=H�=sE�,탾kFg������}������ic��=ǭS��p�6���A��K�4´���=��Et�툾�����,"��?�>ލy�V~&>x}?u%?�_�>� >>�>��> ��\T��l{���)>��>į
?�?L֟>��C>&�Q��/�wFŽgJ����=w�q=4��=�=x�˽��I�c+�	pR�������<oڃ=} ;�'����=+E�=�)�> �3�Ā#���=0*�졌��=�$>�N���Yw>�:������������(遾�"�=�0=G>��=��>�9�>�+D=����}4=V
�i�
���<�!p=֐G��C�>���<��ɾd������v����U��ɽ��
?sV�>�^?
$A?b�>l����P�>E]�h9��ё��Y�/?>aV�>�n>�c���Q,���\��Q�99[�JM̾O�<ī�=6���J1���=Dh>>�f>�i>AcH>Nu�?%��б=�~�>�j>$2�>Q��>��!>@��=���^���
��Gn�����c��X�>�i3>���=SI�9f���Ⱦ=G�U򧽍�{>�Lu>x��>��>6"�>��>ȝ����<�f8D=>�<.4��B�\�s�>��8r���(�Xi=A��CfB�^���ս�	N��˽e�꽛8�s�����>��>ڼ,:=�V?q0?��?�n�>Fj�>���=��>�UӼ�K�=�=�>T�?
@�>��>���>�a��E��l�4F-=��=��=(0�>o�>�9L�Ľnf�=n�:R)>���=�:U<�5X��%a<�=B�q���=�)�> �3�Ā#���=0*�졌��=�$>�N���Yw>�:������������(遾�"�=�0=G>��=��>�9�>�+D=����}4=V
�i�
���<�!p=֐G��C�>���<��ɾd������v����U��ɽ��
?sV�>�^?
$A?b�>l����P�>E]�h9��ё��Y�/?>aV�>�n>�c���Q,���\��Q�99[�JM̾O�<ī�=6���J1���=Dh>>�f>�i>AcH>Nu�?%��б=�~�>�j>$2�>Q��>��!>@��=���^���
��Gn�����c��X�>�i3>���=SI�9f���Ⱦ=G�U򧽍�{>�Lu>x��>��>6"�>��>ȝ����<�f8D=>�<.4��B�\�s�>��8r���(�Xi=A��CfB�^���ս�	N��˽e�꽛8�s�����>��>ڼ,:=�V?q0?��?�n�>Fj�>���=��>�UӼ�K�=�=�>T�?
@�>��>���>�a��E��l�4F-=��=��=(0�>o�>�9L�Ľnf�=n�:R)>���=�:U<�5X��%a<�=B�q���=y�Ľ�|��U7������8�C	Ӿ�t��!�>��!�>D]>y���|�Ӿ�H�׾�G���뮾����
>�|�>���>H�;�F7����r��-��T�>�OF��΅>��˽�+F>����ߔ��u�����<-"��e��'��>t�[���Q?��H?�">yG���5f��}�0�i��?�=p�q>S�R>@k�>xC"��<��J���X��L��\���u�S��<�Pq>ؾ0�_�>�>m�=���=7 콉H>/�d��&R���V��QM>(L�=�=�>S>�8S>����3�
�vM���@���c��n��V�
��=a,O���˽���c���!�����2�e>�o\>�(>T��>s�;<����<�=�h9��	�l����{x�[�"����
�ξ�1=�����=z� �x-�����|��PV������Ӿ�
�9܎�w�?������E�>�Z?��?��?]-�>#L�=l�%�1�@̸=HE>]F�>�K?}�>�?�+�>��9��'=#D'��v�<X]�=�
�=�4�=�>Z$
��[}<'ZP���J>L�[�=��$>+y�=^��=v��=�r�=��>���>�C�d�0>k�o�	$�OC��pQ����>��>����F��E%ǽ��ھ�O��%�8����<)6��U>��f>���>�/�><m���н9�������V�E>=�R=��b��<l=k7���kH�8%� !�C㽫�?�����g�>��>&�@?r?�>?Cc���r/����[Q��饾���P۩�wL�>�g�3�9���B���r�|ks�wry��f��^5<��>K���'0���>��_��;>4,>��.>��O�-%!>l�}>>/�>I|�>ʍ�>��`>4���Q���ҿ�咿�]�y�I�{��k܀��/�=%p:�H�=sC>
�������<���|�>3�>/u�=K?E>���> A�>i]z���Ǿ| z>����M�����*��`�)�������=��ɽ�� ���`� H������
�V�@�"��=Xe�+m?�f]>�x+�� >��G?r�Y?��<?0��>���=Jtt����>V�3> }?	?v��>;�?g�"?�[�>@g�>�����O� j%<�b&>���=]͕=$�=*�L��ڹ�F�>���=g(ν�Z�ژ�=�=W����P=����Ǽy�Ľ�|��U7������8�C	Ӿ�t��!�>��!�>D]>y���|�Ӿ�H�׾�G���뮾����
>�|�>���>H�;�F7����r��-��T�>�OF��΅>��˽�+F>����ߔ��u�����<-"��e��'��>t�[���Q?��H?�">yG���5f��}�0�i��?�=p�q>S�R>@k�>xC"��<��J���X��L��\���u�S��<�Pq>ؾ0�_�>�>m�=���=7 콉H>/�d��&R���V��QM>(L�=�=�>S>�8S>����3�
�vM���@���c��n��V�
��=a,O���˽���c���!�����2�e>�o\>�(>T��>s�;<����<�=�h9��	�l����{x�[�"����
�ξ�1=�����=z� �x-�����|��PV������Ӿ�
�9܎�w�?������E�>�Z?��?��?]-�>#L�=l�%�1�@̸=HE>]F�>�K?}�>�?�+�>��9��'=#D'��v�<X]�=�
�=�4�=�>Z$
��[}<'ZP���J>L�[�=��$>+y�=^��=v��=�r�=��>���>�C�d�0>k�o�	$�OC��pQ����>��>����F��E%ǽ��ھ�O��%�8����<)6��U>��f>���>�/�><m���н9�������V�E>=�R=��b��<l=k7���kH�8%� !�C㽫�?�����g�>��>&�@?r?�>?Cc���r/����[Q��饾���P۩�wL�>�g�3�9���B���r�|ks�wry��f��^5<��>K���'0���>��_��;>4,>��.>��O�-%!>l�}>>/�>I|�>ʍ�>��`>4���Q���ҿ�咿�]�y�I�{��k܀��/�=%p:�H�=sC>
�������<���|�>3�>/u�=K?E>���> A�>i]z���Ǿ| z>����M�����*��`�)�������=��ɽ�� ���`� H������
�V�@�"��=Xe�+m?�f]>�x+�� >��G?r�Y?��<?0��>���=Jtt����>V�3> }?	?v��>;�?g�"?�[�>@g�>�����O� j%<�b&>���=]͕=$�=*�L��ڹ�F�>���=g(ν�Z�ژ�=�=W����P=����Ǽ���>�C�d�0>k�o�	$�OC��pQ����>��>����F��E%ǽ��ھ�O��%�8����<)6��U>��f>���>�/�><m���н9�������V�E>=�R=��b��<l=k7���kH�8%� !�C㽫�?�����g�>��>&�@?r?�>?Cc���r/����[Q��饾���P۩�wL�>�g�3�9���B���r�|ks�wry��f��^5<��>K���'0���>��_��;>4,>��.>��O�-%!>l�}>>/�>I|�>ʍ�>��`>4���Q���ҿ�咿�]�y�I�{��k܀��/�=%p:�H�=sC>
�������<���|�>3�>/u�=K?E>���> A�>i]z���Ǿ| z>����M�����*��`�)�������=��ɽ�� ���`� H������
�V�@�"��=Xe�+m?�f]>�x+�� >��G?r�Y?��<?0��>���=Jtt����>V�3> }?	?v��>;�?g�"?�[�>@g�>�����O� j%<�b&>���=]͕=$�=*�L��ڹ�F�>���=g(ν�Z�ژ�=�=W����P=����Ǽ�(A?]쉼ymU���R�W�>���0U��-�>��q>��>���C�n>����3�������>��?�L>�w>#6�sc�=9�ȼO1]��j��
~#���>��*ǽ��->a�D>�#�=��|����=�\���>f���O>��>��]?���>�ę>��=�;0�������Ձ�*���9mB��K4>gQ>��5�뾝���H��T�s4����ny>�>=��罦V>ޗ�<+�	>�"�='>3�>)8:��Y��7�=LAW>l��>��>)H��so�=R|Ѿ��ֿ���k�;��)�� ��<���=T��=����T�2:M��cR�r���K,����>��?���>�(�<�ŭ�
����{Ľ�|�����=.:��+���a:YS��Kb��1����E�;Az$��<�������<(&l�8�Ď��QGE��L��>$��=D��>��j>(4)?:&?w[?�5J>��V>T`⽊��>��߽�?,��>H?�7,?��?D�>D���`\����=��Wy<(C4;�z�=�-
>�I=Kٰ=XǙ=�QO��*����4�e'=�}=~Ю=L��=��@=b�;>Y�#?��;��8��>���x�_�>Z9=P�?2��=�e=ܴA�rv���!	��* �Oj���ܾ������>v$?��F>��=%�B����\[��ѝ:��j>����>6;��i��V��&=���<lv���j�U��|$�i�=�ph>`U�'? 	�>�\">]�=�����=&�۽���F���kܽk>\�>�pl��a��O���X�Ǿ�z	�ԏʾ��nh�>t���|���G>����S����O�=w�J>�k ��>Q�v���ν�V�=�>5��=��>Z:	����qxٿ�ʵ�x�Q����"��zj�=̓=,5���.�웑=�
�df=�|;NA>I��>�M�>X�C>��H����k��B����=_�1�׾�ف����r"�S���T�(>����ж�$�>Dj�^e�~���y�eu�ɿ<�Ҹ�=��=K��>)e�>�?)�>�O�>��	�$��>BՒ�5��>����E�>+?x!?�?�#?y{�=�s^��P�����P<>ِ=D��="�>��=�_<=�C�=��&>��r<0eD��c��b�d=�˃>��?>>]>�(A?]쉼ymU���R�W�>���0U��-�>��q>��>���C�n>����3�������>��?�L>�w>#6�sc�=9�ȼO1]��j��
~#���>��*ǽ��->a�D>�#�=��|����=�\���>f���O>��>��]?���>�ę>��=�;0�������Ձ�*���9mB��K4>gQ>��5�뾝���H��T�s4����ny>�>=��罦V>ޗ�<+�	>�"�='>3�>)8:��Y��7�=LAW>l��>��>)H��so�=R|Ѿ��ֿ���k�;��)�� ��<���=T��=����T�2:M��cR�r���K,����>��?���>�(�<�ŭ�
����{Ľ�|�����=.:��+���a:YS��Kb��1����E�;Az$��<�������<(&l�8�Ď��QGE��L��>$��=D��>��j>(4)?:&?w[?�5J>��V>T`⽊��>��߽�?,��>H?�7,?��?D�>D���`\����=��Wy<(C4;�z�=�-
>�I=Kٰ=XǙ=�QO��*����4�e'=�}=~Ю=L��=��@=b�;>��3?�A�G�;�5�˽f��2��b`����>��>T4>��`>�춽RվT:�5��L���)ټ=hx	?�#1?/�>+©>ƫ�2�̼��,=qJ%�C�L>�F$�z0�����M<�V�>0�O>�*.�����1�������w�=�$
>�8>KJA?�=4>==c>ԩ�=���}�*F�e��6�˺c����Ư=��%��ʼ{��B �pi�<��2�.��_�T�>>�>6�=u�v=&e���ܽx`>>� s=%�>G�=B���ʐ=���>��n>��=�C>A1���ۗ���п�"�������D��< ��lm=/�R�ܤv>6��Ȟ� ��m ���\>k<�>U��>6{�=�����m1�(#9=�D��É��Ӻ��c���A���: =�.��jӵ<�b�`Ƴ�3A��졽4��B�#���OJ�95X�(*���X�E$d>�MW>��$?+M�>�/?�� ?զ:?�j=f� >�R��n�>).@>�>I�>w*?�5G?"�?��W>��<ji-�l}��J&�u��a�彽=ٳ�=nTx��x�=�L8�r1�=�=�,�=�k�;���=i}�=ntC��_�=��&>δ??�����&�P�`3=�4
x��>�'?";c>G�W=��T>@
���D�q�(���߾���>.?e8?���>�1y>t%�>��]�����>��G�a=�_m����<���=��;4�q>�bO��4Z���H�k�6��Az=�Am>��=G���?��`>T֦>�C=���p� ��I��;��s�ν|������>IH>��D��˾]4������k����՛�2Q�=z�P=^=�k��HM=��=�%>"�/>�g<�*f��&9���=��t=��>F�/�a�b���'�(9 �nlϿ ح���˽�k����̽�8>�q�=i��2���_�>K�����W��=��>�&>���=��꽻C+��P2<5�޾a���q�h>�r=���-���T�������j��"c�ʉ=��q��1 �W�վ�kϽ0l��b���_���_o�<r��>��?��>	>D?�7?��><>��2>�o7��­=��8>��?�?�M?��R>�[�=֛��X ��� �:�<�}�<P��<���=H�d>�H�=�#=�R���=N>�u^�]�o=��y>�+z="v>�[!>�Q�=��=�?��l�������5�B�U�о8G$>&M�<ű�у=̝���&y��Ć�� �2>>:@>��r>rҕ>7��>ﲩ>��>ھ����J�g�@��>⦒>˜�=�Ƈ>ʱD=n{=�=�\=�!>��R=�5�=>�<=�^Ż�7F��Q>��6?��/?ߙ5?P䳽�	Ѿ���Ф��fD�CGn<�n>y��>�{x>���Ѡþ�s���w��x���j���M>�;�>�%;>�=�iּ�@Z��H���v�<�O����!�]��=��>�.>�@>&�<�2����潸�S�j�ȿ	頿�4�_�� �>�s�=B���`���e<-?�K�-�W:���R�ʑ�b����n���>��=�ȼbK���ܽ+��=�z�v_�O�c������+L��G���J߼(��])��H�ھH6A��p"�Iua��"�����{%�����=�@�>R�>��>ZJ?Җ�>�>��b>�~;>�d�����>��J>��>��>/>�d=�k�����]:����ὣ�!���i=���=�{>��M׼*j�=߂ӽ,��=��=݇=)��=W�����5��@�<T=�M> �>� ?�vs�0᥾]'��ʾ�.=���=xu�>���<��=C�I/�8���,�=)c4>Z>�=�y�>�d�>=z�>ݩ�=��� ���G�=-@�=�|�=��E>ʜ��K��;;�=.�>Shl>��f=0�:��^���E�Q��4f@=���=y�]?��?D]Y?��������"�5S���ȾL�+IU�|�>�{��q*�����S,����2��80�����p�>���>��>���=�Y5��>����h�=����y�T� �-5#�ag�<pe�>",y>(��=d���v���οu�8�׾N!T�`�>� �>ӂ���q";�ҽ�~>��L����FOV�����	�.�=<P���H ����9�.Z6����ߞ�����",���'�r�w���'��齂UO<἖�����S#�g-���:[�g������;�����7�<� �>��`>���>_�>T��>L��=Iu���6�=���>��ڽ����)�>���>@N�>7h>�	�>��>ҩA>	�Ԁs�-O��ڀ>��=]r�l�<4�e>�=�<s�-�j��=��Q>�3�R����Sd���(�=\�">��=gPĻf�!?�B����;�վ6`Ծ���I&���h=��)���=�y��k�=��<t�e=�/�=ۖ�<*f�>d��>/��>��}>��z>Y�>����;�^I�a��<�>�v�<e >�����嶼�s!��r<=�y�=�i�=TJ��QxϽ��٣���_�z�}?d�*?l�9?�����%�����`��;���u����>�~~>aD��V }����hؾ�4(���c��.�f.��X�>V�=>���=Ɋ�>�����V�(�.�ֵ�E�Imb>C�$��}=���;V7�=�p1=����x-=8w��Vݿ�b��=婾o0�����=E?>��⽪L>�͸�Srv��u'��v�P������9��I�ɷ�=�=;y�� h�<���"�߾h�����t��M`����ѽ�����;�JھAC1�G�,��=�t�rZȼ�t����}A=Z���b�1>�ݾ>��^>f6? ]�>�`�>�a@>qZ�>S��=ގ�>9k���=lʳ=0]R<�l:>��Q��r�=���$my�E�2��P>ϱ,����=`�>�6�=�b'>�>Y��=�e�=��A>Б�<Ґ�������a�= �_>��^>��?��l�������5�B�U�о8G$>&M�<ű�у=̝���&y��Ć�� �2>>:@>��r>rҕ>7��>ﲩ>��>ھ����J�g�@��>⦒>˜�=�Ƈ>ʱD=n{=�=�\=�!>��R=�5�=>�<=�^Ż�7F��Q>��6?��/?ߙ5?P䳽�	Ѿ���Ф��fD�CGn<�n>y��>�{x>���Ѡþ�s���w��x���j���M>�;�>�%;>�=�iּ�@Z��H���v�<�O����!�]��=��>�.>�@>&�<�2����潸�S�j�ȿ	頿�4�_�� �>�s�=B���`���e<-?�K�-�W:���R�ʑ�b����n���>��=�ȼbK���ܽ+��=�z�v_�O�c������+L��G���J߼(��])��H�ھH6A��p"�Iua��"�����{%�����=�@�>R�>��>ZJ?Җ�>�>��b>�~;>�d�����>��J>��>��>/>�d=�k�����]:����ὣ�!���i=���=�{>��M׼*j�=߂ӽ,��=��=݇=)��=W�����5��@�<T=�M> �>�*?��þ��)�P}�\�ھ����z<�N>��=�y�=ְ����/=�%
>=V:>{�=�jE>/��>!�?��>��;>�;j>/%Z��C�E��������7=�5>h�����;�ž=�R=lM.={I��xA���@�L��e�����<2�?<�?�s_?������)��*/�V��
�&��1=���>�F<��B|��u���뙾ɯ���+���Y�Ė��)�����=�s�>��>^;�>@m9>�lr�t-���><�e=��u>x=�=��=�>�a->si�=�c�=*�)������ؿ�<P� >�PϽ��s>%��=��콠���S�������#3��~k��G������ez���ѽ�ҥ�Y�s�q?�`�	<����-=��!�ܘ�N}��2���9&�6j���P�Vs��M�@�Խ^Ʊ�K���=��ܽ(��������=\o>�S�>ĕ�>�.??> ?Xj>	�>+ƀ>���=�L�>���>i=C#�<�Q>:l[>*3�>\r��=f�H�ؽM =��Z(<!W�<�˔<Eo.>�U�>_��<n�E>WMb=�:��[������<�P�=��_=�'=��%>���=��>��>���(:���?�(��g�4�>��=2��6�H ��,�����wr��o>��>\��=0��:�ɒ>P��>��U�;�g���/>.�p��!�=�� =6�V�qav=yC��=�^j=���=���!&)���^�Y�P�᳍���>Eg5?7?I�	?%r��)�L���O�~�;���W
�>�5?�9>o+���پ�}7�m�Q���_�O�:�> �gњ�x�>�y�>_v�=��k>�����	��w���E�;%�e>e�=ő1>XI=���=u&�=�o�=aZ=�>:쿎���#X���)��3/v>��G>W��>�M�=M��<η�=��=F�>��M>���=�I=��=j>��~=q���z=�騈;ћ�|��Wr�x��d��f�q=;e��1_������I#�퇽� ӽ�N������O"���˽xc�>	�|���2>�z�>�5?��?rD?U��9<�-�>��>)ү=03�>O%T>�R>��=e?#=��>>�>�;�%̄<k�=���;�L=֜=��>,�W=��=�Ҽmi���LĽ�Ky�M���=��>G6>7^>���=B�;>!{A>���=�y����_zѾu9���?޽�z�̑-��./��6�v���T �>��>�ƕ>�Pl���}>���>rf��b��'T>7��|�=T�9�(T����>�i��*�<��a�P��*�M��	6�%#8�Á/���Z��6>>?� �>��>� �����l�,˾y��9����Q>f�>ڮ�>i�������=��##���>�����;�+&>\ہ���=�P=�5���/ �r-M��/=��;��.>Ĺ�=��>���>���>��Q=���
%ɾ�;��v����\r��
�����3�g*>}�<ﱽ��}�0�����<I�<�G�=�I">��<\>>��=��=���==y�����?�%>�}0�>����;K�����=@B��8A���h��վ�R7��s\��e��EG6�Sԙ��x��;���k�>IBƼ�c@����>�A3?� ?-w?��s�k2>|��>�H�>��>���>X�>���>�z�=���L�=<�>�|C���G��+�=��>ࠎ=� >�06>���>B�=����~=q=$>�=�6��_�Ir=��>B�>�)�>=��>���>͝a�2b<���E��J'����D��=yN�=`��=���u!�!&&�J �N�ž�?���=� �>���={��>WΊ>���=�m�=[�h��fr���6=8��=�`�=����K���
�<e��Z�s#�=C����=? )�ɛ�>��0?27?�?)޽]�ݾ7��ܪ1����d�+&�=���<*<9?2����67�2<�Y �1U"���;�b:>��>DY�=�`3>^>Ȼ��=�ډ�J�H�A炾]��=*�>��>���>H �=+���9]ҽ�(��d���8�ƿ�D�����H�M�=�R>�ݝ>ۊ>� >��ǽ��>ρj>�||>��$>��>��>�&>,�1=X��زоq:��'9���{~�D��D�)�P�t�P�=b��	����^���#���z��Cr�:����.e��m�%�x=	a?7.�<�.=��>�_=?\�:?�C2?N-v=
�Y��W9>���>7��>�>��>�?�b�>��#>��=&l�=J�;�`!�	��={��=$�u<~p>���=�S�==S�ѩ,>�>,�/��ؽĆֽ7o+<^c�S*>�5>:d�>�?qh�>~$1�XB��1�>�'�9�H��⛾&�ľ23�L�Q�ôU���I�#c>J<�>rr�>g(>_�*>X+>3�>�5	?�d���CL�^��=��n��{~<ȫ9�K`��Eb`=�ߠ<7��LSi=��c=�?�X�o�l�*�⽵�v���>|�m?�R�>s�>7�<"����f%�3��˽�j�>��>:�c>jP� ��?)�~a��u��LJ���@�DA��^�>���>W�E>7�=u�=&Xc��K=���#=1�3=�h$����<٨J>L�E>mv�=���=J��(AͿ7���~�K������M|���>3��>�4�>)��={��>�z�<�I>> z>���;놵=)u'>�ߥ>|��>3�>9�&�����<Q0׽cǾ��<�܉��C#��ý�n;��������T�ː�RqԼX��<-%���Rƽqz��X��>���=���>�6?M?��?Z�$?���>X	�>���>��?��>�O�>2z��k��k����=t�%>�O�=cJ0�R�"��Fɽ�^.�M`�=\u�={�>d�=P��=���=�P=D��=R�>�<=���=�e�=_J >�ʓ=9�>��>���>��&� ;��D`�vK&��'/�8��RR���m�/�D�bSQ���F�q�@�D>u��>_��>�	�����>B�>�e�>	5���	��""=����u��(��{��`G���ٽ\�=��=���XQO�1��@�t���A�����>��=?O�?�i�>���<��ϾO��E�G���#Ξ�E�}>V��>G��>H$��K�
���ʶl��[I�-R�����MT��e�>�o�>��V>��G>7��=}Y,<�*���ih��Є>�T�R�T�'�$==�y>�QC>u�=M�<�R���ؿ�՛��~��ݾ�>��>�h�>E��>ح�>���>_��;p��=��=��{>�x�=q�^=	c�=��>,Z�=x�c��lg���<��g{����g�:z����1=$���d���yɽ���*!�^/���X7�
�����˽߭��D���>	hŽ��B>=J>?�n2?��?|�:?1s>e¤=3��>�?���>���>��'>�/n<����F�=��>�z>ә0�c�������I���?=�˫=��R>Y�=�� >D�_=Nd˼��=`R(=�>dr�=��=��5>I�v=!�c>O��>�S>;A����bV��CپvY���V>ߏ�=���=�S��</��\þN#�X�]=fl=��t>��>�\x>rl�>K��>��#�!��^߽F=���<���=c2w>�&}>q�?���ezk<�"<_޳=�"�=
����f�����Ay>lֹ>�-?u)�>x��>CC��-Z�֒`�������׭O��?�C�>j��>+Q�{t)�FE�����(��9p�= i�=)��lK)�~SQ>l;�_�=��[=ێ�<~��=�j#>_L>���>%�1>�� =��A=v��=�=Q?��v�ʿ�ۨ��u ��([>�>�7�>�o>i4r>����:��[��AݾB�G�����̇-��f�p����
���+9��r�� 󩾻h�=x��;�E��p���I��>�ܽ��5��Ȏ�+����9���㒾{�-c�1���ߜ"�2Z���1ܽ'n�>N�>66>>��=v�>��?�?�>{ݩ>�Ƹ>vz?�݄�w�|>�����=V�>Qi�>�X���#.>.�9���*���>���>�>29u>#�>��5���c���+��>��Z=��Q��U`�����Aν�>_@V>��>��>3
�=�0��B�����ؾ�4�y��K��>�^��4x��f۾K�]� ��\z4���o���>���>�/�>�	>z'�>��&>5����裾��Q�'o0>��C�w=)���'�>Z�W���L>wj�>/ >#����=��߳
���B>�1>���>�X/? �?��>b[
�4^�	C'�p�1�������;��=NpY>.�=�,Ƚ�,��R&��Ӿ�M<%̍=��?=��=���>�`���"��=ʼS��ߌ��sW���=�<�=c����1b<d?7>=��=`�= '>�s���̿[_����9��)�mCt>���>��=Y����r�N���μ������=e$I>�҄>;��=�>>��3���ݺ݊��P�F��p��F/��1��
��1"��T�~΀�CY������"��\[��qH��h*�-��l9��J���_����>��>#>��=��=adl>�u?*�>�H�>m�Y>�o�>`�=�3�>����3��X�5���(��
o=\v��!ӽ�ƼM�j>�F>ia3>w��<�O>�>P<���> 9�=JҨ>� h��������ި����%����=�v;>Y�<�B?�!�=�׮�ʣ�X�����̾⾜�!=�q��h�0�����r�=V������=1�V>G�>��>=?��Y>�N[>kf�>��վ;N��j7�=� ,��4���Q=��H;Յ=��<���=:X1>p��<B5S��}2��̽I�=�>�=�a>��?~D�>�4�>�w�=��後�ɾ�
��@��^4���@=K{>��=������]���7�����ʾ�GV"�/�>*�U>�\�>�==*l����=X��=�=�UR�$��>�6��=L�|=��3>H#>�CX>.��7��Dֿŏ��J�����_���{�>��6>#��)J��V��y�ʽ; ���@�)=D�x=c�=�P�a��]�½\�P�},�>rt�9�����NF�.�(����L�a�y����������������]��]�H�n��P��C�l�Y>�K�>%�=l(�>zJ�>�Q�>�??|�J>F#?���>ީ??�����>?���\�#�^U>Y�=.���<=�ԽK0`�}c�=e�9>b�t=w�\>ɺ�=W��;Mq�=2�>`��=�x��޼�]�;�v�=��V=�~�=E�>c�=:8�<�xc>`�
�C�����j��c��!�>'���d����rҾV.�� ʾ��<u��>b�>�a�>�Q�>�*�>��>�P=��Ͼ��>>�>z1)���=��>l-W>�^��0�O>���>��%>�N���+��!�����L�<́>�?j�?�r�>�?�tOپ�j�����D�������=�8>[�>+���X����ܾ˃�*��� p��#���'6>�+9>��=!`�=v�O<�@���!�=g��q�'>���u�>��H>���>ԙP>�ڻ=vl
�2�7�Lਿ�H���0����Q��4,�1����n�>2�<���������oE�8B,��2��;��=�h<���=�P�=ǻ�=��>��#�����I���/W�/��
�����1R�T���9���~��r���w����۝��0�O�1�>�iL�vp��oO�>ZN�<X�>���>E&?��?��>�
�Iٔ>v��=7A�>i�=�>�l>_ة>�^2����1��Ӭ����=[,��� ">;0�>U�=�j>���>�!=�u�<�=`<D>n�<��ܽg���+��=�o6=q(�=�n>N�z=�b�>
s=�:��Js¾�!���p�]���JO>��q�(���nɾ9��Ɠ���a�΋k���N>�w|=���>�̈́>��d>���>�w�I��.�r>�5�=<��=�ț�D���ݖ>� =��\=E��=��==�fs�w�Y=�-��՟��W��!��>JK?�
�>q:�>�`���d���(����\����=�?>�Cf>:.A>i3��M��WCվ��ɾe��"���'��F�
>�y�>��g>5<='3�<PE=�ߤ;�>�G)�|1~>$W&��I&>3��=��=H@�=M�=��������@�(�Ŀp����	����=�}c>ft>�a��m�н�Y��8�O�� �����-��c���*W#��4�<�^(�W%'��8�>�a[��5=�A�<���[���ʾ�C��Χ��uþr���WF7<�P��j�̽.�L�]e����t��;��^���l>��>��>.�e>%"�>���>�o�>(r���b�>{�>^��>�1�=B�>��>zB�>�e�=ݾ�=rC�^��:�|�������=�0n>QQ���>͂=W��=8.O>����0A�=��{�9��V��3�=ĦM�}&
>݉�=K�>?�9?J%�>D�ܾ��E'ƾ�2�������&E>��x��1�7�v�����=��ԑ�fR����i>m�>��>)駾��f>g�i>�3���=2�b�D=�޻��=?u=�Y��F���">�D�Q�+���=��b>�Pf>�>�3��n>�+?�*W?��>M,þ��݊� 5������X�=pq�:59>�/��{V�	����M����	V�]g<=|���=�Oq>->��7=��|YJ>=;Ľ�+>���<!�X=+�~>��~>��>�@j=�>8��N�I����>�=�6���򝿮XӾX���c�>*�->��=2s�=@`��T�>�.�̐M�*-�>��N��.J>r
ɻ���;ֽ��)\>�N��|��(=|�׽��Z���1�\>������z5���i���t���&t�N���zQ��1�Ȕ��:��}��4�.�
�=>���>
U>~w,?��>p9?�ٳ>��A>S&?s �����>i��>�>�?D��>�CI>=0w�P�>k޼P�,��+>��.>^\�=X�p>B�
�"�#=�D1><��=╞<���W�����A�'���'<p�U<@=>�o>�� ?TZ4>�Nپ���[]�I�ག��{p?�T��YnB��~�t­������M�>�X�>$^I>3�>8�T�ۉ>��>��ǐ�/>�Dl��1�< \�>"��=��0��+�=s�ȼ ������=�]">3f>:��>�¬��=���q=���>mQ?G�?΁��\�޾���,��W��#@>�V���S��P�����s���ʹ0��%��!Ӿ1$Ǿ	O�=�2:>"G�>�B,>�ν����0��=�[�R�Z=�[�>�<>5>p�>>h=���߼Ʌ�O���c>�F>c�ҿ�V����v��A����8�X#�=
��=�x����[�u>ձ�V=�	�==a\=�G���;��be�=�3>���>���������<A��@w��Ph��\@�W��=[j���K̽\���ጾe�W��ʉ�eMb���3��f�R,n�+3���'�>���>5�M�|��>U�)?�\�>4��>�'=p�>�%���>Q��>���>�6�>eLk>��v>Y�@>����
�>ZS罣af�t>d[�>Rz�=�TT>�X*��Ù�l�<�tĻ2E�q��=���<7��=��<�n����͵��q�>�??���=Yr����'���d�M�iA?X���-�H̚���Ҿ�i��*/߾I�ͽ�ʠ���>���>FQ���>>w>�<z�=D\K=�+����>���\2,����<㦍=�*<@��>��>%E=�!~>���=b���Ix��H>�/?�?�&?&���S�ȓ���2�kDҾS��=_qs<̀�=��=)c��"���2~�������'��_����h�dC}>C�>R�����v��4j���\�<�ۓ>Mp�2#�=���>k��eݬ>�>B�X���ｐ��=�|>��ݿ� ����j�����᰽����L�o-,�c��u7H>��þ�������ƌ}<��ݻ��(��a߽�2�2��=�@=�G��H>��.�囑�\TN��	��9�a=�����9����n)��\@��Ⱦ�?�Ꝑ��n��c��d�ཫ0�=�y>h��>�F&?�R?���>���>��־��?1����g
?P��>m�>��?��p>�	�>�^=��c=�>�^���"�����<n�k��$�=q��=9'�<����=G�=?��<�����3�߽�#���~�;c˓=+.	>��=Eg?/�0�k飾��C�1�_�
>��>"�?xv=r��y�1�Zu�TF��7����n��>��p���H@�>ǀ�>Kʵ>I�>��� ��$5>oƼ�7S=Y�r<y�=2�߽֌C>Xa>����>�"�>��]>�n>ɕ�B3��8�=��?�'?��?A&;:[�侄������K@�sKJ;�U��XJJ=��@�����ʪ߾�D���{�߾�4o�1�����<c��>�y>�D��`<9�A=�����,=)1;7��h�=m�>���=<��=���5r��j��;�,W=�Kҿ���������ξ�3�;[^�.o7�Ⱥ�%
4��T>�I�m(�R����<�F�=��9<�>�:=��y�,�~�lh��>P����i�r��<+���z=�@��K�ա��)��p�N�-낾E	��kG�`����T��8�����g>}�?Y��<l��>��(?M��=�W�=�1�ޒ�=A#��K�>�� >#�<��>�]�>��>�8>� C�vJ�\1�
I5�
"�>��{>�Y��]H�=#�%=p> ��S{<�5�=��t=/h����<},Q����|磽�$�=~��>y��<��#?_.>������ɿ�ZԽ��>�? ?Rz7�vv���u¾Ŵ?��'����5%�<����~q�=�">��o>��r>��>m颾Ո��E�=����=�K"=�K��_����8=VI	>P("���=�=b.>���=���9)*�ŒU>�=?�?��?�V���C5�{n+�=����!=\H��=�K��p9H�BOﾕ�Ⱦ���������x��rz���.��}?{>V#�>LZ!����<N/ ��������>�9=%��>N!>��>�ƃ>{�r�ν��=ɰ">��п�1����=���c�=O�>'�P�����;ž:��>����&2�p���^�h@8:F���U:��a=�j>�a�)Q�b��=������]�b���U���=Ӛ����<$���b���l�νL�X�	�!�~���g���~���I>�X�>Ir�=z�?�22?���>��B>qO���?�gl�g�?��>�ͣ>B��>�Wm>�t�>\�w= ���-�L�s�A�&��=��3>���=
J >!$�<�o=	�=s+d<��Q��m�;q���y��f�=��Tk=P�3=h./>�h0>C�C>�?>t^��c��p��o(�ɔ������#��n��T@���E��e@��L1��3L�Ԓ.�	�ؾg��>�t2?Q��=���>0��=v�W�*�U=]��,����T�:�r��ז�)
�=r�<��W���"�ڗ��!z����5��M&>�R�=Ӱ>�[(?a�\?��B?���T�X��g	��f���o�-w�<G��>�:�=�>?
 ��*��ԥ��?پ��,���!�����;粖>��>�Й>�;<-��EP>�l>v'�=���=��>\��>���>�4�>;5�>O�>����+��t��������˯��/�0���ŽB_>t�}��;}
��ļ�|���4됾��-��;��>����dG+�"?�T{	?.ľ���otm�B��!���~�O����9�M�����v�¾�?��Z��E�ӗ�4��<꤁���Ӿ�X���[�>㼼8:>���<�?ŏ?f�?�F?�/0?��i>��>#?)��>�q
?<?=i?��?x�V>����9L�?(�������ދ�P޽�	�<��7>C8,=�ϼ�R;fg�<5����y�'���K�I,�9tbG=
�=��=C�C>�?>t^��c��p��o(�ɔ������#��n��T@���E��e@��L1��3L�Ԓ.�	�ؾg��>�t2?Q��=���>0��=v�W�*�U=]��,����T�:�r��ז�)
�=r�<��W���"�ڗ��!z����5��M&>�R�=Ӱ>�[(?a�\?��B?���T�X��g	��f���o�-w�<G��>�:�=�>?
 ��*��ԥ��?پ��,���!�����;粖>��>�Й>�;<-��EP>�l>v'�=���=��>\��>���>�4�>;5�>O�>����+��t��������˯��/�0���ŽB_>t�}��;}
��ļ�|���4됾��-��;��>����dG+�"?�T{	?.ľ���otm�B��!���~�O����9�M�����v�¾�?��Z��E�ӗ�4��<꤁���Ӿ�X���[�>㼼8:>���<�?ŏ?f�?�F?�/0?��i>��>#?)��>�q
?<?=i?��?x�V>����9L�?(�������ދ�P޽�	�<��7>C8,=�ϼ�R;fg�<5����y�'���K�I,�9tbG=
�=��=p[���N�=��ܾ�%���ξ[��<:�����R�7�=�%���Q�Y�G�R�P�(��"E��>��f<�2?7�1?lw�=�ƣ>��������<JB2�>^5��o��t>���,�r�P;4ȴ�r�齱	�]��0T
�[���g���N?��r?Ŕ5?;f��f�{�ז	�2\���k���!����>�=NO>=�,	�g��_����־�VM��$�N�>?��=2��=#�=#O>���=0՘���[>n_I>$9�<
^�>�f�>��4>�*�=�۽>�׬>nUt>Ǩ$����I��7(���R%�����'wu����<�CZ��սbe��rY��R�!��S���)-�$>[v�=�1�=��=��<���=+�!�F��jϪ�oܿ��5ƾ(�]�L{;GA|��M���ξy�Ͼ����7��P꠾.����������HM�����ZI?�U���C�K�
>P>�><��>F	)?��	?t'?[v�>�3�>z�?H�?&��>��?�?)�>An�<?i��~�=^��
��=�?���ȼ���;�bf=Gk=B�x=�=�S���
c��V@<H��=&�4<�C;
�"=q(�=J��=WqV>?��S�"�!
����D��🅾ɳ|>��3���hѾK�P�g�;���_.���Q@�>�$���=�0�>�}>�>f�s�(��)�=��< �2; E��G�*������>��k��ܼDNd��>�����.a���$>FY>y����o?�,?@ ?yq�  ��9ξZ�x��x���>,����W�����6���%��о-~ܾ�쿾2��=,�f>��6>���=Yz6=\��=�W���u�<�H>�>�aC>}7M>�ϙ>��>���>���>=v>��[�m�n������Lޗ���A��u���; ���@=n6��a6=�=J��\��9*�L������>��=<B">@��<2��$M~����!ା}��3e�!�˾���:�Ծ�)\��$���=�������Q���_���-��E�����1E���a�S���>�pf�
�>�S�=��-?��6?��?j��>��>&�>ӳ_>͙�>�?	v�>��?�?�
?���>�T=BS�;7����g.>��=�H�=���=�>���>1c�=��=�@s�.�<�1C=0��wj=�=��=��>4�L>p[���N�=��ܾ�%���ξ[��<:�����R�7�=�%���Q�Y�G�R�P�(��"E��>��f<�2?7�1?lw�=�ƣ>��������<JB2�>^5��o��t>���,�r�P;4ȴ�r�齱	�]��0T
�[���g���N?��r?Ŕ5?;f��f�{�ז	�2\���k���!����>�=NO>=�,	�g��_����־�VM��$�N�>?��=2��=#�=#O>���=0՘���[>n_I>$9�<
^�>�f�>��4>�*�=�۽>�׬>nUt>Ǩ$����I��7(���R%�����'wu����<�CZ��սbe��rY��R�!��S���)-�$>[v�=�1�=��=��<���=+�!�F��jϪ�oܿ��5ƾ(�]�L{;GA|��M���ξy�Ͼ����7��P꠾.����������HM�����ZI?�U���C�K�
>P>�><��>F	)?��	?t'?[v�>�3�>z�?H�?&��>��?�?)�>An�<?i��~�=^��
��=�?���ȼ���;�bf=Gk=B�x=�=�S���
c��V@<H��=&�4<�C;
�"=q(�=J��=��!?k��>��S�����&��с�]����S�Z)d>@:�>���
#I��RE��<�w1O���⾾�>�.��a�>��>"V!�����L=�0齁�#�>���?
>��<3_u�����Al��
��<7qѽ��$:�	ƽߘ�>:5?ܹ�>�B1? N��
�*�EJ�``��v'=�]�=8g.>X=�>�Z>������Ծj�#���}3	�_K����,>e=bT> ���[=.+�<4JT�9ez�}�7>H
�7B>�!�>[.t=�3�>�.y>��!;<�<n�r���u�J6����JH۾��龳��>�����lE��ѩھc4�����s�~�=�Q�>���>*��>���>a>�d>��ӻn���/�=��I2��9E��-ེ��<���B���߄�W"���j=oh��_B�񓭽Ht	�R�����ý��c��_�>��R>fh>�jL>̂%?b5-?�?��>JS�=����1$?���>&K?���>��>�yD>
=T�9�C�I<��Z�͊L� e�=VX�=g�=p�>l�0>&�#���S;���ø;k7ν[�\=Vđ=c%-=�<����=>>(�6>؃�>��!>&6�������#������P���>�~/�e��>b��&�ɾ���M|��l�o�c�\��<r�>�h=f*>��>�τ�����>�}޽(���z>�<W�hkh��5���#����q���<���RÇ���C=�)A�S�(��x>��?kD?�4?�ꑾ�8����Q(V�+���r=a����=��%�<Ѿ��پ]]l�����þ�@��+=�{	>��O=��X���*;�� >���#/T>O�>�����=&D�>G�>�dd>}:�>嵇=�JF��O�j�/�<��|�����8Ⓘ�2����>9^�=ʶ������-�<|������T]>��>��>�`�>5�=@`'>���>i��
����G>E�w=*�&��.=�_D;�PB����-�4�>Fz޾��ۼ�氹[�ʾ4����W@����w���6_<[q�>NT{>�M�94�<==	[?e0?�?E)B����>N߹��m�>��>��?`�?���>I��>e�Y>�"������{7>���`����=0(H>C��<�Ĵ=��>|����<2 �<�N�>�b��I}<���=pXW=ĩ=�Y>�R5>�?>s�?�KY>*C���`���S^��J(��@���?��<k�>_$�}�'��LL�g����"�d]>V��>n��>#Y|��|�>�s�>M�|�4ƞ�E��>/+@�A��=�ط=4Z�Ʋ5��hk=w��<��x��l����o>Ԑ$=5t��l���]>�u;?;��>��?����OT%����v�!���߾��=���KU>(Y�<�}�4����u7�RFؾ_u$�^�ƾc�	�2��=��l>��&�%�x;�y>s������<�.�=�A�T�T=)}>�ï>���>�y>K;3���Z��
�S��£��������h꾴� ��%>���=�:n�p�Ľ*_$=��˽��=pNh>RȊ>^e�>(&	>�A�=���=Z�?W�	��Ѿ�eӼ���M���ې��s����e=�½�Ĥ>p��H�0�XRM�z�h���e��;�l3�K����1�BBQ>YIQ=)�Y>8l>\�4?d%?��?�Qʽ��E>�����?���>'��>�?5��>m�=*[��D\�D� �(4��ē;�;��=j�<>��K=5>G�=�^�Xp�=`"(=�>>9J�?%�=���=hWP<���=�>[V>��z>�"?������ھ�w�=X�վF���,Ͼ��>�ϾB1g>���P���$������u*>z�>�<�(Y>LX�\�>���>�"���f�Ԋ6>@���	żq�>��C=M'{���[=��6>gܚ��ݩ�����]�G��������f�
<�>N�5?�6�>@T�>�=���� ���e��ZA���_�bY�=F+�>RT�<>&�C����L`7�3�#�:ؾf U���2>��G>B�>tA>�i�<q��<�岽��=�&q_>m��Y[�=�l�=_~t>�&>�l>�g�����sӿ�ӯ���c�Ei��1���H�>�=��E����J_���ٽo7#���k>ew�>g>D9>���>8��=N�&>�
���Ͼ�+>��^�x漾f�\�������=I��{�W=Ǧ���� ���%�Ty̽����<Z��>�G�WD(=X�=v?��>!��=�j?C/ ?�[?+g>��?��b���,?��u>���>q�H=$�oH�y�=�T� �>(u��T���=ޘ�=�����e5>��>O	�[��=�z�<PI�=IL���ƒ=�V�<%���!�=q6�=���=�b=��?s��1Ǿ�=Q~�����=�>�r�����=?����^ɗ�Â=�9>��>�M>��N>���>��>��M>�'��/�H�8��=Ž�ZC���=�����=��8>��=�1�������yU�X�#�&��=�a�;] >Ns2?��	?�*�>�a >9㭾P.��~�;B�����
>��K>s�=�/�=M틾�5վ)�#�Ҵ�p������Ϳ��W�>=�~>7��>;g8>!�=���{K���>�9��թ�=�Zf�2ʼ=�.>b��>���>·>-M'���|�{fۿ�������=���!�=��=�R��~a��F]��X����� ��� >�&W=��+���ٽĹ��i�n�Z�}>Ai��ԁ>�5$=�d�V���5�B�d=�%�@R>�@Ծ��e��F���	x	���5���L�����!�:�D=*7#?��=>I'�.� ?�x=?t�-?ϫ����?��D�2A ?y��>���>�<1�2�
�!�~YU>�B�>
U;��ɤ�������=��H$Z����=1�>Q��;����U���rt����=jk=�z*<���`fB=.L�;�m�=x'�>�"�����H�D<�N����xЎ��~<5�������B��B<���7�=���=ޜ�>Ҡ�=���(f.>$X�>�L�>����ML����>t�H�c��l�=>\.��d�=TXt�8<��}�ҷ�`�>1��=O�;��=��6��o>J^?��*?]/_?�Y��g�������!�������>?�<Qs>F�����ξ����޾�m��tZ^��M^=ex�=��~��������iy�\,6�?�1>��>�WW>��>|�o>��>��k>t]/=�	�����,�������ƿq���.���\'�j�=k�>�.�>��p�0���Vg�b?��@�=����������������<X,�>����Z��a<p�����ž���<�sv��4��ol��ǳ���l���
������\���������.�d�_��5�p�;�
?�?j��_����#?A9�=�Y�=K��>=�?�D�>J�>�Y�>�E�>�yc>T��>b�\>ye�>�h>Td��"���#=ϋ�>�ha>iV�=G�=P��>�J��Z�L��5�=�� >׀
>�{��Q$鼐"���|=g`K>0t
=2�>7�>�D�=�n���t�����Z�������t=k8������*�)���K�n���f>�U�>��?p=�m�Vf�>�#w>��>���#_�WT >��l�p>I>���t���&Y��ͽ�1Ƚ׽1��M�{�H=ħ>@�e=�:�<��>7�C?�U$?�?v(Z� ��h)������M�=��>>qV>t�>��|>�b��Ǿ��C*�Q��@��F�R��&w=J2%>�ٶ�|�d�=�:�q��&��> ��<Y��:�,�=��@>g�>#Wy>d�K>�';��r�[s%�O-��\벿�1��\T��̻��BE� |�>�^>1�нR��=�'m>Z�u>:��?����<��b���܃���>� ?fי>��u�k���U�� uC=�Z��4m�����E��ob��E4��i둾�T+��H��y/��}ݽ�E˽��?�gN=�nd��P+�><�>�5�>B�$>��F?9��>�P?Ufj>��>�f>�v>�%R>b�(>>�1 >�侽L���%�)����(���|�����>���>\�&=@��>�->�ǝ����=N\�>n6�>2o�=d�M�8
�<��2�Xԕ=�;Y==3Q>��z>x'�>�"�����H�D<�N����xЎ��~<5�������B��B<���7�=���=ޜ�>Ҡ�=���(f.>$X�>�L�>����ML����>t�H�c��l�=>\.��d�=TXt�8<��}�ҷ�`�>1��=O�;��=��6��o>J^?��*?]/_?�Y��g�������!�������>?�<Qs>F�����ξ����޾�m��tZ^��M^=ex�=��~��������iy�\,6�?�1>��>�WW>��>|�o>��>��k>t]/=�	�����,�������ƿq���.���\'�j�=k�>�.�>��p�0���Vg�b?��@�=����������������<X,�>����Z��a<p�����ž���<�sv��4��ol��ǳ���l���
������\���������.�d�_��5�p�;�
?�?j��_����#?A9�=�Y�=K��>=�?�D�>J�>�Y�>�E�>�yc>T��>b�\>ye�>�h>Td��"���#=ϋ�>�ha>iV�=G�=P��>�J��Z�L��5�=�� >׀
>�{��Q$鼐"���|=g`K>0t
=2�>7�>�D�=�n���t�����Z�������t=k8������*�)���K�n���f>�U�>��?p=�m�Vf�>�#w>��>���#_�WT >��l�p>I>���t���&Y��ͽ�1Ƚ׽1��M�{�H=ħ>@�e=�:�<��>7�C?�U$?�?v(Z� ��h)������M�=��>>qV>t�>��|>�b��Ǿ��C*�Q��@��F�R��&w=J2%>�ٶ�|�d�=�:�q��&��> ��<Y��:�,�=��@>g�>#Wy>d�K>�';��r�[s%�O-��\벿�1��\T��̻��BE� |�>�^>1�нR��=�'m>Z�u>:��?����<��b���܃���>� ?fי>��u�k���U�� uC=�Z��4m�����E��ob��E4��i둾�T+��H��y/��}ݽ�E˽��?�gN=�nd��P+�><�>�5�>B�$>��F?9��>�P?Ufj>��>�f>�v>�%R>b�(>>�1 >�侽L���%�)����(���|�����>���>\�&=@��>�->�ǝ����=N\�>n6�>2o�=d�M�8
�<��2�Xԕ=�;Y==3Q>��z>7�>�D�=�n���t�����Z�������t=k8������*�)���K�n���f>�U�>��?p=�m�Vf�>�#w>��>���#_�WT >��l�p>I>���t���&Y��ͽ�1Ƚ׽1��M�{�H=ħ>@�e=�:�<��>7�C?�U$?�?v(Z� ��h)������M�=��>>qV>t�>��|>�b��Ǿ��C*�Q��@��F�R��&w=J2%>�ٶ�|�d�=�:�q��&��> ��<Y��:�,�=��@>g�>#Wy>d�K>�';��r�[s%�O-��\벿�1��\T��̻��BE� |�>�^>1�нR��=�'m>Z�u>:��?����<��b���܃���>� ?fי>��u�k���U�� uC=�Z��4m�����E��ob��E4��i둾�T+��H��y/��}ݽ�E˽��?�gN=�nd��P+�><�>�5�>B�$>��F?9��>�P?Ufj>��>�f>�v>�%R>b�(>>�1 >�侽L���%�)����(���|�����>���>\�&=@��>�->�ǝ����=N\�>n6�>2o�=d�M�8
�<��2�Xԕ=�;Y==3Q>��z>Į�>�R>�mپ�(�H�0��񣾛��]��>ƚ����>�s��h��B�)�޾a{���վ�\�e�̾���u�>�;�>���6�b�͚n�%\&��� >�=�u�=�мH��<kq�C�S>S1�>u1W�g�O<c�
��E������>�"??y�@?�d�>�i��6��T5��$��Q���(;����=`d>��>��b�ߑ������'�ܘ
����/d��$>�D�>~f.>��>���)� ����=�t��D�I�<Y:>\˕>�{�<���;��d�Ex=>�[��(��Y)�x\��r��ȉ¾���׺���>�==��c�Խue�=?��J��8��0����>3�,>��i>�o�=s�T>9랾=?����>0�0`���	-�f����%�\�f��Fx����ҽ�Ͻ�￾������ڛ��Gc�H���'��>t0�� >H��>�7
?�7?��?@R*>4n�>�x���>>�>|<(�9��>#�>s��>g��>�t?sK�>�T�å��e�=�J>��=�>�=��=����
�<��=�O�=��Q������#��
?�=y�=2�?�=_:�>r�>�6>�S5��|*�p(W�j�C���I�>����>��.^�JR�=B�#�������V�0`���ӾXm�>�/�>���=��!��AE��-ٽ�?���;����R���_�����>���={T%>�^����=[��s�򚊾��>{=?�xf?N�?e��I��L�F8@��h��S>68>�05>:{>����2��*:��3;��:�-�ꬢ��~<>%��=6VO=�=>�b=4��<�zw>�>eX�;,�w>��=�/t����=��N>�B>�?�=X6!>�~�;�{���ᠿ��V��^��|�=ȲѼh�#>�X�<Ċ�	e�����xØ��|��&�=�#�>L��>���>��>�_�>N�?�9��meM�ɼYۑ��s8�W���"����=0Ͼ��8��cM���X��.�UF�����-k��{�S?R�>x�>�z>�&:?�?��?+2c=;@? .��j?�e?��E>���>Q��>��>S�?��>K�>�0�]$�kT��o�=�S`>�a�=T�=>�]�;�M:=F��������\<l|���M�;��H=9��=v�=�>��B>Į�>�R>�mپ�(�H�0��񣾛��]��>ƚ����>�s��h��B�)�޾a{���վ�\�e�̾���u�>�;�>���6�b�͚n�%\&��� >�=�u�=�мH��<kq�C�S>S1�>u1W�g�O<c�
��E������>�"??y�@?�d�>�i��6��T5��$��Q���(;����=`d>��>��b�ߑ������'�ܘ
����/d��$>�D�>~f.>��>���)� ����=�t��D�I�<Y:>\˕>�{�<���;��d�Ex=>�[��(��Y)�x\��r��ȉ¾���׺���>�==��c�Խue�=?��J��8��0����>3�,>��i>�o�=s�T>9랾=?����>0�0`���	-�f����%�\�f��Fx����ҽ�Ͻ�￾������ڛ��Gc�H���'��>t0�� >H��>�7
?�7?��?@R*>4n�>�x���>>�>|<(�9��>#�>s��>g��>�t?sK�>�T�å��e�=�J>��=�>�=��=����
�<��=�O�=��Q������#��
?�=y�=2�?�=_:�>r�>�6>�S5��|*�p(W�j�C���I�>����>��.^�JR�=B�#�������V�0`���ӾXm�>�/�>���=��!��AE��-ٽ�?���;����R���_�����>���={T%>�^����=[��s�򚊾��>{=?�xf?N�?e��I��L�F8@��h��S>68>�05>:{>����2��*:��3;��:�-�ꬢ��~<>%��=6VO=�=>�b=4��<�zw>�>eX�;,�w>��=�/t����=��N>�B>�?�=X6!>�~�;�{���ᠿ��V��^��|�=ȲѼh�#>�X�<Ċ�	e�����xØ��|��&�=�#�>L��>���>��>�_�>N�?�9��meM�ɼYۑ��s8�W���"����=0Ͼ��8��cM���X��.�UF�����-k��{�S?R�>x�>�z>�&:?�?��?+2c=;@? .��j?�e?��E>���>Q��>��>S�?��>K�>�0�]$�kT��o�=�S`>�a�=T�=>�]�;�M:=F��������\<l|���M�;��H=9��=v�=�>��B>Į�>�R>�mپ�(�H�0��񣾛��]��>ƚ����>�s��h��B�)�޾a{���վ�\�e�̾���u�>�;�>���6�b�͚n�%\&��� >�=�u�=�мH��<kq�C�S>S1�>u1W�g�O<c�
��E������>�"??y�@?�d�>�i��6��T5��$��Q���(;����=`d>��>��b�ߑ������'�ܘ
����/d��$>�D�>~f.>��>���)� ����=�t��D�I�<Y:>\˕>�{�<���;��d�Ex=>�[��(��Y)�x\��r��ȉ¾���׺���>�==��c�Խue�=?��J��8��0����>3�,>��i>�o�=s�T>9랾=?����>0�0`���	-�f����%�\�f��Fx����ҽ�Ͻ�￾������ڛ��Gc�H���'��>t0�� >H��>�7
?�7?��?@R*>4n�>�x���>>�>|<(�9��>#�>s��>g��>�t?sK�>�T�å��e�=�J>��=�>�=��=����
�<��=�O�=��Q������#��
?�=y�=2�?�=_:�>��>\��:ob�����B��P�iCd;\��>�W�<?��=Ԍ ��Ǟ=�Ж�xϏ�A=����i=i蘽�Q>f`c�i�>�s?�D=�x�G��>�&���PR��Ի�m��>�=c�%<x�j�M��=L�&=���(C�����=ٖ�=hp�=��r���I??�o�>��쾲7@��/M�Ec����:��E=U�H�Ҿ`N2����YG���k��6i� �1�_�`<}%�=���=��I�4ؖ�U�>U�>�S>3�N>��p=ﾸ=�U<;��=Y>4k�>W�>圼=�e;=�y�y�߿܌����a7�dQ ��%�=��=����������&��=��Vwt�����䭭=�׵=*	i>�ܦ=��=�:>L��w>�������|�q'��̾j�������=� �;P
����=���n��eu��hi��&���%���d�Ž?������ç\>8�3?z$?K�>My�>���>�a�;w�>���=^��>h�?[ֺ>�>��?%�>���>lR���]����~O>���=�D	=ç�=v��� h9�����4#>��I=`�,�=��;2d�=%;�;���<Z��=��>\��:ob�����B��P�iCd;\��>�W�<?��=Ԍ ��Ǟ=�Ж�xϏ�A=����i=i蘽�Q>f`c�i�>�s?�D=�x�G��>�&���PR��Ի�m��>�=c�%<x�j�M��=L�&=���(C�����=ٖ�=hp�=��r���I??�o�>��쾲7@��/M�Ec����:��E=U�H�Ҿ`N2����YG���k��6i� �1�_�`<}%�=���=��I�4ؖ�U�>U�>�S>3�N>��p=ﾸ=�U<;��=Y>4k�>W�>圼=�e;=�y�y�߿܌����a7�dQ ��%�=��=����������&��=��Vwt�����䭭=�׵=*	i>�ܦ=��=�:>L��w>�������|�q'��̾j�������=� �;P
����=���n��eu��hi��&���%���d�Ž?������ç\>8�3?z$?K�>My�>���>�a�;w�>���=^��>h�?[ֺ>�>��?%�>���>lR���]����~O>���=�D	=ç�=v��� h9�����4#>��I=`�,�=��;2d�=%;�;���<Z��=��>\��:ob�����B��P�iCd;\��>�W�<?��=Ԍ ��Ǟ=�Ж�xϏ�A=����i=i蘽�Q>f`c�i�>�s?�D=�x�G��>�&���PR��Ի�m��>�=c�%<x�j�M��=L�&=���(C�����=ٖ�=hp�=��r���I??�o�>��쾲7@��/M�Ec����:��E=U�H�Ҿ`N2����YG���k��6i� �1�_�`<}%�=���=��I�4ؖ�U�>U�>�S>3�N>��p=ﾸ=�U<;��=Y>4k�>W�>圼=�e;=�y�y�߿܌����a7�dQ ��%�=��=����������&��=��Vwt�����䭭=�׵=*	i>�ܦ=��=�:>L��w>�������|�q'��̾j�������=� �;P
����=���n��eu��hi��&���%���d�Ž?������ç\>8�3?z$?K�>My�>���>�a�;w�>���=^��>h�?[ֺ>�>��?%�>���>lR���]����~O>���=�D	=ç�=v��� h9�����4#>��I=`�,�=��;2d�=%;�;���<Z��=�5>��;���Uξ*A�s���1�_��=c��<���=*�J�\�2҉��9�<��;�!����F�O��6=�'!>��>����&z�����g�;��4>P0>A�+>C>�}�^5t�g�S��e��p�
��Y��e�=h/�="�@>�g��7>O� ?�>�7�����Ce=�u���==xϽA��v��=.��� ������&:���1�����X=�ߠ=�[�=�&�-_�=j�>��=8����l#��vH=�ق�?`�=�J4�X�> §>�a�>�ez>��}�X���_��ࢋ�a灾)	���,=R?������Y���w���Q�=�t�����6�7���=��A=8j[=_<�0�<��=�Aξ�}X�=���e5��]Ӿ�	ھ/�;_o߽Kнe:�}���gC���+S�d�X�o�����������SP�䰏���>o*b>��t��=j�?wd,?Z�'?Ł�>�ƽ8�=ӳ�>���=���>D�>�?�-?@,?AI�>���z���.��>+�>���>�a`>,�
>�=Tq=��)�c��U_M>�b@>5���yս;����a��h�=b,>��J>F:v���;�~�a����L�������3/>JY�>[�O>}��mϾ�5=
"�=��������M�M8ݽ�-)��:J>|�=6:�g����|�>X��<,;��YE�=M��!̘�ƴ����#>C�;�߽�`� ��<�J��ʾ����`=<h<Fj�>A'?��?�-��{���1�ڕ���%־i.z�v+K>@T>�}O<�`��gT��q�_��f�!��0���w�=#��=_�J�B^D��6=^_ �XE$�eP���ɲ�Q��p?>��>�kr>a��>�A�=0M=h?�^=���������T��� ����þQ�]�^*����=K���6^����=!��r���?6�]�ƻ^QU�@�W��޽�=�Z�=)^��L� �ˈؽ�mJ�k���ƾ����tO����{��C�����K0e���������=�NT��
�M��`�8?�{�=7mG>�>��?��?q��>�ǋ=�B��z_3�8��>��>�I�<�J=u=�>JF�>��>�|�>�p>$?��72m��.>�a�=>za�)V�=��>zl��ּ>Z	>��2=ݛ޽M���;6����<�7�\�=��>�,;>1J<y�Ͻ�=	����P
��)ƾ(9��mBc=ʀl��>�����ٷ��㾡�;��[��y�}���+��lA<��-���>J�>�]��Oz����.��;'�*��<@�,��q>ǉ>�~>Ʃ=g�c�}�Q�UZ2�Rm1>~�>��0�>l��z�6?�ђ>�x>4a��L&�>���.�z����m��o�=�)��/+/�*�����ԾS�3��2�Г!�P��6��=;.=j��>�/>� �=P�3>`�W>���>Z2Q>��n�vs<��&>��q>>�q>�M�>� �>�
*=�P�	P$>����眩�������3�Z�=Ѡ�=c�3�pL��@�rQ)��F�݉c�!W4��E>��q=ȡ�>Ay�=��0=e\>�0$��ž�ȹ� �P�N�ʾ#ǾY���7��j�y�B���׾u�ž<|ƾ����\���d�� ��_��܈�����>ϯd<Q�>�i]>��?��;?�93?� ?��?�|��"?>�
�>�t�>���>�?b?��!?U��>�A�>r�=��ٽf�����>~p>7D>jP�=���U;��<7��=0ӽ��^�w�'<��B�`3=��=�1>% �=W��>D�	>�ɵ��� ��yJ��=b>5�$�E1>���>�բ>�ɾ�y��f}�����v�/�����������=5f?NJ�>0��>��a�i�O�R��<@5R�*c���И�*���C�=u�̽��J���h>f�P��K<��}��ζ�N�B>ҹv>J��>�1?ָ>7��>���(�"Ͼ�8K�dǸ�>?�=5ꃾޣ\>�f�=���Q��Y��m
�����^���	*��4�=�<L>��=�#=�P���
�=���=�w�z�x�J��>��|>�(�=J��>�
?-�x>g��>Qm��k�#�M��J������?��iބ;��=�N>��=�彌�ɽ�kӽ�3[��*����>�U�>���>Az�<_t�<Ks�=���ҕ̾ �d�;�'��r߾3�ֽ�
��
�<��ཌྷo >�י��"ȼ7C���'�)1�O	+��Ų�bN��������>����>O�?c>?
{)>�V2?FD�>a�<-�����?=��>6 �>��%?��)?��?��:?p��>�ਾ��T�Si��8?�=J3�=M�,>Q�l=ێ	>p�>�cz>lW:����s�H����'ǽ�Ȅ=�>=/�
>cG>1J<y�Ͻ�=	����P
��)ƾ(9��mBc=ʀl��>�����ٷ��㾡�;��[��y�}���+��lA<��-���>J�>�]��Oz����.��;'�*��<@�,��q>ǉ>�~>Ʃ=g�c�}�Q�UZ2�Rm1>~�>��0�>l��z�6?�ђ>�x>4a��L&�>���.�z����m��o�=�)��/+/�*�����ԾS�3��2�Г!�P��6��=;.=j��>�/>� �=P�3>`�W>���>Z2Q>��n�vs<��&>��q>>�q>�M�>� �>�
*=�P�	P$>����眩�������3�Z�=Ѡ�=c�3�pL��@�rQ)��F�݉c�!W4��E>��q=ȡ�>Ay�=��0=e\>�0$��ž�ȹ� �P�N�ʾ#ǾY���7��j�y�B���׾u�ž<|ƾ����\���d�� ��_��܈�����>ϯd<Q�>�i]>��?��;?�93?� ?��?�|��"?>�
�>�t�>���>�?b?��!?U��>�A�>r�=��ٽf�����>~p>7D>jP�=���U;��<7��=0ӽ��^�w�'<��B�`3=��=�1>% �=W��>D�	>�ɵ��� ��yJ��=b>5�$�E1>���>�բ>�ɾ�y��f}�����v�/�����������=5f?NJ�>0��>��a�i�O�R��<@5R�*c���И�*���C�=u�̽��J���h>f�P��K<��}��ζ�N�B>ҹv>J��>�1?ָ>7��>���(�"Ͼ�8K�dǸ�>?�=5ꃾޣ\>�f�=���Q��Y��m
�����^���	*��4�=�<L>��=�#=�P���
�=���=�w�z�x�J��>��|>�(�=J��>�
?-�x>g��>Qm��k�#�M��J������?��iބ;��=�N>��=�彌�ɽ�kӽ�3[��*����>�U�>���>Az�<_t�<Ks�=���ҕ̾ �d�;�'��r߾3�ֽ�
��
�<��ཌྷo >�י��"ȼ7C���'�)1�O	+��Ų�bN��������>����>O�?c>?
{)>�V2?FD�>a�<-�����?=��>6 �>��%?��)?��?��:?p��>�ਾ��T�Si��8?�=J3�=M�,>Q�l=ێ	>p�>�cz>lW:����s�H����'ǽ�Ȅ=�>=/�
>cG>/�?�f�>+h��b�ʓC��^���$�|��}�=��[>��;c�������j���=�H^��<A	�Wf�+� ?c?�>�w�>Fu����e��������=��(=�X�=�O]=I0�=Y�,��:	�>��Y�Y��<i��rý�<�>cbV>��>C�9?N?.�>�>�R��$b�c%l�#��@U\>�Ƚ��K��y�����*о��%��e�R�:��u��sV�kF>���=�x����>;cѽOr�@�T����<�Q�G�7>�0=��ѽ ɖ>��>���>�W�>�3{�������ڒ������߽z=r��<�p>�m�>pB�����{���P9;>l�=G?�>7��>�n�>�W�>⦟>Җ�<��Y���D���=�S"���y3��@|��ء�R|��f�e.���	��A���������ѩ�b����-t���>C�>�R>��>�?�?�>4?yv>j��>8�Ž� >�z�>.S�>ʸ�>��?�?��$?��>�¾?k�����>#��>�m|>�9�=�OM>!2>(؁=�׃�]�>+�=�
�=�=��b7���\�=���=� H>��g>)w>w�=�Cػ�/��qb�U��c��1'�>>���>{�w�oy߾�!�:WE�o-E�I��v���*�>	L%?�ض>mP?���n>ڦ��lG�u������:>~!̽4f0>@%�=��)��<��Ҧ�W���އ�s`~�J
�>��>QP_?�m+?��?�É�.<��0.�\P�r>���'��f�>�(>�A>k;��ao�]�����c�yн��r�3��=�f= ��aJ�>xG�>�b�>F����u�=�����X=>+d�>���>3�>Jpq>g>�ꏾ�9�t׿�I����l���>�Bg>#��>��<��>-$���^?��7�	G���,��%�)>E� ?e��=��>%W�>Z@��HӒ�)���e��<��ܼ�C�<�Y���L>�v��x�V=�6��/�HN"���ݽﾼP�μg���> ��G�B��>��9>�>>��>6!?��?yH?�e
��J�>8o�:��;4}�>JX�>з?��>gq0?�:�>o#��WFC�6��F�-�wt��c��G����/=M�>\}H>�Q=>)�>�&�=�蹽Z�����WRX=�=�W�=��>�G7>���>��A>X��>��n8L���������hQ�>�K<e��>�"�O}%�o��?�5��kD�S��8��9]?;�?I:�>���>������Q�D>�,��s�<�N�sI��o(=E*��ռ6��pݎ��5�/FӾ)�C���>��f>�ϒ>�"?��?F�>f��d��8�*�ҥ-��`���=Mvs>��E���[>LVW���X�P���@�9❾a|�<v&%><� >��߼��'=��=l��@�n�z$��&��
�8>r�>5�>^�>�(�>�I�>?�>�\��5���7߿�����7����������M>����F�=80�>�5R������>B�>$d�>Q�>y�>p��>(�>��8�����թ���:>�;X=j���m�<�����ޕ��� ��U2��B��&(��
��pɚ�=4��hA!=�S��q\��aBӽi��>>n�'>R��>��O?�s?�?A?2^<��!�?�þ�_ҽt�>8��<���>jk?���>��>�|���Z��/���M�r��<��ӻ�>>or��P>�)P>Ĵ�=hS�=��B=K�����<sd8����<׃�=lͻ�5q>ۊ>>�>kf�=eB�#2���c���޾�M�"��>,��=�/?���C�P����G�2�0�P�վ�!>�i�>�?��>�a
?|���aC6�3�=���4&�BTe�xNL�rc> %>֜f>6=-��RX��������oyX��m>6E�=m�[>�"&?��>Ȫ>�>p�ɉ%���G�����Қ��Z��lQ>�q�>{ά>~0�{W������ktȾ�������I(�t��;BK�>�*�=�z/>�:l>ɉ>c����M��H�z��=� ???��>v�>�A>A|������\�QΪ��Y���Ӿ�;5��o�=�F=�*YO=v��>��=��=w� �蹃�:�.<P�A=,��>~>�ڧ<"c>����VI�D�P>^��=)`��T�+�(�� ��(�i�
Lݽ+�b�ݑ��V����i���ֱ�v�.��b���XR��.ڷ>xm�=}4�=��>��-?�?~�5?d	W�|�ѽ�g�������P<:�6>�4?��>�2�>��?�^�<Lׂ��H�R���ȼaB#�;v�=}4>�e>��L>� >�k�<�:U��m�4��K��9��݆�=0��=��C>��z>3"�>�f>��<���]J�����cľN�>|�F�D��>J��Ҕ_�M�F�����0�#j�����>A�>0�?�>� ?-���{u]�<?9>Aȵ��J��_=l�b�=½6>�w>���X�l���Ke��U����w~>�Ix>�_�>�??7�E>��>��%���:�ɁB�:�,��,=]�F����=4j�>�"�%rȽ�>���I���S�)U��
l���j=CC��W�=͖h>�>�u�<d���@�<GT��Z�g=��4��:>r��>��?�Z>���=��?�,'���׿4좿��h�۽|�=���~><�$>KJ$>ޝ>��b��E�O���=��%>V��=�D�>�t�>p� =RZ$=3ɞ�~t��t��=���a�%���ӾR�����/L)��R�� C�keϽq	l�5l���;R�$�y����� C����>zW�=\_n=���>v�A?߯<?�<?�� ��E��j�����=��(��?�=��>d�>|,�>�?#�^=�"�}�lb��}Bu>/9�=<�=� �>.k�>J�n>���Ϫ�<2Q��Ӡ4=���=	��]���x>f�=��>���>��>Q->|D�>�"��o�����̾�G�>P,���'?�P�N�>]���r_A�D�-�d����3�l�>���>8b�>��?���LG!�VFC=#!������������ɽқ�Y����=����tK�ހ'�wNm�����<b�=��=���>�O?�*�>�u>���7�%��F�������F�N�=�8�=�@�>�s(���>����׾|t.�`Ҿ�Ľ_�<�\[=e�'>�n�>6��>Ô@>�!���=�v�r��>�����!>1ś>�p�>K�m>��>���O.̾Y�ܿ�¡�Q��-��wr��{�=��R���ʼz��$��=Q�?���銾�p>LJX>$:Q>]�0�Dl�=I|�>b��9И��a>�霽gE ��'��o��6��ώ��[5>�=v��c<�؟<PH��[I�/���ǾSc���Ƽ2��>�P	�)a��� ?��N?.rC?�Q?��,=:��>-���$!��>����<f��><y>�K?+G?�8�=�E˾O\B�� I�m/��>s=Oި<��D;Pc�=�z�>�	>?�	<�������;�1/���Ʌ��L�=q�=�>C+6>�?T���#>P镾M��>�h��]k�>yv%��|�>�ž�,�%1�|~L��z&�d���UϾ$]�>h)>�d�>"Hn>�^�
�4������\��+9=�㴼v1�=��=?�>1*�����?O�=@�b�U���ݪ;C{>>��>���>��?ƫ�>�T?,�{�M��l?c��׾|��V����
��l��櫡:����zݾ�O���3��1��>[¬�?$�>�
>��=P�>�/l>Z����{�4:h�����z���v<�R�=�=��>.��>"��=w��������m������F; �β��̓�=�?�([����Ͼ8ş�Qe��˘z��熽��>�B{>�Hs>�ԕ=Q���i�3�{�FDj��:>BfA�	��3��V���@r>0�l��XV���s���<P�n�F(ƾ�y�=��dJ����!�'�f��E�=��>Zn��M>�;?at,?tW?X��?��5�H�
?$��>��9?�.<?*i5?@0?��1?���<�=*��紽�h�.�S=&l=��	����=�8�=��@�1>�c�=z�ؼ�|c<�_�=L7�=�>Q�=��=��=l`>ũ?vS�=�(�<��z��b�~ھ6Ul�7*�>��^��?�6>g��=q'�D��>�%�w������q\!=�?<G�>II>*D�޿��#��=���7d�;(3�����FYC>�5n>$ކ>�̜=5��=Ӿ7�q��c���Chؼd*>�R�>��?b� ?�J?����;��i��ǩ�����)�>a�
>�y>�n��25��q���*�2N���A���z�X�Ŭ�>�1m=ڿ>`Y�=��ʽ��=��>	&8��۲������$�e�}<� �n�=X
�=�!�=C3t�?Uq�Keؿ����S��!S������zfK��d������8��s#%�	�s�����>sA>5Х>�h >Z�>!�I�Hf�UΎ��H�=���p��������w�я��k����ٓ��p��yK� 7���ν
�9�#�4
��:?��?��9">��>�)p��U>M�F?�;>?)�.?���=)?�þ�x�E>�]���.2?I�>?�#?��%?��(?�l�>������߾6�*Xx=OMۼk��;$G�=M�{=�1���O2>��|=���<̏��=��=�$\=|��= �=�b=U�=��=��,?C*�������pE������������>����V�%?K��,�+>V����|l%��.�z#`�>I�?i��>ML�>�ƾ)L[>�x��z7�!˽<Q/H<D@Լ_�;>�B�>}tϽ~:s>��'=5ݯ�3����JJ�)h�<$*=�Ȕ>=9!?7?��9?�e��"q�����ھ@w��_ͧ=���ݺ,�%>i�'��=��~�վMa7�f{)������Ȝ�F�j>g�>)E�=&\�>\�<�gW�!u�<S���
��zda�J?1>��N=`p)<h0c>��>H[,�WM�,jп]����ΒN�df9����=�Ƞ�0���#R�=�ľ����'�O�ޖ-�y��=
ӷ>[��>6�=�&�5����["߾��/>�V����4�-�.��}���⼈(k��r.=�t���;>�{H�@���Y3������M^R��@��R���� >�d(?3E=��?�oL?�7?��? �<��%?lԾ�?�nY���>8�?�=?>�-?�?���>t�3�_;��D���R=L����u�=o��=��=�2��n�=�RF�4-=��%��غPW��F$;���<$��=v>>�=��'?W6���nA��E���ľ�q��P�'>XX�>�)1�1Ȗ>䌛���=�a��%���(�Qz����>~X�><��>K@�>�FM>���{�c>�;�=d>h����<=�V�=[+�=�4�=��>s�i��g>3�T�EPr�jjK>��6>b^�>�x"?qi+?��>u��W2��LL�j��oIѾ�$�>`�>��?~�u������@�Z�	�H�VA�}B�=�d7�{ݮ>��۽$	��t�>������ =Z'>q���7轱���w��<�=L��9�>�����Y>��>�Ff���w��gܿ������;� ��F�髴;�糽��Ѿ�u��z�����$վ�N.�A+�>ˋ>�rY>����#C�����_�U�Z� ���J>��g�x	��i���{N��o.�bH�������w���+=����A�	<βa�J2뽟+d���`���i�+�g=җ?T�p����>R�M?a:?Aw�>t��>]�?�S�My�>�\��H?�%?a�D?%9?��>�>yΌ��ٽ�ڞR=�H��r�+<��>��p=��=�.>a<7�=���B���侼W�=B�=(P�=j6�=�B>��?W��=H�5>%�7�Xd�ؿ1�����O{5> ((�K�>>k��T�>��D����^����(��56��2)��p���>w̲>��{������/�������8>�/>ν3��Q֡=�*i��Gx�t5N��в=i�L����Ny��Ż�� )z>[�?�c?�b�>����7�Y���Fɾʓ(��ւ>y鳽.��>��e>����*�� �9�2�Ly1�ʍ����>n�>�"�=���=��<7~�=t�q<��>�
/>�|�>�$�>7�>�)J>��>�1S>���=m��=\F1��ֿs඿��
�*ܾ�X��	��n�����Tn�=��Z��U��*2پ�G>�>��=��?>O�m>Ϟ'>�0t>*惾YzZ�B��<pN��z=�_����=<��}�j���O��jC�g}���~����@������ｚ�1���������!�>M��>��A�nh$?'�P?\ZE?�2?�Z>W�.?!���5?
C*� �?��=^�? �?-�?��&?[��>�s$���<� ��=��=���=O�[>�8��Q�v�j>]Y��1��Q@]�Uy�=!_���D��T��,�=���=
�=R/�>S	>�+W��ݥ����K����×�XԔ=V��& �<])��	H��0���&�{\5��qݾ��j�6U�>���>�Y�>!�?u���mA�t�>�����s�+>%� >돀>B��<����=Qp�W������e׾g'K���]>C$�>)\�>?�?� 8?�'-?C���K#�-�$�}?��4�ž��>�Ճ>��>;)�'D.�Ae��F0���?�7�#⵽��=!��={fI>Ⱥ�=xL��u�>�>�>pO�=��
��!H��ђ=�F�>Sn�>���>٫>��>���=�߉�{$����+����� ]��������=�3���Mq�UN>����d���G=�`�>2%�=�_>�"�>`�>Y �>�0`�����#�}�����3ޑ�Ҿ����-̾�C�2�ʾ���)ea�E.��?�+n�>�r�W�6�,�q.���><_ο>`u>�]������62?�?�Z?���>N?�%�0��>�I�>�h�>(�?k�=?�q?[�?�+/>��H���߽I?��͂=�a>�kd=x�'>��>ܙ��*>�B��񚩽0³<�܂���N�pFJ��*@>�[�=~�$>�4�>���>��>[t���z���`۾�*��3����>��,��=[t��3��OYb����q���-�vM辀%�2�>�ֺ>�?�嫾�0콀�
=����«(>�fG=�
	�ڊz������SL�1B�t~�M�ڽ��i=៓��d���ٽ���>:S
?�uM?z��>����ن��,�t�*�ߨ�8ng>4
b�'^A=�-�=4�P�	�Ӿ���|��$����]j��)Y�ӛ>�1>Q�>$�>�8!�A^>��>�>hc^�$=]>l�@>�i�>|+j>A_\���<쬚=�1��(R��j��=�־x5-�~�I�޳��O�=�k���������ӧ��5O����K>&��>��>咙>s�>��>��>O�������:���:��D����+��=���",���\�x�*��X��i�����Aν���_S#���,��8
�ޱν�M�>�+;�R\�C�a>�`0?ڪG?5W?�#�>�-?@ْ�yp�>��[>�#�>.��>M�?e�3?x�"?���>Z��ԃ��Խ&>Żq �<k�˽F��<��@>4S��@�=j�<S><��D�ؽ=z��`�O��I�=��2>Ca�=מ�=�
>c�㩾;�=��?�����!Xu���>�н�>@3f���2��Ϛ�����B��I��<3ZF���&���="��>���>]v��Q�Y�J��<�w��m�=�G>�ѭ����nED=߹>�u�tn{>Rq�>�|ҽ�뎾.�J����YF�>A=?��d?	�>���=7�����������7������E�>X��5Ҿ�	����D�N$���2�h6�������"�H�'>5�>�C>�_>��;���c�>�-�&�r��J�<uԭ>U�>b-�=�j���Qr>�ː=�c=��߿-���|E�ʗ|��r��kb=a�d�?*���ϰ>k��>�M{��O��5ʇ>.Ǟ>�2i�Y>>��>�3<>5��=̻ξ���C|v�kB�;���(*�������I�>Կ=����"���S�/�q��^����N�K{1=�-��`c���Y�>b�=C�f���ѽ���>wu?d1?LY�1�\>�E�ж�>q�<@J3>���>i�?��>���>�v�>���=4H���!̽�=��=�}y=��=���=��W��_\�=�a>A�½+����r���ܽJ�=1b����P>F�=�>%?�`?�D�����,�^��_���b?S�x7�>�r���>>F��t]�`�]�԰��$����"B뽧xn>�<�>�׾����.�=Eg>�1=䤅>Wԑ<mu���Fq��_4�y���������=�R=�Ī��8a����k�>��?kR�?�>??=��nf��)�Ǹo���J�>�>z���9�����</G���;* ;��T{���F�N��<���� �>ՙ->E�7>��=��i>㟭�9��=�R>�����=���>�[B>�N�<{��=��H>uW�fG����ҿY?���8I��r�ub����Vzx=�+���=�T��!f��\!>�N>IwĽ��]=� �=��=I�>�-�>c�K�ք���4}=�z��ʹ���z�Mٙ��c��^���t{��\ýS7/���u�ƕd��^��Mݽ�Ê�l�ս�6��>�2��Qݾ���<>0_?�g?�J?|��>+�5?��=�y>%y����>yT	?��>��>N�<?��"?���>n��i:����<�N>�M=M�ż�����8�<�>�h=$4�=n�=�$c=<��=�:�x��?�?����=+W>:?Y��=���$�I�":��^���1E���?q��=, t>Vی��"0>����F���DTɾ�Y��[u�>p��> P�>��r>�௾�؉���n>ZSY�?��<�>�b̽}\	>�)(�of�>C�I>�."�R��h�Q���;����=�o�>�(??�??v��>:S��us��/c/��Q�ժ	�nx�=�d�n�<˝�=�I׽0�8(����7G��L��ن]�8��=�>�'�=k ��<^>��<#�!���$>�����E�=�q=�����P\�=t�f>v$�>�!ݺ�(��m��)]ݿ�괿jt-�<S��>�e�=m>{�J�v�����'�z>��������6�>�
�>�9�>X�=�a�>sr|>�,�#M��K�V���E鳾�呾��۾���M���w��:�Z͟=
J��3������)۩�T2
��Y]�q�`���3>�>Sх=�*O=7?�,E?�`@?��=��?�����=>sؽG�>���>�5?�3?�.?a�>{0���B�1ȥ�Zh�=A�V>�=�">Oυ>%�ɽK�>R	=�lL>Slg������=R�߼f��=o�=KM�>s�>��>c`>.�ξ��;��!Z*�;�Ѿf�?_���=_�:����7
�0k]����=�@m¾#f���$��G���ܗ>�č>����۬��1HJ>�ٿ�܀�>̀�=��p�0TO=���;��=;&+=Rq�=�j��_�p>>/4>�y}->�->
&?�?k8>?�-��p�#��Z��x� ��P�7�H���`�G���Fs��#�~p�����Q1�|�c�!��Y�=Z�N>�Bi���>�܃>���<�=C�4<�y=�><4�n�@r>.�>���`!>�E>7Ľ�1ӿ�\��x��ž��7o�z�^>��,���B�f ��Z���rn�>L��� ��o"�<��H>2���J�Gd��%���o�z���o�5>M�=n��6�ǽD���c\�Ԋ �����gv����r<�ۿ��L����A�� ��ǳ��?a��↾���>���>��>�&5����>���>��?����tTZ>=��>�V�>A��>��?�s�>(i>N�(?m?�?�z�>#)i������h�=6D'=w�����,@��@.w=�u�>P��fE�=�½b��<�Ȧ��
v<h����к;��O=9�?=b��>��>\���d ;��A��踾���`�>�R'�C�c�q����uJ��[7��e�h 4���++��/��(g�0�>E��>˾������>@ὼ��N��>��$��1��f�ֽjݙ��o�>ZT>����|̵�Q$>�W=����!@>J�#?���>4�*?5|�s�9���˾}���y����Ƚ7��=w�;U)G>Y������Ǿ�{۾U�*�4��������.=�����^�8�=c�7=/�缉�K�Srl>^Cn>�;>�`r>���uG��N�$>�>�qn=�	�=�98>l��i¿�M6�l���8=߮�>��=������	�y"	?�b��6�۾]a1�pY�=A�7?�ف>~ƽ�c��걆��Fͽjn]��r>�/>��Ӿ����iIN��6K�����sû����ߠ�����I��B+=�H��3}�U�6�������>O�Q>��="��=�5?�x?��>F`Ƽ]�>N���J>��>+M�>KY�=D�J=�Y>Β�>@�>;]�>��`��EW�&m�>�s>��<���=���=(�̪>QN>e��==���y�:�M�$0���=���05��H<Z�=f���T��=�r<��=�I�s��h��/�>>��i�>�֓����=���j��FǾց=��3�I�b>1���#�>i��>����m�I�l�ͅϾ�B����?=
��<����D�>͕d=���=�ӥ="�a>~�M���Ⱦ��5�
��.�>�D?���>��?��R��b�E�3
�c�M�+��q�.>7�>�n׾�I�x���q�ӀU���O��T�o���=�o��mg�?�>*�=�J>	 >�4�=��C��J�����P�C�o>�ia>�b�=��{>�*��B�=oMٿ�Ѩ��rC��۾ܝ���"v>����|PC>���>ϑ�dc�{���e�>�Hս�����>���>y��>��O����㒷���^=��t=Mt;;���鎝�d/���=-�=�7��L��<����&�c�HԌ�k]�_Lt;��=�wm�y�?_|>�B�2�p��F6?�<?o�+?�c+�����!>� �>���=l�>��1?m0O?8�?�R?`�>4�?CI$�� 	��	5>Ҽ>8�8=k>��ʼtk%�4->���*��F��#>2R���/�[�O=Y�<�es=m�=«�>=>
`���*���0�,/���c(�p�?+�>������yC��s�%����P-���>�־$����ı�_<4>��B>Z�ǾD�W����=������>>�n�=�����_A�ꍝ�+棽�$��L�=a1��kp�<��/=z�D�k2~>0�~>�)0?��?��O?l��2�%V������������h7>|
8���>	����b2��E%�ju�L+"���f�$o�C�=�{��a� iH>l�5==
��w�=�e���&�=R��>" �=1��>�Z�>ۓ�>w䡽�z{�#f>p):�=ӿ�"��<^��p3����:��>��|��ژ���@�AFK>��N�d��=e�>�ʵ��Q�<�n����ź�U�>mq@>�>�	���Om>*�[=Q��d�<mG��4쬽%���=�m*�4�p��L.�;��GF�4�彾���A�l���ʾ���>8�>É�Q��:��_?��?�M?\�#���ػ�E~>B�>^]?n��>õ ?o��>V7?��D?�"�>���>��tJW��a�>]ڌ=*þ=��L>���=NA�"��>�О=�y�W��=��=+S�����<>��N>\��=�A�;���>R`>�-ƾ#X2�E�>��@�*����?z\�g=�����a��9`�E[��E;��f�y:��^JI��R��>���>��m�p���3=ysY����=��>�!�;u!�I��=�O(�������(�T�;��%��HT=��ͽOƎ��6�>��>?�X1?s�Q?gD���$8��Z+�U���8���`� r��P���C���^(�F+ؾ��F��E���E�x{����7�׀>�b�=격=��T=��7=tw���=��>�>4s!=	~�>Н�>B��;��$>
WW=nHd=���=��ƿ�ͧ�_'þ�c&�5���A�>x
J>;C=�B�>h��=k>��O|�=$�!>/��>"�>�î=t�i>ӊ/>�r�>Ə���L��X
=Hه��x����;��Z6��8&�ռ����=�h���⏽��!��0�<�K�_ ����w�y,�4��>��>�Ƈ>]�">�_�=\�k?�-?���>����t������>�&(?�E	?��?p^�>�,>7#?�5?�E?�C�>p!P�?C1��w�>�>��3>��>�:��K2����=�5��{W�����=8�K�˽[>v��=lO�=��
>�'>5�>�Gn��}�����0��þ����i�>K/A���>��½0�{[�?� ��)'�'���Ӿi��>���>��>+�>4���>�f�=�dU�,�ri�<v?�=̌˽5G?��4�=S/=���4���iӺ�W<�@�;a<;~v>�1?�[�>,?�O���%���)3;���=���>��J=Ѯ��i�����p;�>ĝ�͜3�)4��۽1�=um>��l>��=q�e:C�>�>���8K=�Ak=�Y>l�>˔>���>@��>���=�d�<�?�r�[�������h>��N��|Y�Z�}>ŵ�<�O>5����A�vX*��,�R� ������'�=Q�>�!=�_�>��>���q��d�����>^}7��è���=� 辦w�:��#�J)���x㾼a��񃠾=zl�"�;��?�Qo���T���;��>A�>n���5�>T�?��>�\?N����&�>JGҾ^���^�>s]�>�9?b%?�r�>�~�>�ST��� � ���Ȑ2���L�Ӽ9"��Ux�=�^_>K�=�1n��L�=la�=}���u�Լ�UB�ǩy��""=3�=� �>�{n>��+�����h뾴I1�G��B�̾,G>��2?�㾊�$<�2���TH�-�̜������Dc�=�u�>�E~>���>ƞ�>�fĽ���<�#;�6�19������ǥ�L�>��=!�a<������W=��� W��~舾�Tq���:����>h� ?��?q?<_\�	���� ����h�r�D�����Q>��׻|b\<��@��a�bӾ�%�{��1��HV�\d|>h��=���=��=S�>�p�M�^���>��.�|s=�fU���:>�/�=��>?��=W�b�� A���="�ٿ�+���%���+��"���ʢ���>K�#>��?�����ƺX���	�n�=��y�JB���7n>�e�>�G�>j��>�aǾC�x��G��鎾�7������][�8�7=<3�!�6���߁��2E�^�+M���U�&��<`7��3ʽ��>�o�>��=��q>
??��?O�`>CJ�S
?�
={>!^�=��>���>��?�@�>X��>/�=��>���C	���L�?B=�C,=��z�E<>�GZ>vq��@>�~z>GCv>Q8�<��
�=���(>�3�>|T�>���==�=>�{���_����P����HI�	3�pG�>3e�Ԯ�>�=���|���:��lN���DS=�Č=��>�~=(G�>���>�6���{Ǿ�wX<c�ټOf㽌�>Dg��`>y%>�o��Be=ţ�=g�1;�}�[��=Ҝb>���t>!�%?�D ?�n?f������Ü>�=
��}">���01�>Nm�>��=�R�I�*��"�ޞZ� pԾ��%���=Ye>}C>��=�s�>���=_-:�n1�>=����Ƀ����=t�k>I'>/f>���<m���Qѽ�~B>�8�'B�����V��z�Ӿ�&���9d>�/S>��2=>'��L��=�D=ȍ�<�2�<�E5�~��=��S����=w��>����}+��p=:𪼍�?����倾哳������9`���c��0(�����\�����
���6��۔��ln�<�?���>�OS��=&q?C�>'��>&�$�5�>�X?�J͊<u/4=���<��>�?�ʕ>�Z�>�u�>vg=g�����B��l�=I3>��|;�[Z��)�=L��=K�=?ή�~��=�N=���L����<��=�G=X'/=qi=�>���j�Z��X��.��4��{�?-���-�=�����4���e��h���?�=�E!>���&!��νQ�>��>���#�c�|�y>��<բ�8�>�+y�Y:���H=֎�=B��=L���={ �=M`&���I=����vBl>�?��&?�]�>����A�B�\�Mz��N��)�>Y�>�>�O>�8��5 ���Q��#��(��SX�<p�<�]�=ϐ =㰅=���<ql��9ݼo<��>9�3=�.�=�*>�8�=j�Q>n�@���ܽ��=@f�;$���#���ї�?n���n�+v��r� >��>�:=�U�=�h���EY��ʾZľ��<UO��2�=C?�=�=w��>z���8���}�=��۽N���H���o��=�����ռ�}���^�끧�Lᕾ-���U�C��pɾ�����|�0��>.Q ?�n=�K	?A;?O�/?���>�ے�Ӑ�>�ƾ[��=��>��>�L4?DZ�>���>Q	?���>��	��fF�j�Ľ��f>�^>P1��D�>�/�>my]�i�>Fw>"T�=���O�x=?P=�ļc��<��m>�;>�A�>!o���վ��;N�����O/[>m4>D
?���^���Bwʾ��羵�B>�}�������<��.>��>�t?= ��>_�>౽<�����=���Ϝ�/s�=�0��)QE>sP������$t==6������V*��;w�^�=�5ȽK�v>�?���>%��>������<jL�P� �M�!��?Fv7>Ao\>r⽒����x�ʚ�B�7��WA�{v1��V����>� >֜l=Ο�=/{<x��=m<9&/>|�^��l�<R�$=��V�{3=��>�l>�>?�C<�z �5|޿�������iE�6h��1Y~���`>#ϲ=U>�~�^W������<8�H=��W� �>��>�S>��`>\߆��6��	���9���羝�>���Ž1-��b�n6:�F� �b��=%c�﮾�\����<da=�q�<��	��?���>�hv>j�m>��?�#R>�r>?`��@�>%�&�)�>1��>�Xӽ�r$?*k?��?zWY>a{�=��żދ@�U-���=l̲=�_.��>�5>��'��UX>�ܱ=�[=����v�;>(�(>X�ݽ��}<i>6i�=��V>��?��=f����1g=�@>�y�ﾎeƽ���>��ʾϊ>��_����͢��׾��G-�Z�>�a�><Ű>魋>�j>�;X>�R���b��y�<L������=Fz>ݨ�=�&^=��r=[+V�� �=���=1��=�����O�=��/>�z�=�=�?��?o��>�>>㭒��s#�����kԼ�~:4��>�O�>���=�i�M�ժ?��(A�,����\��ֽs�=H�>��=��==5i=�Ȁ=�oO�:_���'�G�l�H3�>�L��a���ߠl=U֠="<���95�t�����H���G'��Z����d>�͊>H�{>�V<�m>_pr��lὄ�=�
�>���>���>ޱL>'�8���>Ka�=�`%��p=3>nW����&t����̾$�i�I/!���j��'w<9Zd�Nj��eT��yH�����w��~��N R><>Pa>��p�0�?�Z?��
?�B�d�>x���Cܼ��w>[p�>�a�>�N�>~�q>\�A>���<<;X�&��_d����>�g=�g�=�;�>&�4=�o=o��L�=�ǣ=ʲ �&��=���=�l��J�=2'!>`kE>upM>L��>����,��{��AH��0~߽ym��26�>����������d�>賽��>/�=]f=P� >�+>,]#>�1I>��j>�QɾN���.b=�2�=�U]��
�<�=03+��r�;�ֽI��zZ=�v>��=��T>��R=߾9>���<�-?��,?� ?H�=�d���X9�>���:���Y�=�f=>�M��ཊ��B����B�������n�e�d�P�ѽ�}>���=��`>�F=�,����=Ht8=��=%�<><s+>:>͆=�f�=x�=Ct�'��1Dm�ptӿ뇿3�<�@��=�D�=П�=�8&��냽��[>\�k=��������S��ﯰ�W�=(7�CoN���?�KL�=�o�=w:*>K��:&���`ɾmҾ��:=$��,٢=6꙾�p�A0���_V�������X��A����'=	�.W`>v�$>>�3�>1[�>��>��>�Lƽ�P>�n��,q>s�>�8�>�H1>��~>�>�w>>K��=#i�kå�~w>�=��/�UV�=i5�>��½ŭ�=�s>2A�=��D=?��=�*=��X<*1��
�Y1$=8:&��H?����¥��i��=�ۯ�����mh�í�[f�<Π=��h>�=">���=��L�]�M>,J�H�����f�%��>!'z>4�ʾW��=Q�I<Gp>���{R<fu����L��=`�<R�=�y�x�����l>��H>j0�=.�r�
?>��G?ܕ�>�M?�|��T7�����$�����6��<:7��܀=N9� ���$�����❾Eҽ�&����<�"�>�.潗yT>�d%�W0��M{[���>�^>ԑ�<O�=���׋���P>p3�h��o�b��M��̿�R���X>����>��>�ߘ>7��;�l>o��=y���ep9�Q>�����=^�>���=� ���B>�4y>��:���<��1>G<��"T���&n�}i5��,��HB�ȽC�@��D�NOw�����(V�XD(�mh��^Ӝ������<>.��>��>K>�r??�%!?�?� ?�y�>�{ �7 
>�M�A+=�CY=oF>`���ܔ�>�}�<�V��	 ��l6���>ͻfD='�=:��>?0>k�>>��>��"�^����>{\>ga>*-�Dl6>�]{>���=O�?b�޽k� �gV�������c���L>���U��tAE>O'N>���>��>�ʀ��ݝ>G�y>y߀��Ӥ����<��>Ǒ�ɠ*>I�0��-�<J����Q2��<��څ=	<{F�=�S_�_�����>Ɏ%>�4>NŦ=EE�<]��>�4�>ڼ�>jM?� 쾸�6�ƸH�-�4�|1x����>Ԏ�>>��>��u>�ǾC��x�k��
��Q-�O0>�����0 ��!/>˴���>3���q�_V�=B�=�+&��"/>Կ��fT>!;b="Bx>���.Q<F{һ� �wɿ�B����>.2�g�>Rܠ:@�>$q���>�>�⊼�0�m�}��J�-b>>�>/>��ħ�ǘd>C,m�zގ>�a��l=k~V�:���\o��^����zŽ��P��7�9ی!�b��#����Y�\�h�4����Wz�`!ｄ���`z>��??[�>���>fZ;?�� ?��$?}:>?��>e��X�X ������ڬ����>mP��L��>�I�>$�)>�Ԑ�o����>>��d�>�e>��X>�g>-(�=��[>�,��ײ��:+=31�=s��=��,������	��a��
�=@�>-O��Wھ�ƾ����5о��|����*���-D�=���u�=��?>*%�>֨���>>�Ԁ=��0>B9.=�g>(d�=��7���� �A��=��O�1���
�����=���=���<V����=�>���=8�=�f:,v=�<X>���>T��>�"?��D���0�O��-~��A��r�>2��>Ճz>���>��Ӿ�-����)7۾�	.�-�`ኾ{�<��1>�I�=Б�>0���g�>�*l��df>�J'>'=��=�k�=6�X�H?j>wj=	����=�cټ�п�����M�>�b��>y>�2�>�[ĽX�&>j�>�[���\��s˰��Ց��S�:�><�Lq�����=���>u�T��HA>���=��UN��*������|U�S���>y�|O�i�<�&�*�Z���H��b�9,��?�ؽ�:�>�o?;T;�^>ɱ)?��>#(�>��7>H3�>lL���y�;U���U���m�X��=m���-�>�l5>��{�o��,ع��ǖ>�mG>ĩC>d@>R�=b_�>\A>�ZA�_5=$��<Ȋ=X�����v��5ǽ�d�=��"����t�>�!�>�(�������)�hL���}��8��>���>f��=�1q��ʾ���v��}$���>rk>�W>���=���>��>�`>��J=.o����qC=J�R>Z�	� z�=kQ)=���Hǘ����ô?����>��ý�V�>h�>���=�%?L�X?v�p>�N�)����b�tHW�]���C��>�Z)?
���>g�p>��&�?D[��nP�zf���%&>�2\>����k���*3>�O�/��R&;}�>�m<��_=�>���>	�>��>|
>uT�<i�(�����8$��i���\��<�T�7>[L�=�%��1ǽ�P��q���2�����{���ü���=�<>�X�=�?����*}"�Ǹ�<)�$����� �o�����|HI�$��lֽ�˽���q���g\��Z����S�����]�X���n�>{�@��I,��z�>�OW?R'?��8?�s�>���=��X�%���X��>8�$�.>?'.�>�n�>8��>��>y��f~n��.�ѐD=�h�=�'>B;%>c:*�@���qżH�������K����=�Iٻ	���Q�;�j�>���X�>��=��O=����n�-�FNj�R�ɾn��>�_�����>敥>�i���ײ�c���G��5�Q��T��O1�y{(���>�A?��ҽ!ɶ=ހ������
4�j�1��7,�"���N>�Z<�\>=\�;G����ʽ�	>8#.>9�9>OS�>,?�>��"?Y�Ҿj�e��[����L�>��<�,�>�u+?�Z/<Q��s8��M�7�#B7� ]=�l%���"=#�.>sg/=Fn��gSH>�!>��=�D5>puY>El��x�ýs�=�N�=&�C>��>�~�>ç�=��=fQٽ?ٿ���)ھ�W��7콦�6>{�A>��b���m�PD=�`���Lν���ͷʾ��ý!t1���R�J�i�3�=�Ⱦ�~���a=
���I�ӈ�_������A����=�P%=vK2�ٜξ�V������������r�V�X��Op>��%=Ә�=�!v>�<?��?�'?Ե[<V}D>~�����
�%�>�>;?���>c(?v?3?���>mǽ�{���j�;>�m=b�6>�p�=M�%>�P�Ĭ=�^=s~���O=Vb:=�м>���C��"x<�6ҽ�:�<`�$=�W�Ǻ-�$�2��Q�0ƾ�����$�>ƞ���N>Q=��m��Ql�d;����Cž^7�����%���8��> �?T�==s?=Ɂ������&q���9�������`�,i�>!<����+�%��籾wނ��3�D^��<�>�G�>��7?EO�>l�=I�Ԗ�ܾD�J��zdݽO�[;�>H�?>����8���򾸰2�� c�P�e�T� �D=��>�uL<���;D >^5>50>�8>/�/>���qټ0r=�9>�!F>���>O�>�/>V>-����#׿%ԭ�r7�p�.�=��>��<�K�����=�_�=U	�(P1��)�>}
�=y2m����_̀>u��=P�#���ƾ��ƾ=����P�����!��Y�x#�����U�=�FV�\�ǽI�<����Lt�����]�]�Ľ�9�����>�{%>�̀=��>w?]@�>,L??������">EP���꼔T>[4>{�?�6?{>?�?[�?�7�>|�㽰Um�x)B�X�<���>��$>�?�>�k�H´=���=n1�����,л'aM�e��iI�7O=��=`h�=��|>��p���\�⡓�s��w$K�2�����ƾ_�#>*�r>+=[�.4߾�p��|����XѾ�;>�zi��RU����>@;�>�ھ�����¾tӘ�����|��~ƕ=�T>w0�=��{>΢�=&���m��Yξ*{
�7��|�<���>�%?�Ӕ>��>s���7$��M�/U��L ���g<��>Vo>>�ɽ�7������=�T���D�U����=y��=��>��V����=|L�=D�8�19�>��R>��Ľ�<@�W=~�>Ru�>�x�>���>�[X>�^s=>�I��3�?୿�%���C����Ù��M��<��=<z�=
�>�V�=�-
��N �(�'��jW<#	�=2��=��5��ٽI3����!>�%�&�ľF��͚Ͼ5��0&˾:.H��9�a3��%�N�Ç���d��'���#��i���W��Ƃ>3|�=�=��>)]!? `�>L�?B#->zP�>,���žj��=�>�?�?��?r�>��	?fһ>����th�ґ�=z�1>��>�=<>1��>�X�����9�<*"�������?��<7�6=Rw�=S�S>�f>j9>��>u >LR��z���C��$.��캾�b�=��r��0]=��=��p���ξ�Ͼ%t�䗭�}�G6�����jg�>Z�>?:���u�<.|W�(	��>��T@�x��>l����:W=j�>>�x���T%��%������=�2>9�&��j�>�B?_�=h\ >�̺��'O��+?�z�����������87>z�?Д#>V@!�y�����C8��0�\�����=8S�>��<�FW��5�=�1>�S����H�5H,���=3��=�x=�{>�n!>ω�>[dZ>��U=�n@�4�<��ݿ*����\�=|��h֩����=D�6�B�^>|k���>�\H>�m�o�=jWm�*�}�
�=��g��C1i�|
���5�i��>�x��L��M�l��8>zT(�������н	է����.��x龱�ͽO,���E�Z����*�>O���m���>��(?���>(T)?,Ӡ=���>��=�ԋ�Yt����=s�?�?���>��	?o�?.��>����2���3g<��=`�>�E=��>��2=�����%X�� ����T<&�&�"k�<Ǒ�=���;�P�n�]��3>W�>ɛI����_'���*4���ݾ�f{�R��>>]>^>�Қ���w�V�)��d ��������f9þ��d�g{a>���>b?�Wp��O�cVG���g��nJ�9�>�P>�?�=��<�^>��U=� �i\��n�.�U��x�<B�M>R��>S�+?�?���>X�Q���پ�5=�7>�kؾ���=I�>0=O0>��پ��!�.�P�3��P�4���w+�=�/�=�׎<�:f`�>�J�=�a�묦�8A��>�9����>�_���%>���>%�>��a>��>�g˽�ߵ�V���W\���\��$>���l�?S>�E?>�����]<�t+=��� A��v����j>�M�>���>��]>�C2>0RK>a�վc��d���� ��U��?:�
k����p�߽�$�;>�"��6u���о��Ľu=�d��N�����
��	��q�>0��>o7�>h�>��M?��>��>f%N��c�=��}�0�>0�?jH!?�?���>��!>�+?W��>e˽�Lƽr񇾟��=��= 2
>�3>���>�$�>�>)�<�$���=5�>W�>谤<��>�.�=��=E�">4��>�|>�=�:��q/O�8������@�>E�r�jmT>��>���f��.h"�ba��������6mH�:䀾�}�>�L�>��^�� ��~L�=�����o=���>��]����=>!��-]2=��1=6�a�b={B����=�=C>��=)�>�7?;�I?%��>lf�����{?�����UǾap�=ƕ*>����R��2���0�P�?�)�E��hS�(}ξ�D�=#��>��޽@ŽyL�=��X��?��Q����3`���=�_p=�\�=�㉽ߦ$=���=x�>��">_D|�Q����տx�����f���t���=_�}=�_�=$2�������=�����=�L?�ʘ>�52�K�1<z�(>�c>J����\��)VX>�������m�=�����|=m5��`�������o��W���<
���k��)�����YG��j�>�>8�'��!�>�dV?A��>W�(?����>��+u��`�=>46�=OC�>��?c�7?F�6?���>i$q>Jٲ�p,x���y=qz}>��>�b�=;�>#8��IR=A��F=�ʂ=��<#��=�`�=X�"=A�d:S33��=~�>��j=�D�> 9��;#���^�q5��c�?��k�;�|�W�h���>m'���"�)o��膾G���=q�М�a�>�\?7���X���i�I�f
~�vx��*�H��|�>��^>��1>҈�=��t��`��0R$�-�P> �ս��P>��F>���>#�X?��?��>��)�5�5�X��h��MV���>z�6=;f�L؊>��,�"'�wG��?�e>N��M��'̽�g�=�b=�~>��=��>�t��>��=�2)��f�W��=������/��>��?!�=a/�>- H�;����ڿ�VӘ��G���^��&$�=m�F=ܵ�=�c,�_�پ�-1���4����>i0�>?��=O  �ڽV���>��>�ڽ��P�_�|>�������7<����	a>5ҽ�?���F��G�����}h��OZ��F���>�[ug������>���=���7w�>�n.?47�>��*?�g��`�>&U�>���>vM�=X����E�>�?�$?H} ?���>���=Z��	��V��<���=��K>N>�:�=]ɮ�R^���r��[j����<�D�=��-=UO½&Ky���@���=���=�g�>��>Su/=Y���m�.��<�;��R��?���~����PA���ݾ_?�9BB�dA0:'$r�|�;,#�=��>���>���o�_�=V���J��P`y>A;ӽ >�u>���=��V�J�!�����>����V+�5��>���>bG0?�G?.O7?��r�����d���۾c�۾;1�<J�=���=��>�����=��-�_3�x�3��p���5=�ޛ>Y�w�c�w�M������	�=F��c��=k=�&�=hA0>�*]>��>b�>�����y>��:>܂������xP��]�1���"��p���J����=�nپm���
$>M��>�E>���>i' ?b>�>Y>>��>���)�I�7���ޑ���k=�;h�Q�Zy缱�j�lļyO$�\#%�u�$�>���8x�ɍ�R����6��w��\uc��[�;��>��a>�W&���N>v?��?��I?�>��4?�V���<���o�U~����6=5��>{�>�?��#?�&?�����B��=�c>X�	>x�=��B>����4��=�e~Ž ��hݼC��=�^H���q=Q��=cd-=�[T�7��=[d�#Y4��2���Wᾎ���$���N�>+�żh����z�=t��67��2���B�=:�=�"��s���z%����>�=\>o?<>�߼M����N�t*��{�=se=���=���>�(f�h�Q=�@�= >�C=��,>_i�=bf�>��B?s:K?M��>��Ծ��2�1�_���ξK	5�nrR=��>��e>o"6�7b��!�����S 8���8��%�zU�<��>��=�'�9�����%�j0U=&�Ǽ[�h=���<�b��:�}�sT~>�֠=��>=�����=34�< �2�dWڿp���I��x���H(�V<=�V:>��̽3쾥8��D�F������0H�_�5>��=�Tk>�e�=�^�=|f`>N�V�t�����=
 A=N(5���=�����-k�=L|�_���н{E����_�FL��d܁�IT��Se[��ֹ��D���>TŌ=�@�;�->�Z,?_��>$�&?����Ǹ>D[I>ß���O>F�#?T)$>��>�0=>8_�>�R�>���>�j��o��9����;5XJ>d�=?*�=��ν��
�������/>�-�=���Q���?�3֧�G�޽D�	��=�=0f�>��X>�/Ծ~p�F�.����̼�>�m����T>џ�<'b)�Wu�,2z��>>�5>|�F>��T>��Ľ8-�>6�>����.E0�c�8� (��"e>[�5�L=ot1=!��>��켊���Ň���0=3=lνV�?>Ț�>�!�>�;?p��>��?R�˾?��^�L�15�����X�>i��;j�'>b��>�F��J-�;f�-Y>��>�^Y��f����'�=�ܱ=9B�<��>�=\�=/�b>�V�=���8H=�#�" d>�&�>�$z>r�=��>�A¼p����ο������r=Īξ%7�=H�=�p<�^��=k�!��IG�d��ǟ!��an>�ѽ=���<�=�r�=nV󽱍�>2
��ۘ�>�㊽�󍾌|��U����|��UT>J����T=׋=s>���W� <��������ھ�iO>�� >�<ۘ�>�bS?/d1?2�B?ɦ>��+?]G����>�=��=�|?
�>J��>���>Y9�>�z�>�ێ��$��>M>>�q�=��>z�W=�	���-=?�@��+���`�<�V���ɢ<�j �D&=��8�	�t=/�	>qW�>�$�=+}���}k���7�Cڵ�wE���:�>�+��Ǒ�>�s�cP�{Ž�៾�<=?�W�Lnǽ�f�T�6�q,>DU�>���锚='���ã���>�>ޮ�z��=P��U�>�u��l��=��=�($��|>��=�I=���=_��>�M?�j�>���>�����/�oK�#���~z����Av�>�
�>>h >��	��kξ�"�7��Z9��v����jz\>��{=H!��r+I>����^�=9�t>cd<=F`�F��=+>y=���=��>��$>�3�<^y>u����)���ԿLw���{>4��p�=�A>���<��g��3Y�����&�
Ç>~�D��_=�M�ٽQ��N|����=���؞�>��+��<�>�LU��I��'����w���=�Z]��X�=���87>pN���ɼ�}>Ǖ`�Fߤ���j�c;�I�!>�+�>kgV�S�u>(T<?B�?S*?/E4��Y:??N�&ۺ>��V�J�=�? ��>��>ʏ?Cx�>�i	?�I���L�������F�A��>׶$>V�!����xu<�9#=Lw���=�䯽 �>z� d<��<��>�f}>���>M��t������I��T���{�����>$�ܾ�y">6���bt���ӾI�޾�鋽^������q��
o�錞>4��>�$ľP�ۼV���nFN��)�>��F�ֻ>c�h>{a=�oI��Ac~>��m>�K�=��#>��*>�"�>�zu=���>Z�?���>�0�>�,�(=��kb������[&��ʧ=u�`>�C�>��<����c�<t�e�N���>�?2��=b=��>�'E���R��W>�����?"�>w��(V��:D>Q��=�ֆ�}�<��;>~75�^��=5�e��T|��^Կ]����Q�O�Ծ~�/>��>��O=�O�=j}���d>\�	�W�ϼ�>�*�<�Mh���
�N��= �=<h�>��*����'�>�0������~=�l���<>eO��E��=6@׽�z���	��g�Q�,�������79r�׉K����>2��>��e�>��?�ؾ>*P9?ᷠ��6?�h��֗�>6܄��f�=��$?�e?.?�*!?�?�[�>��@�����H�;>�c>k�>��4>s��;�{	�5�>�ӽ��s��	=a�y=H?�@���͇��ĈW�gG7��tT>�X?�2m>K�¾\��w�	�xா�X�UN ?�þ�d�i���B���:�/����V��UM����+�{��	��>�(�>������5;&�� ν*�D> H>�!>fe+���v>� =yC̽A(l>��>*XS>6en>�� >�o�?G�>4�?�?D��>͒����,n�G�Ӿ����>_BQ<
f�>s�=7����+��V��X}J�v�P�^} �#ȃ=[R�>�+��e�F��T>�����~���=f��=�Y�˥/�X��ύ�Hom��E<�V�ǌ�<��?<�v��38Ͽ���[���� '��k�< ��<=7վ�,���=�#��\�=X�?F�>���=^��=��=��8��i��G�S�@��]t>�l�$k߾����
��>4�u*��7��=ƶJ�����z�>�\�T��?�$3��/�Ҿ�n~����>,gK>5�=��>��/?�$?�2?rF�<�=?C�R�J��>����y�����>���>M�	?�*?Yv?��>�8 �U���.,>W6
>� !>���>��[>�8�\h:;T�ӝW�a<=I~>A�;���o�;����%�=�6> ��>����Ԛ�񜑾j�������|>�@P�X�'��Ö��(~���p��끾b37�##w����ͦ�<}W=�>ʘy>�g�( � 1�;_u=��������2����>=t�=��=���=��ռa���h�g^|��75�-r��Nq>�>Z�?X�?�H���ž�0��.��9��1�>;�<�Y��N�=�NԾ��W����&��
��R���H=g>�u���	���>�ɶ����+�>77=�Z�4*k=z����x=Q�+���A>on ��Ƙ����<����ܿ(���� �U��?�+>�=���>�{'����<I��<����vS ��l<�>���=&��=x��>�i�=u�>ܷ�^o�J��=%�<#޾�J����㨽�F���|>�����˼�&�;�;���%A��d_�Nԣ�5i���1Y����>�p�>�;Q�A�#�'4?%��>���>X��>,p?��:��>��>p�;Z�?ǁ?9�?�*?�>;�\=�?_�L7|��s>_c>�\x��p�=j��>'Ħ���~>�|�=���=��:��$���>�
�cAi>=��>�2X>�ޗ>#�?���=�&��E��ˀR�P���Ԃ?���~����>����{�^�la�*T0���5�c�*�^�*��!?�[�>G
�>�]���<7a��Ϯh������z��J�!��'>�#f�#�@�;�$��[�<چ�f��Xn��LR<:��>/�W?�o�>�I?�����;���f��u$�[�=��[%� �=f��=®��ѓ"����5Ծ
j�Z�8�rvG��TӽY�A>U'>4\�NMc>�=4�>��=d��>/��ư<:��>��>���>�vp>a��>ތm>���=�i]� 3ѿ4碿�g����"�bY.>
lk>3M>�J=�TT��O�݋�]�r�[t��u�v��/x>�ڙ>�ׯ�w1n�.�=;� ��`�N�6>׹������*�R�� �=�S7��1�<��#�}Mѽ��ʽ�5ؽ�m �ŭ��p[�&����	2�>�1I>�ٛ>�љ>��?p]?J.?p۝����>���>�������>�w?��,?6s?���>P5? ?3˃��(˽��N�h5�=m<� >[>I�=
>��S��w>�୼�$���?Ի�K�<���t����
>��>+>��>���<�>�������{��ɾ ̍>d���������z!>>h@��*��78 �ܾ]����=�1�>^F�>�6�>���u�� �/��Nϼ�����s��>�~���,�=�W����B�j��OR����ۻ��_=r��>⍪>�q+?f=�=T+?�Wu�I�	�������f*� V���p>�
>���=������p�!5��xN��ef�{�n�+�=�B>W��=-uG>z�=_e->p�n=<�����k�=����{>���>��>���>]��>�X��w�ݾ@�ҿ�����ý���3;�>=^�>�ā�{��F�ʾ�.3>a����-��¬=�I�> �>H:>�8(>����6ѽ�R�>�s��f�>* :>F�q����I�[������m���t����i`�=�5ٽD����R���J��a�֬þ�w��Kf>��>�U�>�E�<�*�>z2/>'!/?�;�>�`�>�s�>�:�=���
/�>�?�7?ɵ?kJ ?%�>n/&�Q�ξ�|�UD>\�b��pż�[>���=I�>��>1O��T��{R��R�m>�Ń=�&>/�><�k>鹭=	B�>t���w�o�ݹ��Vz���2�btž_��>w�ʾ�Cy��
��a�#�'��w�\A��$F���x�=�4���;���>�>����hF�=\n =�J��鑽!�����ԽN<��)�0>6 �>�r��	��t��z��-IL�v�=�D>t�>�&?�m�=�~?.�ξ�[���@��־�`�Ljž��>���>������<� �F�j9�=0ӾC=�>*]=��=h�\�@5S>��g=mB>�&<a�9>4��<0�y��H�=�J$��h�>}2j>q��>W�E>2>{ ��	���5Pο�3��ξ��{�C��-=LZq�x��>�����<ѥ�>P�����%�>�:"?�C�>���=h�L�4�>�1>��f�r�����=x�s�p����G��@������=�-k�Y��X�p�0jཿ��rh�A��<�P����NOѽ4 ����> t�>�4�>�\�>~m.?Ln?�\!?�5�=�b�>]ɠ=�1�=l��=$v�>m;�>� ?��3?��H?"�N>��׾�6'�5`Q���>����W�+>�h"=MN�>X�F��j>�*�>�Zd��@ҽ���=���=47T�:'�=p�E><̑>P�Q>�7?�>_ ���N���;�֟ž�������=���������_�,=$Z�W�5��8��?��A0���<���>hܝ>X��>�7��#/=?��Z9�� ���=,"W=� )��	]>�bA=�x��c$,���A��++�)�����>�V >y�>��0?��	?]�?v�����ʾ}�#��K�bT���?�#��=�~h��@="ž����7�x�f�N������<t��=��=]x���`>�o�>6/���6�XoE>]�q�7pf���R�<�=^�>F�><�)>�d>�ϰ���ξ��ȿLۤ��������[ե>��n��D��	+x�bK��>^:���妾��=V��>!��>� �>�S�><��>Z�w>�6w���9�F=�}*=�p���0�C�Q�rC�g�c�+�^������]��2�0;e��eM��C��f��*Q����Z����>DGO>` �>��9��{�>@9/?J�S?JO??u��=�:k>*q�>�_?�h�>_�?�q ?��?�>��E��޷���<���	>R����=��<g<�>Q�,=�Sb��OE>S3=��R>%1>��Y>�>��(=i f=�X�>n$�>��?���>d�����=/�����Q��̀?�{r>� 澤��b���W���4����߾��N��� ?;�>��>a�G�N��=h�>�*��,�ѻ�,l<tڞ=�#����½���<_F$����A�\����6�=��<�p>��>?43?ͅA?.����M�K0�|7��㚾y�R^K����$���阕�n$~��a��*&���<�*���Q��;(�L<�>��E<�0*�0��=[]#�kr޽<:�{�>+o�>�q->3�>�>�B?�b>�z>���!ZI�a�ҿH5��c��"t� �j�=VC�CC�Wxý��==��>H%ƽ¹
>y��>4tn>�=�:˽���>1��;��|�Іr�f�,��� >�{���C��&붽�!3�?,};{p�Q����=`��ih�b��&8��<Z��˽ ��+>)�	�%��>!hc�>�!>���=�݇>7�J?�,J?#�0��.ڽ��>���>N>��>�?68�>��<?m: ?�>E�'�_��mC� �:�d+�0c��uE���=J�X=��>�l�=���ܚ�<>̒<_0���0��'�<!ļ��=�_'>_G�=)%�vH4�����-�5߾ dپΜ�>Q� ��_>��>G��L�����ފ���l�y��B�E>�8�>���>4��>x$������d��F;i��M�OS��U�>��H>�.����/=�jp>�_>�X�=�˶=K: >�~�N�`���=�f??��?�ݔ�4����ھe���g���ս,>��=K�ܼ=8&�iͭ�����L�Ͼoyн4H �N��=�\=�
�=��W>I�=���Ŋ�<X��>e*+������]�=��y2�=�XE��}�=u����F���ڿS���=�=_¾�>�<�l�>�X}<q���?�L8E���{�Fϒ�}�(��ko���w����=��Խ���==s9��Jڽʸ>n�׽�{����J�>\�����R�M�(��q�߽�1 ��w�{�K��h�Q���Օ���n��0��*�>�^�>�]
�n>�'�>�8�>��>�C=��>T���r/��f>�j>��>p�>|i�>�r?*F�<�T��k�P���U�W�>C(*=d�O>�Q=ْj>�t=�jr��]��,�>�0x;>���@��';�ń=0O�"�>�M�=�*L>`g�=�Ͼ��¾#�� �� 9�>�p>��B>�R��t�k=׾�\5�֭�����1˩�(i'>���;h�>��>۵�2u�`����M�=�=N�O���=��">�G�=n�ݼfu=mE]>��<lH�=��;I}=�=`Hh> K?��>�?]K>���2,�	<���н��� �G>�~>Z����'1�RV�3�)���ξ�ؾ��i>���Ü�����>[�^>��=�c����� z=�f����:��>}�!��/�=���=4`>>f�=;�>����"���l忀�ÿJKq�㮾��4�;�Q>tK�<tz侅�ӾA�P��������!S�jO��+�2�bA�=�)�>�~�>7=�^>��Y>-@�>u���y|���򂾌����9<wE��E$���Ⱦ:Fa= ］!qr�*3R��������¾z�e��K�>�v�>�e�>m�>z�>���>;�>��U����=�`>[Ǐ>`�<���>>M�>?��>�8?30�>0��Ǽ1�P��&�b������=��>�_=*�Z>��::�=���\B�<��<����������g�o<���<q(>]�>>���>��>��H�۾����޾x�/�{ȩ>㳸XS�>��e>������=�(�{�ʾ�F���B���$�>���>l6�>nޚ>�׿���K���>,E�.f�Cj=��=gx�>��[
>�.�>�ny>����*�U=�0�>9u]=��!�5XS>?�9?UB0?58<w����5��!��9=������ ��=�t>�,A��౾Z�ھ�JľX��#�q������=[�;>�$#>S>>h��=:�=J��'�=}�W���'��p[��EB<�.w�ŭ>䄻�B�<�w�lw�N$��H����ب�����.>8�0?� ��~����&��}~�����@��bݾ�_��p�>�2=m���YϽ���=�����/���@=[�:����YY�|�]�B�e#˽Lu�f�B�ˋ7�����R��MI�F!��j���s,۽�?|��>	w㼙���`��>'�>`bm>P�>�^�>$]>�펽�P�>R�>�	?�W>/��>�*?������Z����G�/U3>�Y>#71�䯤=UÙ>�	�=�[齞�����)>%**>��r�Խ���">3wI=�T�Q��=�0�>D�>�6>�W�����c���.��������>[m����<R�B�R୽*��.{��Of̾����ޯ����P�>���>N�>�q��Qľ( Ͻ�c���%�=ϊ�>r4&�d�>�>�<ټ>�Tr>},�>�'>��>���=��=�\��Z�>�1"?;�1?�5?��/���,��𽾟�`zӽ�%\���ּծ<nro>�p�"A������M�J���(��7M潗��=�0<=�..>���>�F�=�=�����z�>?c���潱�?�E�=�νIv2�c;#���>�է=gq%���Կ�ݲ�s =�xQ���뢵>E�$>���|h�=��;���=$g���"�U���?'�=I����>�>}�����˽L��=�+	��^n�o� ������2ܽO S�����6���hс��ݽ�O�6��d��K��!5����8�'��>���>��<&�Ľ.��>�c�>��>��w>�>�!>�[=}�>��>�H�>_�{>�?��>�(�=Ș"=e�.?��E�>M�~>/���a=���=N� =Zd�;|	5�,G�>Hu>�<�A"����>���=n�����<�e>�v>�<m���`3¾u�U�i�<�D���[Y�>�U���,�>�!����=T�J=�!��y���d�k�9<%M�ǳ���^�>*�>dl�����?俼A��=����j�TУ=,��=����ӝ=/��bT��P��Ļ���˽v��=;>h�>�5(?Q6?�)��և��nM���N�=:�澓#~��*��J������*���ξ>!��CV>��N�3		=װk>Y��<��>��=[�=�P >��=�b	�y>R�}2�=��V>��=�c:�\�>�w=��۽��Y����ɇ��x�<I�h��F>���=�G����/��]���rF>���>���>ap�>��>���>[�񼗙W�W�Q���Cǽ"Z������@Ɍ��x����C�-�D� �t
7=��<}߽6��� �t��I���}a��u�{�>��r>V��=z@���@�>�g?�>�>%�����>�d>ҧ�>�S�>pʸ��H�>n6�>�w�>k�=aW�,R�&��)h��8�=U1>�K�<���<�=_�:�B��<	��:.�	�vר<��= ����!L>A�>�=D�9=��=�1(?n߭<�=Ⱦa<�\
�e����=`��@�h�9G��uٜ�˾�IM��q8�iǏ��K+>��>h~�>k5k>ut�>�����<�Z|��j��<ͅ�_ܻy.=T�_���=M?�=�H�={�<��%<�@��x(�0J;�_�m����>:�r?���>�s>�LC>��2�i ��l��&�=&LK��yH>���>��>�)P��0ľ�
���GD�h`���Ӫ=k��>@��>{�n>X�B���s>����
�=���=�U��<�Zr=��i>���=��P>��nc�l�������f)q������=�>j�u��B��Ո�=U�g��t���GU=[xf��\�����=�V� s	��ϳ�����w����=��۽��4�w����n� �	���ۻ���G&�؞�
���8����2����<kP��Fk��҆�=O>>��q>�5?��>4�	?�@?��8?Z��=�<9>N1>��>�>Wr>e$0> �>si>��>��໬����sl����=�F�=Rx!��=��S>Z�T>�x<E�6=�X�<򞁽�۽�M�<0o�<������=ET�>+,>�h?���{b���ʍ>T�����O:��g}�.��Y���������������?��=o�[>���=���=���>J�>���>,/��,�%��������\L]��Ɣ=Dk�<�%R>��t<��=��e>E�K�ǻi����BX� �=��,�~��>�D2?<?O_�>S�j��R辳`H�PV��Km�=��=9r>h�>7^,>D�h��پM��������.�ν�pB>e�=�潩�J>�6>3yt�x����3<�ս�
�:��^�M{�>�ʯ>mT�>u,C>wkܼc���t̸��T{����<�GƜ>$?�>GԽ����f\	���>�>%澼q�ż~�F=��l<0��=��"�6b��D>��۾���=F�	��'�����$&ڽ�p�I����2���(��^M�n��ô�3!*�i�<��r�y�/��� ��pP>�g�>�"�>S�=F��>���>�&�>�Tz>u��>��=.�ʺIs]=Q��>��l>��=�HڼV7��%{:>\8��9��Z �gj>B�]>��>L�=)��>fO>:�w<y�����=�=3������Ҡ�=���<��=z>�ב>��?`ӯ<�ھc=�����E����`���b޷�.2׾:�N�ž�����/=�[D>��w>�8<\��=��>���>���>3����*����=�L
�Je%��=�>^.�=���=vI0=?��=�F �S��<�ゼ��������q�jtx>��5?�r�>�?f��s��1������༥��=E�)>{K{>�>5啾R����` �c��������I>�Q>+½ͼ�>��+>�E=� ��gI&9*�<#���/�$OL>��e>�->p?*>���=������
Ϳ\\��@8������'&>h�n>FK=�6�Q%�;�6�>���>�H=��˾q���s-=>�=�s^��W�Lbb�JU�gZ�V]8=#���˾�B�K~������୽ m�����R����S~���ހ��=���?��Jl=ĶR>.t�>v��>Ec�=~��>d"?ȍ�>	��>e�>�,>�� >�Hl>�
?��>��9�q4��\UZ>��>Z)����aB�˂_>��w>g~ѹ�t>�ͯ>��=`�׽�?żc�>ۓ<�����<Wr�;����M
>Y�>�g�=΁?}cB>��	�� ���6�!��f��� �&�>��Ӂ�H�b���1�������5� 6��^�U>l�=(\>���>�^|>���>��������k�<�\��"����r=�u�=��$<�a>��->AIk>f��#������q�}{h���>*��>��E?)��>��.=��<�~ɽX����g����,X>��>?b�>�?6���ھk��(��[��v׾�=�t)s��~>�9�>�}>��M<��V�#���䲦����qV��{�,b�=,�r>쨨>��/>��)>tP��˿����ѿښ���/�=�K������>B]�>w��=a�+����=��/�H�I����%���q=�9[<�5@>G�>$#=�z��1��F]>t��l�s�B�u�`�l��D�:���~5�!����1��� �E�½�&������˽ԛb�����AM�>O�\>\q�>�]�>o�?�t�>�2�>� =(>{��=���=w��<\4�>�l�>1ll>�<�=�1(>csC=Z޽r���j��
>+��=sCY<Fl�=���>>qp�</w^>W=�ýX,R�u�Y�����*н�T>��>xd�=�� ?�e=*�ˆ����/��<����ݾ�խ<�*�����>~Ͼ஺��XȾ��=i�>��>,���qoc>{�?@�\>i`�>������N���=Ф�;���E�>�>�=:�)=А�=<��=�"�=ܾB�h������G�gڡ��=``=>}SE?'��>��v>��O>z��X��b���\L��~�=Q8>���>��>U݀��� �r��N��n$'�����3�	��۲=F��>�kX>��">qڼ}m��%b�<+>�ۇ�+�<����M>�r8> 	�>d]>��g>YO��4���g:�n����f+�
�9�;V�=˷�=_����G~4��;�t<��`������=�e�=_�0=�*�=�|�s���4�G�(���1�=�uh���#08�I�T:f�9�k��伆��?50�
�����w�!��l�ƽ�?�B�b��Ͻ�I>)�?���>`E5?Q?��?��>g�j>m�>[��>W��>"�>z<t��N�=�X>E�#<'�Ͼ�ҽ
0~��?>�fe>3ܹ<��\=��a>T�[�S��+}����=�	�����"���!=`.�=�j==c�8>8�>��>����GdW�lܑ���𽝱`=.�?���G�u��־
"1������š��<��� ��
��wQ��Ճ�:�>y�>�cf��<_A'<�lj>��=/t>��H�.E��g��d��n8�}|>�?N�6��'.��;��D�=��/>�R:?1�l?��a?ˍ��"o�����e1��̾=�׾.��>��G>�����,%�4��Rc���b��o���=x9;>�^��/�ýڊ༣�uL�Ş8��j�=.�=��>��>a��>��>K�0>�$�>���=�lռ���MԿ�\���B��6��5>�½ׇ�1�p���}������U����s�*�R=�4�=��;��>�?3\?o�?�sȾ�6J�P���{���н��<��kY�괠�&�Ͻ�6н�v��FU�	R>�ջ�D�N��Ƚ�,E���ͽ����[q?�a�>�o��m��E�>'�??�^/?�#�>r	�>���>��'=?۫=�,�>Bp?[�?��?�j�>i�>��=GY�WC4���w=��>��*=YY�=V}�=�>��=Rh>�=������J���j<x>H~�=I�= K�=	�һ�v���ʺ�j���ܾ���==>��O>ާ��?�|��Ehž�X��O%�e?��νHÅ>�	�=���>��>�E�$��<m�=�w"�t���;ʙf�bo�=0��>wC�=ʁ=���� 2�3н����DO=s�E>#����`?UK%?춑>��.jX�k�t�=�-�jO� ��\�>�O�>�>V�v�p?��r1���^���X��	���=$S�>��:��(q�I�<�Y�Qq����=�dB>*��=��>5��>���>p~�>b>`>�f)���>�A뼻dA�/\ӿl���o�:�g��*��=�:$>���=�=$o4>Վ=����NǱ�1����_1P��Y�>�5>�,�=��Q=�O����ݦ���&>����>>��Ca��B�h6��Bt�A�~�8�����֤��f=P��D�#Z�uj���J���-?�>�H� �<�L?$p�>���>��t>C)�>y��>R��=P3=�R>���>�,�>�~�>8	?t�>���>Z�N���!��߾=:�=���=�e9>�]!>�=��=p���U,��;�O��z�
���I=T�=ϛ6���o�n�;��>����GdW�lܑ���𽝱`=.�?���G�u��־
"1������š��<��� ��
��wQ��Ճ�:�>y�>�cf��<_A'<�lj>��=/t>��H�.E��g��d��n8�}|>�?N�6��'.��;��D�=��/>�R:?1�l?��a?ˍ��"o�����e1��̾=�׾.��>��G>�����,%�4��Rc���b��o���=x9;>�^��/�ýڊ༣�uL�Ş8��j�=.�=��>��>a��>��>K�0>�$�>���=�lռ���MԿ�\���B��6��5>�½ׇ�1�p���}������U����s�*�R=�4�=��;��>�?3\?o�?�sȾ�6J�P���{���н��<��kY�괠�&�Ͻ�6н�v��FU�	R>�ջ�D�N��Ƚ�,E���ͽ����[q?�a�>�o��m��E�>'�??�^/?�#�>r	�>���>��'=?۫=�,�>Bp?[�?��?�j�>i�>��=GY�WC4���w=��>��*=YY�=V}�=�>��=Rh>�=������J���j<x>H~�=I�= K�=���zY���ʽ��Z���T��E ����� D>$��]L��;,A>��b�$�u%�8$�1�_�����<���>u3�>��?r2� �L�y -���KW�=.(>ꨮ�\�*=��0>��<�9=�g��?�=��:������p=�����:���<?X�>0�P>L�T�0"A�;2���B�?(����t���w>�u�>4_�= �]�cu��<��=��X�N�3���R�@=P�=| >�@a��䥻$�>��:��%7�*Ĝ>�vl>�5W�ki>���>L�><�d>-�>�rp>d-ڽ�]�Kή�6$��!C/���$���>ˆ�>;}��=��<:z���
��H���C���x�&�yՈ=`�U>s��=��=��Ҽ�|ξ&�'�FJ��I(�~���4�(�O��?:��6ݽ�h�����d�����#����3�y��r��e�{����=k�>�E>D�L>��>}��>t��>r�?�?>fB(>���>�u������5�>��?ӈ�>���>(L�>���>�3��0LT�)R�1�A>k��>�5r>�>Ƨ=s� �U��=����=r�=�r.�	� �j�Q�^3��"Q��>%����<X��=V/��W�޾��޾5#F�Y�@���ـ��?kЍ>�hݾL�/>G�R>gn��0'�� �����}rʾ0�S�B��>���=�W>�m���)7����<�yQ����6&>
+�<���LK=�P}=}ϯ=^<��=!�l{�=�*<�������ō�O�/?_��>��>�=�*��1�U��\�qq%�=�KM>�}>V��ɩ��mҾ�� �(hM��	�>�=B�G>KD�=ڡ��am�=7z�>�EG<�@��	=�%�=˛��b@�=zrD>�>���>�T>l�>L�>�%���塨��N��@i��㬾 D��ܪ;��D=�Iս�D��Ľ��A"
����=�'�=@�y=`K�;~��=��=f3�v�ھ�ɶ�,�=�Ǿ����Ծqr��G�r��}k���:�(�����!���ʴ����Z���H^o�[Θ��j?Ŏi>��}>fݵ=�1�>1t%?��?-���Y�<E �>|�	��)b�{/>�O?��?(��>���>Kh�>SPe�s��=��c9>e��=΀=,�=��>���;�-=�=�A.=H	5���������L�� 3�O<��>�(>Ձ�>Q��>��6��D���X-���k��N(�p+�>��=��y�O^+�pR�=K)A�0�Ǿ���|��^e���y�?j$�9W�>�g��ɾ2X`�0c=M7�<ى��V>��z�I�/>�'�;���>�<>����Tځ="���X��0v�*�{�k>6�?��??S0?3Ä>a{$��r0��F<�@�׾`	_����%�l��Ӿ�������2)��� ��N>{껞닽þ>�1>������ٽ���=����Wj�p�>D:�<a�>��#�
�,>
�>){����>��>nn\=��=;�Կ������о�;�A^���=�m��̊��vt�	T�I��蕇�V�=���>4�4��>:f�>M�*��h+= � ��z���mҽI�a=ȼ��f⧾z>Ͻ9K��o:;�O�C�N�������ίǾӥR��������nd���I��^�<N�?�k:��^��|�=���>�O.?Q�??�S�>}k�>d�>G�?���>��>�)?��>�i?(?���<��:g�m�����>?{]=�=���=:m�=2�G�<�J=�)C���%�X�8���;,����>��$>�U�=���<�1�=*=C��=9����]�����˾﷾��YL�N�M����K����ȾX���h��ki��(i>xҭ>��>U��<�,�>��>S5Q���1��P>?�4=h%�<��=��6�����,߽�K5�՗�<�eȽ�����b=��>�T>�J[�8Q=s
?()?qa�>�Y����J<��!s��q@�l�t2>��x=N$t=�
��%��=9^��(���&�	�� [=ŧ	>q������ז����W�;�K�<���>6k{=b�B>��>]��>(�i>��&>D� FC��:ξ
!'�_#ʿ���C���:�EG� V�=�>�=$ɦ�Z��=�ƃ<ˌ�!X�%�m���"=E5�>��'>X�ǽ�^����9J��������F�=�p���[�6虾Djy�.���Q�J�Ɋv��������	��?�W��׽��r�)���4ݼ8#?�Y�9D�����5�/?�m?�?�Ԑ>O@�=�d�>��?�,�>��?�%?3<�>k>A_�=�]�<�q=�R����ͽ{�_>�%>�w)>^�=��=��<I��Gx}=}�=2��<�
�A��=;h�<[�=̃=G��>��C>D�@������-`��p⊾�뜾��>�푾�=�����W�Q�L��߾�� ��C����ǽ�0>9�g>���>Æ�>T�:��G�]��=OU�<-,�;yiB>]�_��5���/<O�����=�Z�����<�ؘ=��=.�z�^C@����A��> &?�?#?w{�j�̾Ͱ*��x�^"��
��=w���p���?B�������Ҿ�0�V����x���>�@�<��>���=�鯽�䚽)�=�c����=D�>B>�_4>�o >���>cb�>h=�>��,>`�>�����D���Ͽ<Z������Ӥ��f=��=%�*>�Y>�UU>-���w��{=��D��>���<�D�=��(>3ka>��=�˾�3���q
�Ċ��X7o�Qm�jJ����Ծ�;�m׾����:��R���ld�P�H�Ⱦ<��=��E#?9.�>�߲=�[�Hb�>��>�)?��{>��>B0>PZ�>Q��>��?��?#��>�?���>B��������Ӽ�k�R��,0>�ܝ>j�/>'�K=��>�'��:�=߹>��=mm��<��!�0���c�� =���*=ϫ>�B>>��C>D�@������-`��p⊾�뜾��>�푾�=�����W�Q�L��߾�� ��C����ǽ�0>9�g>���>Æ�>T�:��G�]��=OU�<-,�;yiB>]�_��5���/<O�����=�Z�����<�ؘ=��=.�z�^C@����A��> &?�?#?w{�j�̾Ͱ*��x�^"��
��=w���p���?B�������Ҿ�0�V����x���>�@�<��>���=�鯽�䚽)�=�c����=D�>B>�_4>�o >���>cb�>h=�>��,>`�>�����D���Ͽ<Z������Ӥ��f=��=%�*>�Y>�UU>-���w��{=��D��>���<�D�=��(>3ka>��=�˾�3���q
�Ċ��X7o�Qm�jJ����Ծ�;�m׾����:��R���ld�P�H�Ⱦ<��=��E#?9.�>�߲=�[�Hb�>��>�)?��{>��>B0>PZ�>Q��>��?��?#��>�?���>B��������Ӽ�k�R��,0>�ܝ>j�/>'�K=��>�'��:�=߹>��=mm��<��!�0���c�� =���*=ϫ>�B>>(X�>���:~�Z��k꯾E�������U�=�J@>^þ*�a�z�=M�޾HA�s�E���z�Wܪ�M�/=��Z�?��>���>t>�=R�=~&=���A������
�q�b���i���H**�i�p�2��Bİ��I�>eg>cK�>��7?�.W?�D??�>���)]�V����;;q��꽾K����<������@��YX�6�!�Q�����=�+ǼS�0>(�W5����<O
�Q
^�"�>�:�=��=]�>2P}>�>~9[>Sk�>�eh>3^ؽB�׾�������꺛��xH�U"����jH�I�3>�u�=y�
�!�=���ˤ�V�>�>��>+�>��>��a=��=�����Ҍ��������|���3㍾���k�f��݂�Tjg��j�G-�#�=�*�1�8>V��k���rѽ��ѻz��(?ew�>��;a�W��3}>D�^?9�-?�\�>�Ѡ>!�?. -?�+�>�(?Iy?4?�n7?;�?�ݓ�­����}e���=f+V>�Wt>��>��O>&�y<��>��*<�x��k?�K�<��=J��0>�=9�>#*>�s=>�?�AI>q�N���N���ތ�34'�����pO�ɫ˾���b(��+���S0����2�;�{#>&R	>�a��ǖ>X�>ϳn����u9��� =$5=�����n�|h>2wu=�z�>�W>����C�.=�0>r�<�e�=~�U:0��>�P!?�!?��1?�����{¾�Y��迾�.�=�5:ڮ�=/K>x�E��b߾S	��vҾ��m�%n��xF�HE(>��>�1>�@g>�磽��½Q�ɼ4\>�B>�kѣ>V�k�۰�����>ČM<$泽̦E��,6��A��ۿ����1s�	c��F��V�=�%�= ��D���xL;��������I�e>8��>�5>�#�=|�L<�W�>V�����{�*�����pC�Z�������Ž
�9�`p��(w�;�R�,|���f_���)�mG��uE�3�l��K�A>v>z��>A��>�sR>1��>g�$?��>�E#?�3�>�??���>q�?���>�q�=���o"w�~/�<lQ���`��w�=��5=y=t�<Ƣ">B>�=|�6;D��[�eՐ<qv��>`A=���<���=��=��=�wk>�<d>K6�� ��G�n/��L̖�7�������7�㾭����������Jz��;#��a>�M�>�>�>���>o2�>�?��.�1��=:b>��Ţ>�3>�0�ݫ8��>�;T���=�� >�'�=�l�=.T=�Jս�RS>"�?�n�>7/6?�ؽ�n;��R��)����T��=޾O�DA-�a�A>�����a������r�ؾ�������CJF�0��=�n>�J9=�	�yz�-�
>�~�=)��=��>�V�=_
�=u��>{t�>/����٢=�G�n��� �L�޿����x����e�8ҍ�.�<?�}>·k= �|�԰2��4}�����L	����=��3>%{����~?�����¾����/�<�����¾1�о3���c����:��Ȧ��������"���ܖ�5|��HWu��x��/����K�>�]�=�m>7j>H��=B?
�=>�T�>kh$?���>̔ ?�,?�!�>�&?�(?[��>'��4��Zm��ʜF�\uG�`I�>��>{�>��
=6	>��Ҽ���;�����*>c�}�ss���[���=ąC;4O>>U6>��>�wk>�<d>K6�� ��G�n/��L̖�7�������7�㾭����������Jz��;#��a>�M�>�>�>���>o2�>�?��.�1��=:b>��Ţ>�3>�0�ݫ8��>�;T���=�� >�'�=�l�=.T=�Jս�RS>"�?�n�>7/6?�ؽ�n;��R��)����T��=޾O�DA-�a�A>�����a������r�ؾ�������CJF�0��=�n>�J9=�	�yz�-�
>�~�=)��=��>�V�=_
�=u��>{t�>/����٢=�G�n��� �L�޿����x����e�8ҍ�.�<?�}>·k= �|�԰2��4}�����L	����=��3>%{����~?�����¾����/�<�����¾1�о3���c����:��Ȧ��������"���ܖ�5|��HWu��x��/����K�>�]�=�m>7j>H��=B?
�=>�T�>kh$?���>̔ ?�,?�!�>�&?�(?[��>'��4��Zm��ʜF�\uG�`I�>��>{�>��
=6	>��Ҽ���;�����*>c�}�ss���[���=ąC;4O>>U6>��>�wk>�<d>K6�� ��G�n/��L̖�7�������7�㾭����������Jz��;#��a>�M�>�>�>���>o2�>�?��.�1��=:b>��Ţ>�3>�0�ݫ8��>�;T���=�� >�'�=�l�=.T=�Jս�RS>"�?�n�>7/6?�ؽ�n;��R��)����T��=޾O�DA-�a�A>�����a������r�ؾ�������CJF�0��=�n>�J9=�	�yz�-�
>�~�=)��=��>�V�=_
�=u��>{t�>/����٢=�G�n��� �L�޿����x����e�8ҍ�.�<?�}>·k= �|�԰2��4}�����L	����=��3>%{����~?�����¾����/�<�����¾1�о3���c����:��Ȧ��������"���ܖ�5|��HWu��x��/����K�>�]�=�m>7j>H��=B?
�=>�T�>kh$?���>̔ ?�,?�!�>�&?�(?[��>'��4��Zm��ʜF�\uG�`I�>��>{�>��
=6	>��Ҽ���;�����*>c�}�ss���[���=ąC;4O>>U6>��>�&�;9=.�E���P;�Qܫ�r�mH�;H��_���g��O��?��k��]��B	����þ��T��>��>� I>I�/> >���d���3�0� <�ӽr�4=�ϣ=Z�T>�
>�c�=��=��B<�"7#�:������<S0�Ӗ#>��?�?V�(?4�M��`��U��$���v���U�=]:�=B��=�A/>b/{�(�ƾ@��t�����;&W��v�>H=V6�<��>ܩe=$"�<RY���
>��<�ȇ=���=5'�>��>��{>AH�=�=�+A�3BX��P��h��z���/�׾b����u<��V=D���Ѿ���.�v�B��VȽ�9��>�O>9�>YNI=5��<���=[>��L�=��������r�����T6���P�ھ彪�������wT�l�<��H�`�?��#}��I�ǔ�h'�>�`Q>�Pk�8����>',?ࠤ>��o>���>��=>++�>~��>���>YT?�?��
?.G>c󽷝뾄>��Ӳz��ߵ>)�=�&>�l)=c�%>������C�ca��A��Z'Žot���*�n�<�T�=�<�=��>�L�>�,�=1.:���_��vS��e�����'��P��H/�>�w>ek�<�6�bl+��\ �,��D���X��$�>9�>�c�>�z����ۻ_Ċ�YɅ�Y޽j�ڽ+�x>�->�9@>�� >'����<N�}]Ľ��ٽϸ����Q�}>�*�>0�?��s>�?ź����1���2��XھA㔾�`�=Cy����>��K�����S����}K$�t�L�+ڔ�m�C=2�0>#T>^����]I>��=�>*��l`>����3���=�c>�W�>�$�>P��>"��>��=�D,���Ӿrۿ���������;��7�ً&=�w>�).><���̾�]ξ�m���=��S>m�'=u�R>+y�>mWQ>/g�=�.˾
��x�˔C�ч�Kjt�窶���齇�:���C����Ӏ�O�4���O��R)�b�z��?�t����^�¨�>�Y>Q�>7H>7~7?��?�>!?�/a>2 �>�c�3��=��f�Y��>c?��?xR?��?��>�#�Ч˽��T��c	>9�=xt6>�g>�j�>e�ĺ�d���+O<I,���ֵ���qN����p�瓎��ڎ=|�w>�=D>�{?��q=�����ľ(O�8Ty�~���k]�>�t9�Y�ҽ��ͺH�d<`�$��Ⱦ��aX��偎��P>�,|>h۸>ժ�>������`�@Jw�R���@��g.���M�=8ѽ<�ļ=Y >i�}�j$1>��H>�W>��G��!�TW��JF>�s)?/�?� ?�e�;��羺��1�����oؽ�_�=5�=cb�=���>䙾t�>�c��x�}�#��W�/>agq>�� >�>B۾=q%��m�=���=��B��dZ=��1�A�R>��->(�c>�,,=y�P<u���*��ӿ�i�����i��6_<a&>� 6>6EE��<۾Q�=䏻��O=f">���=L*�=��Z>�=$/�LTa=�̚�)�I�1�(>�`=.��ZGk������w�2���inO�`. ��C�/Y��T[�T�о\�4�4�,���B��8E���=[�>Ӗ>a�u>|r6?�Z�>g�?5Q���|�>�=OZ>�ֽF"�>(��>�?���>'^�>��ʼ��-� ���<]�Nb!>�"�=|��=R��={^4>F��=̫�<��=B�>X�D�\fP�/���e�R��t�=tA�=br\>�$?cgq�Y�ܑ޾\�6��ξ��ھ��?�����>yr�>��*�a;�?��g#��}��<�E�d\�>c�>劓>��>[������G�>o�2���������>$�2�xP�g�>����"�==F=(�>��%=�Nϼ>,����O>ǲ?�>s[?����P@�~��v��M*�\n�<�AE>
��=�ؼ�R����+��V����������J�!>?��=皖=p�>	��=gjҽ*ɸ��o>w�E���k=܌�=�>���>AkI>X�9>n���&I�����%������R��ؾy��-?�>�U>�;���þ[_)��%����c���=�)�=��H>�r��^=����эu;M�n)}�S��#�{������xվiED>u�Ⱦm��='�;<G8=���ڀj�Eƚ��x4���w��Ux���C=��>1�w>���>�M?q��>��>mM����+?U�5�(󍾲�>ۻ?p�?��"?~?���>��l������tL��	I���>i]S>��>�<�=(}�>��޼���q�=kR=L����v=�Ͻ�0�=�潯��=��>�xm>�#=?*��>��-�S7����<���2���:�%"<򯏽&�>I���8�>j�G��D�,=o���Ѿ>����0>��>`�R� ��=��>6]U��Xƽ��׽���=�0�=S��=�P�;�x%���꼬�x>�̆>I�1>��=ݯ_�lp�=��3?�<?�&?�����MϾ7�߾�[��T�9Е�������=�#=E@�����z'�����s�پ�XP���%=�G><:j>���=�=9<-D>�ln=S�2>F�>�Qս��5>�E>�"'>i�>A�1>4J=�=���X����ֿ������DoѾ3r��=j��=�o4�;���\����o������Mc��f>j<�=V�I>��>�\>�WF��{>9��=�=����(|���n��q�: ��(V�2җ�z���>���d�Q!��8�2���s�Ɔ<�fj���=��P�2��>��A�O/,?�%?�+?.>��a>�-#�~M�>q��??Sû>.�=���>���>�,>�
%��6���-;��C��<rs^>m=>�<<�윽��<N垼oȼ<	�z�D=����a���?��==��=�U?᭱=vZ�$W�)�9���о҄��?�F<����H�<֩E>/��k�Nb �k������kg>�e>��>�H!=�̼�����D�ż�l���jӕ�_�z=�Vc=��=�Nѽ���ۨ�<�=s�>s�7>�c5<y%��M�=*�#?�'?46?ՆY=+վ[*��_���������a@=S��=;�>�t0��뚾|���:X	�cq�H�N��{��U�>���>l���aZ����=]>�~�<� >����:�UH
>q^>�>0��=Z��*ǽQ���<�z������}=�}n��b>5g�>p�>*W���F� �o=rUW������Z`>c�=>ix>�h>���=X�]���I==��W�4=�yf=.�=��N��*K�IL������Ao�������V�W�=Y5���q�^Qͽ��:�z�$��iý�Br��SY>ê�>��k>��>�v+?~��>�>~3'��R�>Ɯ�<���=7a���j�>���>%z-?�d	?ɭ?�`�=�eT��*��䈌�rMb>�-�=(�M>5�d>]J�>pz�=|R*�����l�=٪��a��=� �v����E�tZ�G݂=V�,>�^(?l��>')��	v������1��>���>,$�������%���6��4�����ļȩ�<���>yb?q	�>8�>{m7��pm��齼�Ƚ���=cp>X@�=Ɠ�=.��=>�r=]�e=N�Ҽ���x<0��;e�p>��.>dl�>��>0/B?��"?�d�>������M����m���;>]*���y>M>`��H>��r���)�+Ѿ{�D=m�$>Z�h>f>0	 >�|�=�;p���=x';2󍽦�>���<);3�>��>�ҫ=�.�=t�:���v�{BͿ״���we�`Y��o��=
��>sN�>�<���e��ť��V�����>�>� �=��c��=�u��jP�a������r]�=B�;�w�t�)#��b��q_־�k �A�����4|�X,��U�D-���^��� ��|���S�<���=#�>�	W�e� ?�K�><W?"��=!#Q>�e>���>�>�E�>�i�>8 ?UG�>-�`>�; =[�O��&�]�����oq>��l>�>˒�>[ڽ�B�=�"x;���)�:���=�1���O=�� >��=ʀ<�S�=��?��=����\M�����v��Û^�/>�>��>�u�Vǡ��?���?��^��2���џ�=�`s>L��> �>@��>��þR���jq�=���������>��4=q�>�]�=΃=[x�:�$=���<Cf�=ʦ�<�F>���=8��=r� ?�J�>���>@]S��}վ0��۞Ǿ٦վW�?�@�=A#�>���>c��=y=��	�ɾZ�3���PB���;��9=�w>app>A�>(�&>�u�=��=n�>iK�����э=έ�]v�>9̲>�K>T�m|_��gT�\Fɿck��pr����|��J�,��>�M>`;�B��4uͽ�s��g��R�>Q��>/�j>4�>Ŀ#>����������8��I�h=Xdx��'���޾���ȓ��-�Ծo����d����=�V����s�;c���!��o��{����*>k<>��>�0�<f�??��>)d�>Ly\>��>_�L>;E�>ŸX=m�=�>{�>j�>�Zk>3\z>r���f׽A����g>�X�==>!q|>L)�>�ܽ��=(�ＭE�<
�;�=�"�
�$�&��3��MX>�,=�2T>�3?�ZH�b��z�����'�+죾g���6�>n��>4�>;�g�-Z��k��
��Y ���=|��>0|�>O�>�Oh>aϽ>�����҇�����'���=m�A>񪵽�4h��M<=�V=D3�<��^=�C�6�n=�l��Du�=�~\=�>0?��?e�>�#e=�ľ�q������"޾Pq<�Ⱥ>�7�>�>P��>^|�: ��� ;��� ���߾������=�dk>;�>(^�>�R��i�>�)�@�O=����ZK^=��l=z<Q��=1�">9��>�*>�$v=7p���yٿ���\�s�8Y��>)�ts�>q">>�:	�![¾��B���g�>K�>t��>`�>Ҡ�<�ʂ���+�V3�>��1�>�u>�Ԟ��/���
���@<s�4�i����3�'��Н0��P;�O����l�Q@������F6�r% �O\�>Wc>5	"="�`?5�>b!?��H>��>�'=�c�>_h>9�7>״�>�E?R��=y�&=c�@>��-��þU���;��=�����޽Ǎ�>��= �p��/>�!�=�p��mP��q�=��;���:�l:�d�y=��5=��n>�$
?���> �[���0ݾeN׾�+����?u��>����,���%�k����������ۥ���e>�L�>�	?Ֆ>#�>�ƻ��Ӕ�m��<Obf=�+>���=bJ:;��9p� >?�=�*�=���_.F�(��G�><̉B>��>���=���>(�?L
�>$j���j�������L�=�ƾ�">�u�>q1>�m�>�[)>u�˽]b��,����1�ྒ�R�g->T=�>z$g>ѵ;�7�\�|<��r����]��<��>��=o�F>�9z>٬�>�۩>�?>�;��An��~]ѿq���9!��?���� >{`�>�@<��T���D@>���׳پo�G=8��>u��>�Sk��y�����7��Ͼ�1ݽq��=�s'<�S ��ɾJ�$�7��/��2��=�����s�u�{�?��g��������U���s��o=���=��>�b}>�r?eE�>1??��z�'	��B��=��@>j�[>���>��}>��>t��>�E>��Ž'�\�r]���}��O�>�>�Lr>>b#>�C>	�<�)_>�U��S�S�]�мI��'�7���=�
�=>�P=@e=|�$>�^(?l��>')��	v������1��>���>,$�������%���6��4�����ļȩ�<���>yb?q	�>8�>{m7��pm��齼�Ƚ���=cp>X@�=Ɠ�=.��=>�r=]�e=N�Ҽ���x<0��;e�p>��.>dl�>��>0/B?��"?�d�>������M����m���;>]*���y>M>`��H>��r���)�+Ѿ{�D=m�$>Z�h>f>0	 >�|�=�;p���=x';2󍽦�>���<);3�>��>�ҫ=�.�=t�:���v�{BͿ״���we�`Y��o��=
��>sN�>�<���e��ť��V�����>�>� �=��c��=�u��jP�a������r]�=B�;�w�t�)#��b��q_־�k �A�����4|�X,��U�D-���^��� ��|���S�<���=#�>�	W�e� ?�K�><W?"��=!#Q>�e>���>�>�E�>�i�>8 ?UG�>-�`>�; =[�O��&�]�����oq>��l>�>˒�>[ڽ�B�=�"x;���)�:���=�1���O=�� >��=ʀ<�S�=
�	  �   �Π�[mb>�Z�{޾�qn�~�I�t��{J=E�K�Q=����Y־G~���=�	>���6!!�y
��U����J?Fl=�N���V�es����>�ޘ>�Ϯ>�^9�[|�ND@�>����=P��>Ū;>����/�qG�av��,s>B?H�h?��r?$��a�Q���[��}�~���z6?v�@>�?�/6>ܠB=r�˾"�V�i��	]�M��>���>�\��مV��1}�ިþ[����>�l?A-�=�8�>	qI?��
?�l?�"<?�*?&�>'� �a��A&?���?�=��Խ[�T�99� F�<�>
�)?�B�.��>��?��?��&?�~Q?�?��>� ��<@����>�a�>�W�Yb��3`>O�J?%��>?;Y?�Ճ?y�=>�}5��ࢾ�ҩ�@t�=�
>��2?�2#?M�?b��>��?��]�R���>�]?L2�?��o?���=V�>���=�G�>�ic>Z�>���>L�?G7,? �w?�S?sy�>f$<)�Ž�~��$.�C��<4����5=�'�<NZL�Dh�]s����=^&,=K@��=����/��ק�O� ��ɧ<�W�>�w>�2��\�8>"��J�����>>�,
�"z��-f��$#9�Nt�=�g�>�< ?6�>5)��e�=�<�>D�>Z��#�&?n$?^F?з+���`���۾N[��{�>�;C?�G�=@xp�����:�r��9=!j?�9[?B8X�������b?��]?+�P=���þr�b�]S�~�O?�
?]	H���>��~?��q?M��>��e��6n�/��:Gb�>Jk����=u�>�E���d��@�>ɘ7?�;�>��b>!l�=P{۾״w��Q���?0��?��?k��?�)*>��n��4�����ao��]?M��>95��T�%?���J���w��
s���ž���D)���d�������b(��!����G�y=�?T�f?T�k?��I?�<���g��F_�� m�X�L�f�̾=�1�*-:�L�Y�YT��s������{�K~x�w
>q�����=��в?ϋ:?��c��>}叾��	���־�!|>�uɾ�J�*��=������<ga;=�g]�A�����d�?���>U׽>S�8?�<X��8��N&���7��8�d�d>p4}>3h>\x�>�<h�3�=�Ö���H��+o���e.�k�c>�nY?8�R?��{?��O�$��CV��3�ެ���ym)>���<�>�\D���P�A7�VA���k��S
�ڞ���H����=�z?h{9>q�E>>��?��?qm�14���wh��a ���<�[�>��V?���>�&>�YH� 6����>�h?��>�>�ܽ�q,�>��ȱc�G�?�e{>���=�|>.hM���A����NS��}jL�=�">� k?��v�~|�)p�>��h?�B*������>q�<yFE�\sھA!Q�Y�>��>��f�-\�>�΋��@��X���\v~��-?�x?�k����*���>�~%?��>�2�>8�?�c�>G���,�=:f?�W?��I?@�9?���>p�=�_��E�ǽH�%��Y'=U��>-�d>���=���=G�)�"�a��.��=�=>�s����)UP<d	�B�;Ϛ�<�$/>����k��v��u='���۾B�ξ�Mӽ5���ǘ����n�|յ�����]#=�Q&=RX����M牾=�L�1��?���?=���;ݾ�p��gD�� �Z��>m +�[�G���������?���Z���'��n3��O}��X\���E�F��>�m��˿	����m6���7?��[?��b?{}ؾ�yL��i�>yk<�=�Ex>�ʾ)�����Ͽ�.���3l?R��>e�˾l�)�vI?1?'�ۢ�>�"�<3��d�o�v���I��>� ??,M��G�ֿ����5U>Bz�?
�@u}A?��(�'���U=�p�>V�	?�?>1�0�r��찾da�>�>�?��?�N=�W�z��S�e?'5<Q�F���ڻ��=k�=*�={u�n�I>SZ�>����A��&ڽ4�4>��>��#� ���2^����<�]>��Խ���5Մ?,{\��f���/��T��U>��T?�*�>O:�=��,?X7H�a}Ͽ�\��*a?�0�?���?%�(?8ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�߅�=h6�ˉ��z���&V�z��=Z��>c�>��,������O��I��W��= ��7ȿbE$��4��C=9*����X�v���|���cH��
��(u��,��T�=�a�=3X>B!�>� R>��X>[R\?��l?���>���=9������L��)�;�����0!��̋��o����ut达i⾍�
��k�>�,Ǿ�]=�!�=2^R�Đ�� ��a��DE�[�.?�p#>
.˾�(M��/<!�ʾ������t��¥�.;d�1�1�m���?�cB?���{W�"�����o����W?�����a���L��=�̴���=��>�9�=���P@3�R�R���G?��?h_Ҿqjl���>v)�=�w >�?��>��l�$��>��T?]Q���~��>�~`=<��>�_�>-/U>8t̾"�Խw	8?��O?�$	�eS~�y��=����o�&�j���W�=c���к9|j>���3`������X��;{Bd?���>!�1���IPz���=v�'=4�?�I?��>��^?j9[?��H�������,����m�T>C�_?n�\??��= q�R`�A���nA?(z?���>p�ǾLr��;��5쾾h?Dys?�M?���<�W������ƾޤ?��k?c\���ם��$��Ӿ��>�(�>�j�>3����b?�U?�Qv�"����g���C;���?�P�?b�?�!�H�̽ڄi>�-?͍>�����;���r=}$��� N>��?�܁�d닿apI�wӾ�VG?���?d�>��A���뾃��=:ؕ��R�?W�?	;���
j<���Ll�Ρ���-�<jl�=@��R�"�x���7��ƾ�
�⮜����q׆>�N@>�T��>2�7�c8��VϿ�慿о��p��Q?�H�>%�˽��x�j��u�e�G�4�H����z��>��>Tm���s��L�z���;� 0ؼ�1�>��Լ�>-%X�e.��%-��U�';?��>6�>�@�>n*��z~����?F����ο�,��e�� Y?�&�?A�?^� ?7_<j�^�S�l��{��l�G?,�r?�Y?;��vG��7K�ݾj?Jc��ZV`�Ӎ4�IE�U>!3?�C�>�-�K�|=�>���>e>6"/�O�ĿIض�o���U��?���? n�l��>[��?^r+?�g��8��Z����*��0�?A?/2>,���n�!��/=��В�.�
?�~0?&u�0�]�_?+�a�N�p���-���ƽ�ۡ>��0��e\�N�����Xe����@y����?N^�?i�?׵�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�j�>K�?���=�� ?]�>� �������=�->�/���>��F?Z��>�b�=�>=��v0��y:�]�C��1���	G��~�>/o?��N?��
>��ʽ����.�]����KǽS%μ����y���ɧ�m~�=o(>˵�=�E���ܾ��?�F� sܿhq����V�u?�>�r?� �i?��IB�=�w[?i�e>�HӾ����1!���D�S�?��?_
?M��D��M�=*�?�o|=�گ���I��l$�K{�>�8?�>������d��
>���?��@$��?}��O%?'��ދ�Z(u�E ��U	��S�=�;?Ȱ��yq>E��>Ef>��p��֡�͓y��> V�?:;�?���>�+g?�k�v�1���<Zӱ>ɅJ?!+
?TѮ��l�����>
n
? �	��׍�u7��bc?�v@c	@��`? ~��zRҿ:���w��������=�=1�#>�̽��=d�Q=��4;�@ü�->��>�w>�̃>��8>u#(>�>�I����#�{��������[8�g���<�N;����Q��=��m��,�Ѿw���PԳ���O��&I�}+�C5���=�k??��{?��g?��?-3�iHC>F}�zt�>c�E�R��>�����t?ƃ? �|?��{>������s�ĵ��hkc���Ⱦ�BY>x�>=�?w��>��'>rY�=�qN>Q�>U�>��=�/�=Τ>���>=��>6��>�ѳ> ��>�@ >���=@o��Τ���k�Y :�`H`=��?���MsN�ͦ��!�������,>�0?���=�[����ʿHq����Y?�TY���#�#��e�;�,?�[?��%>Њ�������u>�����^G�{�>X�l��(�8���>�T!?�f>�$u>{�3��c8���P����Dj|>^36?�趾�K9���u�B�H�Zݾ�<M>ľ>�HC�)h��������zi��k{='v:?΄?0���Ѱ���u�4A��cPR>&\>�=/��=�M>=�b�f�ƽ�H�8%.=���=��^>��?��2>�E�=�
�>���m�C�,R�>��>H#3>�/<?O�"?i�=��%���\����3�ٓc>Ғ�>��>˔>�'R���=�T�>n�h>�K?�9t���*yA�R O>[;��I^�Y)��*��=f������=���=�b
� !B��6=�~?���(䈿��#e���lD?S+?_ �=�F<��"�D ���H��G�?r�@m�?��	��V�?�?�@�?��H��=}�>
׫>�ξ�L��?��Ž6Ǣ�ɔ	�/)#�jS�?��?��/�Zʋ�<l��6>�^%?��Ӿ���>/`��������}�z��k=���>D�F?���G����;�0�?�9?�龓t���ɿ��v�(�>�@�?+��?Q�l��ę��9;����>,�?�Q? g>zܾ;�Z��,�>B?�P?�>�>C\���&�͘?�?�?�?'�9>��?�uW?�=(G>�}5�껾��Fc����>��'>������<�{��<�"�Z?����{�i�d����?*�>5W=�o�>��H�eh۾��W�}Y�����/I�Û?-�C>��4>��(>=5�>�|�>�>+��h�������	�^�K?=��?���3.n�7A�<Q��=/�^�k ?uJ4?�c\�O�ϾϨ>U�\?�?x[?b�>���>���鿿�|���ʖ<��K>y7�>qK�>����0K>>�Ծ:$D�Ws�>�֗>涣�:ھo��Q��$K�>�d!?2��>�֮=� ?��#?|�j>���>�=E�c6���F����>���>~T?ۍ~?��?)��M]3������͡�Wb[��1N>��x?2[?���>����:���x�C�t&H��?��ू?�g?��彂#?w.�?�X??աA?,f>z}�n�׾+����ڀ>��!?����A��M&����~?Q?R��>{4��H�սDּ-���}����?�(\?�@&?v��b+a��¾$6�<�"���U����;�iD���>@�>Ԍ����=>�հ=GNm��D6���f<Im�=��>'�=B.7��v��q?���f҃������i���x�0g>@֢>�	�j��?���Cۀ���ÿPz��,_�C#�?�R�?��?��zw���V?K�?�X�>�?\���n�ھi���y�N�۱��)�y�9K�>D�D���ƾo���mm��y[��+�S�N�|�͝�>�s�>��?L�>�w=K�>�@��Ѱ�?wξk�۾�=p���澺+2��f�^����L���S�;�r˾�N~�
> ڄ����>x|?Q�i>+�V>f�>������>��y>A��>��>n]�>`��=ٜ���iý�	�LR?������'�;�辠����4B?Lmd?D�>
�h����������?Ԅ�?Pn�?u5v>8}h��&+��l?>�>{#���m
?�;=�q��B�<fR����������\��>}9׽�):��M�8_f�#^
?�'?�{��+�̾V׽������+=N�?�"?����E��k���C��J����=7]Ծ�cH�F�!���p�s�� QN�\�q�,���>��'?;�?�	� �5QH�����d�S)�>�?j�>�Ҽ<v�:=��0��}5���h��u��G@S��|?�Wu?�l�>��G?�Z8?�mU?��D?v�>Ա�>q��^��>G�� ��>�g�>(9?�##?u"?Ic�>}� ?�"b>0��5��ֱ;��#?�?�\�>3#�>��>���"Ľ@_~=f���d���^�S�w��=�AԼ�	��%ƽ]�=_�'>�Q:?�ĺ+A�oK �fP�>�L?S1	?�>��9�$7��ɼ�<nA$?��?$>�`���Rc�CǑ��
?IXi?ش;�~����&>�>ta=���3�=��`��^�<�B�����c�p=`>9�o=�p���?<�Ͳ���\��C=���>X�? j�>j}�>��~�������lB�=�|[>�U>w�>�M׾󫊿�^���Th�|dw>���?>��?�U|=�R�=���=-Т��/¾���0������<��?3�%?�]S?�ݐ?Z�:?�"?3�	>��S���2��������?�,?I}�>�����ʾ��Fy3�X�?:T?3a�����9)���¾��Խ��>|]/��4~�	���D�(}�\��<������?���?��A���6�͇�!���`��K�C?��>�X�>��>��)���g���ik;>̇�>IR?�o�>^�M?�%|?��\?g�^>��6�{1��Lᘿ^&�9I3$>��@?��~?��?u�{?f��>�!>��1���p����(��b�k��0�E=)�]>#/�>��> �>��=���諬���>�|��=��l>�s�>�C�>�c�>ɭw>R�<@T?{��>0/���'�������/� �A�?_��?��4?��5=���K�N��u	��S�>6R�?W@�?a�'?M&�d(>��<X������r��>�F�>�ޯ>��#>P�=�R�=?�?b�Ž�
ᾙn��W�~�?�b?<1�=J�ſ�%q��m�����5|<�{��Fld�����sK\�u��=T���c������*\�MN���ْ��o��H���.�z�l��>ϭ�=���=<^�=
��<2�¼r]�<��C=xɋ<�=�;y�-�<��A�����̊�)!��L`<�H=����4Ǿ��{?�SJ?�Q0?9�??�5x>�n>%����>/6}���?�B>ߎ�l����kB��
��<闾�C׾�@Ծ��g��\>7�T�Ň>B�>k��=�g�<��=#Ol=�[�=��� � =#B�=�A�=�Z�=���=�P�=��>j6w?\���߲���4Q��_��:?�8�>E|�=тƾ@?��>>�2��旹��b�-?���?�T�?��?qui�Fc�>_���ێ�Vr�=�����92>���=��2�'��>�J>8���J������4�?^�@E�??�ዿW�Ͽ�b/>w3>�V>��Q��31��RZ�c���X��!?��:�ޘ̾�8�>��=�OݾvlƾȞ4=��7><�e=L���x\�m��=����+G?=�r=`ĉ>�H>Y�=6��a
�=�O>=�_�=�1T>�";����>�)=�B�=~�_>"}$>�`�>w�?q0?�gc?U��>�p��Ѿ���j��>~X�=?\�>6��=W<=>�r�>�K6?aD?��J?���>ڥ�=�>�ө>	-��Sn�R�⾏����e_<@��?�#�?�>���;��B����U�=���̽��?��0?H	?AΟ>Q��4d��v�"��~�;5{�1_K�=��DV���T� ^��q��̨=6��> ��>���>8o>!��=/�9>���>�)�=����
7b<)i���cP=�=��=箎�8�=�K;�!M�����8��/A��u!��=�!=��F=�8��6��>��>O��>��=�(�r-
>��T�ּZ�^*>��v���b�liu�uŃ��	(�m������>%/U>�h.�`ᒿ:�?Tx>�1 >��?�h?&j>�P���S�KR���A��6{�^��>���=W���I��Xm��R�@�1�>Q�Z>`�>�g�>�/�OwC�Şm�Q�辇2�R%�>��9\	=8#��={��ޘ�T���1�X�����=I?�ȃ�ӥμ�w�?l,o?R|t?���>�;�=��F�mY@��ܽ�"����>����?R4,?`�?��!��Z����텠�V��>�*w��A�2f��n3��\ �����!#�>C
��ؾ�%�R쎿%fv����S���m>��Q?#)�?Ѩ�:����:w��H��S�7��>߻�?�~�>p(�>"�I?�r�<DQ��Η��n6>/XS?^��?�??����=쬴�S�>e?	?���?*��?�ss?��?�9��>��;f
!>G7�����=l>fÝ=e��=hM?[q
?m�
?i���+�	�������c�]�|g�<���=ҍ�>�<�>��r>��=,7g=⪢=�1\>y��>�Ï>��d>ڣ>C�>w�q�߾�?o>��>��#?KId>VVS=i��L��K5>��/��=L�0;��=�~O=�AS�#3���j����>�����?3f�>^{ɾ�+?�߾.�$���=�8�>���l/?�3>и�>6��>j!->s7�=��4>wZ>�7Ӿ��>D��0�!���B�+R�w�о�k{>�M���&��y�����GJ�Ob������i��B��W.=��.�<B�? ���N�k���)�i ��k?�
�>�5?����'Ί�7�>�2�>�Ս>�����y��sލ�'��%��?���?�sa>��>%�W?�?�K)�qH8�i�[��r��U@�мb��a������܁���
�
̽��^?��v?&?@?C��<�!|>�&�?��&�\����S�> 0�ۼ<�f3K=:.�>�u�� ak���Ծ=�ž��5�=>ylm?��?B?��L�bAG�*p>?�@?�;9?�}?��5?M@?�Aٽ�N-?�<Q>��?���>5�G?BK?�$$?��m>a{=!G�Ĕż�����Q��w��xjѽ�� ^�=��=��=�}�;�HM=�Js<T����m���m�<�WS�Fn�<~��=}��=0%>
��>��]?�)�>_-�>p�7?d$��~8�ퟮ�\/?/�:=�悾���Kբ��4>5�j?˫?�GZ?'hd>S�A�]B���>��>�%&>�\>;�>Ć��tD��؇=y>�> ��=�dI����3�	��ӑ����<jD>��>��|>\��(�(>,
��� y��ed>pHS�;��r�T���G���1�ŕu���>��K?h�?擙=�龒k���Pf��)?צ<?�]M?�;?�m�=��۾"4:��J�����>�N�<���剢������:��r4:UNs>�g��Xݡ���b>:��C�޾�in��I�u����S=���ǱK=�W�X�׾[��+��=��
>/S��u� ���۪�УI?T�c=G���X
T��J|>�8�>���>ۡ4�Z6{��@��N��W��=ׯ�>�d:>UL���/�C#G���� ��>IA?Sa?�N�?�炾S�p��d@�C%��꥾����?z�>{??s�.>ϭ=ǳ��L�&�e�L=7�/�>,y�>�_���L�v{��/;��%����>+=�>G>u�?"M?yc?"�M?VS*?��>�s�>�eX��ݶ��E&?���?�ׄ=�Խ��T�R9�� F���>��)?/�B����>��?��?��&?�|Q?�?L�>� ��:@�t��>\�>��W��d��]�_>�J?]��>`AY?ك?v>>cu5��Ӣ������:�=�>��2?�/#?-�?ֱ�>�S�>�Ƣ��Q�=���>��b?{<�?M�o?�M�=.�?/�5>}��>�_�=l�>�b�>�n?��N?�s?��I?
�>��<�$�����Y�o�D6\��D�:p�H<z=�-�Q�v���ƹ�<}ݛ;u����	p�����<�~=����;YU�>G�s>�֕��S1>��ľ?D���S@>w����R�������;�Ӎ�=2Z�>�?qx�>��#�(�=x��>iB�>����(?M�?-?(Y
;�b�r�ھ��L��3�>��A?�L�=��l�?���t�u�s�e=��m?@q^?>X������b?i�]?�[�=�\�þ~�b�����O?��
?��G���>��~?��q?>��>��e��9n�����Cb�a�j��Ŷ=�f�>�R���d��;�>�7?�I�>��b>a�=�u۾a�w��o���?��?A �?���?�'*>��n�o3����ړ�NUP?��>�ё��w�>d�!�4$;h$������|�呡�=���6A���]��w)���p�(�#�Ht���[?�!h?Fuy?:�W?�^��Os�ca��}�g�q�D�@D�w�0����T���A��Dg�o����˾@J���
>�v��3;���?Ƞ/?�*��{�>pȥ�G�
�i̾=�D>�״�-{�I.=�ı�8U<o�<�S�{D�5����?�۫>���>�@?;4Y���7��'��E@���޾��8>�g�>�ي>}F�>�$=�yV�z��2�ƾNꏾK���?Uz>H�X?;R?�-p?-!ѽFG'�7u��$�a�˼�V��C�9>B�>y`�>q�P�T"���'��B��Wr�<P��Ӊ�C���=��(?��G>SǞ>��?m��>$���ܞ���y��A)��e�<&��>=�Y?���> Hn> ;���(�+��>��]?�'�>X$�>�O+�qe%�i���$�� >:��>*��>0�>�=i�Qb��:��^��������%>}�M?{}���G����>�gk?��2��>�ĵ>Fi��:���׉ƾ�\��>�(�>���=2�>b�о�����Ɍ�"�_�R)?�M?*꒾��*��@~>�+"?Dy�>�.�>!2�?�3�>�aþ�j(���?��^?U=J?�HA?;�>��=����EȽ��&���,=q��>��Z>m=-��=���`\�}��m�D=�f�=μ�2����<f�����J<�j�<��3>��wHY�����4(�B��^䵾G����׼ܤt��IN�.�t�]��S=1���=�(;>K����<槾�r<�o��?� @^Z׾�񯾊+ſ3f�hop���>�쎾HS��6����0,��?�Q�پ^����p,��;W��Iq�*%�k�?3���5�ǿ0���O�����?��%??v?����P+�00��>��]<��(<CP뾑����̿g٦�R�\?�:�>�D���*�>WWv>��%>P�d>�-��8̐���<ǉ?D3?�b�>�̘���ʿ�ķ�A��=���?E@�yA?��(�b��sV=���>��	?ζ?>�u1��I�9����=�>l;�?G��?�M=A�W��+
��|e?�4<��F�^�޻,��=Wz�=�=%���J>&Y�>�� 8A�f+ܽB�4>�҅>f�"�ُ���^���<=}]>ֽ�0����?"Fn���\��?L�>����U�<#q[?TX�>U 1=�-H?M~V��<ֿ�Ww���`?�q@y��?�i>?�-���_>��M�S?pS?���>h���'��oRn�l:o=I��A��CDi��_�=�H�>n�D>�Q�{�-��u����78�=�P�
ǿ%�:N�b��<�'8�tM�x�齷���P!T�gY���]p��$㽒o�=]a�=�Q>�>(U> �W>7X?�m?��>�>�i���}��G8˾�2}�����Q�#�E���� ����u���߾��	�nH�Z����ƾi�=�흍=ΆR�v���^m!�Tb���E�0
/?��#>��˾�>M�5�<�?ʾ>.��G���0����̾��1�ݥm���?��B?q慿w�V�x���������W?/��'�����
.�=��żJ=�F�>�*�=V��=3���R��/?
#?lܻ�	��4�2>�V
�ѐc<�+?��>V;|<��>��&?e%-�������S>��$>d��>���>[�>a宾C�2�?R=W?$=�����z[�>��ž+�t��{N=� >7*���ּF�R>9�<^J��C�<�ǽ(��<�w?�$�>[�<���U�A�Y����=��O�i��?"�-?��>i�I?��z?R��=Yt�%J�m��q�2���K?[I~?��=�6n<���:[����A?mʒ?��>w�ž���)�����K�>���?B8?���<�"��e������O!P?B�o?�a�5�����H�����>�?���>+I��c�>��7?���T���*����4��5�?�5@�|�?A7T<zQ<��⼯�?F��>�\ �೬��ֽ�����u�v	?���?4��&�;��Aཪ�P?�'�?E��>uVe�ih��{�=@ᕾX�?��?�|��C�d<����l�s�����<�t�=��<�"�����7���ƾη
�b���yv��)��>;X@��H!�>A8��3⿯XϿ�
��A_о�Sq�}�?y�>��Ƚ������j��Eu�եG���H������U�>{�>Q�������>�{��r;����h�>2��$�>��S�~��C����3<�ے>���>e��>6��1۽��ę?"U��Bοꭞ�u��5�X?d`�?4s�?�{?��:<�v�3j{����<#G?��s?*Z?`l%��]��7���j?.3���R`�(�4���D�D�V>{�2?"�>o�,�n�{=U�>��>�>o�.��bĿ5Ӷ�z"�����?���?@��$
�>��?:�+?���\��D���?�*���Y� p@?ML2>e��
�!��&=�ہ����
?�90?�)��J�]�_?+�a�N�p���-���ƽ�ۡ>��0��e\�N�����Xe����@y����?N^�?i�?ҵ�� #�g6%?�>c����8Ǿ��<���>�(�>*N>aH_���u>����:�i	>���?�~�?Qj?���� ����U>
�}?���>��?5�=�4�>-2J>1�!���l��=Q��>%����h�>k~W?�:?��E��VR�i =��.P���>�����*�L���=��?��s?W
�>O���]�<p���@���پS�J=�q�#�"���l�1�B>]��>s��=?���h)���?����ٿ{c������3&?Ǝ�>�u�>���;����&<@�X?|7p>���Pٵ�q����ؽg��?/j�?��?�8侶�Ƚ#Q>���>ʦ�>}*��ҽ9���̮�>fO5?ݐX���������D>W��?v�@6�?Q�]�b|�>�����O���$T���,�Z���x>y� ?]��R>��>�>9�q�����ׄ~�>���?�=�?��>�z?�с�9�8�L��<�$�>��r?�n�>��$=�2�lC�>a��>���W-��z��&,j?�@�@�ip?���(�p�����Ⱦ�����>�a>KOR>�{5�;�=>֥U=��üP�'>@��>f�>d v>��*>��>�u�=0���z�˸��0���۱V�2�`a�Ns@�"��7���X	���;#�����97R�6�սǎr�_T!�y�1<�4>K4?�_g?Q�c?o��>��e���*>Y �Q�=..��vY>�fY>3;P?��X?�6$?B������h�*慿dP�����i؂>u[
>g��>��>!�>0�A��j*>��I>Үy>�$�=)��<��=��Y=�z|>B��>L��>.��=�5>��>�ᴿ�-��ϔj��.t�����+�?�����K��;��g��������=f�-?R=�=�+���)п�﬿�H?cǐ�����&&���=�.?��V?�A>������a���>]��n�m��+�=���hp�z~(���Q>C�?�03>�Et>*l0�>>9�KM��ϴ��?�>p�7?�ƾ{�[���e���U���澩9>���>>�+�9�� ѕ��ҁ�w�h�|W�<��1?�;?�^���n��ۺ{�D雾EOb>�1J>�C�<��=��f>�!�������E���g=���=��q>�/?�-,>�0�=ϋ�>�ڙ�w�P���>�s?>�*>��??C@$?ty
�_꙽���{�.�V�t>v(�>�>�W>ވJ�HF�=��>5�c>�_�z��@��ZC�UUX>K�{��`�i�v��s=���!��=0�=ھ �ŋ?��i&=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ���>M?��$���W��N������<:��>��@?V���ƽ��/��u?��>Ц�pw���Vǿ/Cs�"8�>1��?|�?s�h�U'��CY-�1��>���?]�P?=>��ھ�L:�*˄>\F?�"J?\�>��#�K\�.�#?�*�?˻�?/>>!]�?��~?�?,쌽V�(�����'����x=�ׁ=[�=�O5>6ܾz .������ ~� �M�p#���>��=�>�շ�����5=���'F��.�<t�>�5>$C>^�[>�?���>\�c>��=��۽�ރ�7��{�K?���?
���2n�PO�<T��=�^��&?�I4??m[�V�Ͼ�ը>�\?j?�[?�c�>M��O>��B迿0~��W��<h�K>4�>�H�>�$���FK>��Ծ�4D�jp�>�ϗ>����?ھ�,���M��MB�>�e!?���>�Ѯ=3�.?�/?F�Z>N�>�3��ʌ���W�m�	?V��>�1�>0/C?I�%?�l����E��,���X���33�[Z[>�Tm?;-?��>ݥ��t��L����v]�yۄ��՝?�T�?٥�<�>?��?�x0?���>���>G��Ҹ�%�=�T>7�!?Y���A��L&����}?~P?��>6����ս-5ּ���}����?�(\?g@&?���P,a���¾-4�<�#��U�(��;;vD���>��>㍈����=�>�ְ=�Om�wD6��!g<�n�=��>��=�-7�(~����(?�8&��X��W=%v��[L���>?5^>�*Ⱦ�^a?0w�_n��ǭ��Cm����Oϐ?1�?��?1˽=bp�<�F?�?-?XD�>KJ����뾎Ҿ}t��;'������">{�>$t��}������3���"��������)���>4F�>�n?\G�>*2>vޢ>^E��S\'��������Y�j��#6�'�,���?h�� �@�Hp�X������ך>��<�@��>n�?�uu>FzZ>Z��>6��Z�>5N)>�ph>�*�>�.>��2>{�=���K���qR?����:�'�����M��DvB?C�c?�>#a�	_������?���?�9�?�/u>ҡh��F+�9?B��>�e���
?��?=��軻�< n��/Q�-Z�����j�>Aֽ�9�}�L�g�f��E
?�!?�>��A�̾�ٽF���5YA=}��?�:?�M�7|U��*j�m`�ߛN�'�������ʈ�
�#��e�l�q~w�<�p��s)�竜=��,?��? (��P �`V��_e���N�X��>���>�'X>rΩ>9>��[:�ץC�����N��?i�o?���>nzI?b<?�}P?�eL?`��>�F�>�R���`�>��;���>��>��9?
�-?a%0?�^?X+?�b>3��������ؾQ	?ޢ?8?? �?�����Oý疗�<�h���y�����c�=��<�׽p�t��#T=�S>�??�CD>5C���#�]t�>g�|?ދ�>�i�>!؉���Q��5%<�w?�k-?m�y>�:������MH��5�>��?��������m�0>�N>sb���%���]n=�꽫�5>ԇ��;ؼ�:�����=�-�=����ڼה��7諾�>�3�>��.?̤�>���='��<�K+���J����=K��!>�v������Q��E���pat�A#y>`i�?�B�?7Q�m�=1�=�]��E�������b���Ǯ=І�>?�?�|O?D�?�[?_�	?�6C>.þ꫈�Zz�jO�� f%?U,?v��>i����ʾE�2�3�1�?�Z?;a�����:)�ŏ¾��Խ)�>�[/��/~�_��eD��|������|�����?,��?�A���6��w�����#Y����C?Y �>�Z�><�>��)���g�%��6;>Ì�>vR?�n�>J�M?!X|?��\?��Q>7�a[��/��9�z�>F�<?���?䡍?�w?(��>�z>��1���`�����;��ŀ�.hQ=6�U>�Đ>���>4��>?�=�wƽ�>���o@�OU�=
{j>A�>.�>���>ɋs>��</�G?���>�_��j��=餾�؃�M�>�u�u?���?Y�+?�J=�c�z�E�"g��,(�>�f�?��?X8*?�S���=v�ռ"���7r��>��>��>54�=�+H=��>�.�>��>\��Z�g8��5M���?�F?�=��ſep���p���8�<<����^�g���Bc���=�F��14%�g����]�~���*����[���F���
��_�>��c=i��=���={u�<�����u<��?=�F�<L$=5s��Q�<xU%�F%���j��j�h�< !K=��L��y�qh?�Q?6H?:�5?>)�=��߽���>n��?G�Y>��>y�����U�~�ܾ�j�� }
���k��WP�W����Q>��˽�<
��=��K>p�=c,<�@w>���=؛ �گ�=&ux>���=�@==���:�=ٿ�<�m?�z��@���[nX��ۑ���3?���>��+=�A�'M}?��=�م���ÿ,k���Y�?gL@���?�3?�"��x��>pa���mS>�7�z:ƽl���1�=��?�e?
?�_b>�f:�:̵�Jy���?�P@HNM?�Ғ�O&ǿ�=L��<v >0C��b5�VCo�D�������ǚ&?�_N�Z-���>/(�������о���=�t+>;��8@�g��t��~�<�a��p���v�=���>#�p>��v=�*[�ۮ>�ῼ��>*>�'=li�<�����뾹jj�=֚.>E>���>��?�n0?"sd?U�>�p���Ͼ����>*�=���>�D�=�A>���>�p6?�C? EK?e�>�&�=�_�>Z�>$�-�_�n�}��̊�����<gw�?U�?"5�>aߊ<q�=��m���>�Df��D<?F�0?�9	?���>�U����9Y&���.�#�����4��+=�mr��QU�]���Hm�5�㽯�=�p�>���>��>8Ty>�9>��N>��>��>�6�<p�=ጻ���<� �����="�����<�vż����
v&�@�+�E�����;f��;Z�]<���;���;��>�>�3�>�%<�YӾȭQ>
�n�Rc��b�=+���Y0V���e�uxx����u�ýtq'>��>��[��q��=�?!�>��->�?��p?R>���>PԾ����>	]���,>� �;谾�RI�Aw�8BK��
����>]��>�>��u>?*�*�=�VH=���E5��^�>O����c� x�q�Uk��ٞ����e��X����B?So��|Q�=�Q?�nK?E�?���>�Ì����cV8>/�~���<���2�y��qx���?�J&?,��>m���B��gǾ����>��3�%�S�S�����)��Y@�>���!#�>ܭ���¾��.� E��]⏿�dB��ap�E�>))P?=#�?��O��|�K��*
�fh���a�>�j?ӣ�>,�?\H?���i+ᾁ���%˛=P�j?���?�?��>���=�0���D�>�-	?��?3��?'�s?��?�p��>T��;R� >'Ř����=��>?��=m�=yh?ɇ
?0�
?�t��4�	�������E^����<Nߡ=���>�p�>�r>0�=xg=�~�=C4\>�֞>h�>��d>���>�P�>��پؗ���
?4��=*m>�?���>�̓=R#:�Ͻ���{֫�*�C���h��<?*=[v�:^�e�������>��ǿg�?���>`�ξ�R?�=����+ u>��d>}���.L&?�ߔ>��4>A`>m�>��>%m�>��j>K6��R�%>n!��,�c�h�֣?�1!��Q��>�������;v쾈H�,bW���d�)H���'i�j��e�I�Y�a=�?��&�a����T��>��>��?^M�����<�=��?K�S>I���Ҙ�&'��ȯ���\�?�C�?�1>�>�K?�s?�����ɾy�{�0I���[��tl���y��W�����U+� 7��K?��w?�\?ȋU��Ҙ>�g�?�d�w׾Iz�>l��z7[�7e=��C>zׇ��7���վ&ݭ��`���<�@_?�g�?W�P? �Q�a�$���S�>RC?� "?Z�{?�a\?��P?���;�J?�~�>�r]?䗇>'D\?��x?Ө?>>X[�<F{	� _r����`;g���/��[��Ko�\o�=��t>4�=sF�=�\
>v��=s���)��;R��=��9=Б=6/>�>�:z>YV�>��\?>Q�>�p>iH;?jR��=C�g��1q?�1=zb���dw��3��ޮ��׽�=R\_?غ�?��d?�P>�8�ՐC��>�d�>�� >�f>��>���h�,���=��>��?>ͅ�=�%8�I7c�>��������ߝ.>���>��C>}���}��=��þA��b�>ڛ���� �c�Z�'?A��A��yB�>I:f?|-?�E#>Teؾv����~|�`VC?�,7?�M?�6�?:V�=q���*�)\����+E�>�?�=| þ���������W�-��ls>A�Ѿh���b>ӯ��a޾�~n��J�@���N=u��PW=���C־�X�Q[�=��	>����� ����>Ϊ�_J?�j=�R���rU�Q��9$>ঘ>�>�f9�wow�ol@�����}�=z��>PD;>Ы���$�|G��4�]��>�qH?�s_?�Ӆ?�p��,_�jT��'��L��5���/?��c>�m?�8�>�>��;�O�d���I�� �>�`�>����G�Oe¾��*����>W3�>8�=���>C~G?��?�ql??�@?�?���>�l���p�&?o�?,��=@Yֽ��V���8��tE�&��>x(*?�?>����>�?7�?�'?Q?{?��>  ���?�;D�>�)�>�+X�^����_>)�J?��>�KY?��?dc9>O�4�U#��h����=ݑ>��2?q2"?
P?Bķ>Г�>J���Kځ=��>�c?�*�?H�o?(@�=}�?��1>��>\y�=E֟>���>�'?�eO?��s?��J?a0�>2�<�Э�t���dr�TjL���;-�K<S
{=<)�7@s��� �<\t�;>*��5&���[�!E������m�;x��>K8t>�����1>�]ľ���Pd@>�#��o��������9��z�=��>��?�ϕ>H�#����=��>�v�>��(�'?R?m7?i�C;�b�OھFML���>t)B?f��=�m��y��P�u�b�h=)�m?�_^??�W�Ĉ����b?q�]?v`��=�9�þi�b�K����O?��
?D�G����>
�~?��q?��>��e��4n����PBb�5�j�u϶=|o�>�S���d�8�>�7?�P�>��b>��=Cv۾��w�Qk��2?��?�?c��?a0*>I�n�2���\ݔ��X?*g�>�p��й?L��)x̾c����%h�O��ݧ�����tk���e��O$0��mq��Y��R��=��?}��?rdo?�L?��ܾ[�m�R���_Lp�n{O�S��u<*��;-���F�|A�O�b����|����jt�|	�=l8f�6�M�6��?�P?�!r����>Jᨾ|���ƾm��>Do��?=�:M��k�%�3>��`Q�*����0�/]?W)�>Pj�>�?�<����<��a�� �Č�>���>�I9>�y�>��v>�=������7�����/���Xn>^�W?��G?�gg?��$P*�i������ߊ"�������=��<>S'e>�v��t]�O�.���:���p�V�����u��8�>�6I?��,>�|�>�ݜ?M�>ns���W��[����"�t��22�>��t? Z�>�x�>39�6��m �>�hw?+N�>;6>9��
-��h��m=�?؆>��r>X��>/MT���r�[n|�?4}�|sT��S|=�wr?��O�_M����>)�k?ä��ͱ�=#��>��N-��(ھ����>���>+�=��M>�,��聽�<{��B��1h)?�v?ސ��cS*���}>�3"?�_�>q�>��?(�>��¾�)��K�?Q�^?KSJ?PA?E��>p�=�u��\oȽn�&���-=��>8�Z>��n=��=����\�H��S�B=gܹ=��ɼ/�����<�첼g&Q<zk�<=|3>�5ؿ,KO���˾�����U�
���\ɼ�'A����뽥[�������u���.�DY�G�[��8����i��G�?"��?�B��꼋��Г�X���D��˹>'�s������0����������â��z��i�O���]��1X��g?�ۢ�#�ȿ���y���%?��&?xXd?���<g�Ȏ7�p��=F�(=�~�<d+�q�<Ͽ*�����e?���> ���4�����>��~>�Rt>�ia>d���+��� ��<���>�.?�m�>�9L�N>ͿUw��-\|<^��?��@�|A?��(��쾃V=F��>G�	?=�?>MU1�YI�����R�>[<�?���??tM=��W�f�	��e?nX<��F���ݻ��=�9�=�@=�����J>�U�>|���SA�m=ܽ��4>م>|"����V�^���<��]>��ս�;��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=X���˿�=�8����D=8vn<����B���m��9"���s��U�~�>��X?=��=�%9>�>�@>;�+>��_?`h?1>�>�>�B�ϲ�������k��r"׽����씽Z쫾�Ծ��ؾ\�
������v瞾�9����=��J�Ï�F��o�d�v�P�P+.?�$">~�ȾwvT�{��<$4׾�8��5�����q���˾nV(�z\e�vv�?c
H?7����Y��s��7�U���S?s:��K���r����	>����=���D�>B��=�q�{.�#�G�'�5?�| ?�nƾC��k'>`�����<�(?�6?����P�>�)?����
��v�`>�}>�ۓ>�)�>��*>+>���u���?��W?�7��݋>�0ƾd�c��,2=Q�>/^J�Nc�"V>\1�<�م�P���㮽GiO<��w?an�>�<���?�Ǫ���sD=��ѽ���?L4?���> VP?�_Z?b��=���[\7��^�J�ٽ��L?K
Z?E�N>X��<q�c겾v�C?��v?�6 >;T��Ǝ�]v����#��>�7x?K?�>�� ��6h��+����#� ?RP?�Hf�����ͷ�����'>?\F
?n�X��(�>�8?�-�#0����>�Q�+�?��@�@�ȧ������=�w?M= ?�"������f�C���tA>Ev?᳆���y�-�9�U��'?]�?(	?h��q��:��=z����N�?l��?�-���s]<����k��}��|�<$�=�/���$�c����7���ƾ��
��x�������>�\@��Y��>� 7�'�yϿ�ꅿ(о��q��n?���>�ɽܣ���j��u�e�G�N�H�:��E��>ҡ�=TL3=�,�-t�<�(�i�����>!Ɏ����>�����=�����6�:=$ݞ>�ߜ>â�>�A�$ۉ�N��?�푾��пq0������$?��?G�?53?��=�^=�v�ic=]�d?��<?��T?�{���Ψ<�-��-�j?k_��xU`��4�hHE�6U>�"3?�B�>:�-�p�|=�>���>og>�#/�i�Ŀ�ٶ�H���L��?��?�o����>o��?~s+?�i�8���[����*�Ǟ+��<A?�2>$���D�!�60=�NҒ���
?D~0?8{�c.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?8��>�x?��-=R;?�w!>�n����>����=�v�>Kd��$��>�D?2?�_=�3����(�sI�3F�����0�K���=#@q?�Z?�Tz>f�~������'��E� rx���>u�ľxC-�����FO.>��i>5M>��r�Ä���>�B:���h��7 ��]\C?Y�>B5�>+�E���V���񽿱>?�d>�������ꏿ����Ɨ�?3�?)p?���}�7��y>�z?p<3
���//>����4��=�8?}��=E!��f�}�CW|>n��?��@
@�?�����~�>�Lэ�`���c��V:�s�@>��:?�x�'<J>���>�=��z����� '�� ��>�ͳ?tI�?%s�>]f?H�_���'�`�=ϴ�>E8?�.	?��b=�ܾ9;O>f�?+H�A����[��~X?�@� @Z�`?����B7���,��!��/s���k�<�+�=���>EJ��@��=\K=��Y=[����5>5�>qPn>��q>ӌ5>k%>9^�=.	�����F�������|l��C����޾��1%������B$��7��g����/w��ʾ�-���j��(�p�)>K� >Q"T?��i?iq?F�>�$���
�>�!	�kI>�����b�>Z�:�)Y?{�?])d?���>�hн��U��ܚ��ߊ�Z�^����>.��=���>�:�>��H>g�ͽ#��<��
>�?>C[=��M=.f9=�>8*�> ��>���>vk3>�C<>��>Fϴ��1��g�h��
w�~̽0�?{���S�J��1���9��Φ���h�=Fb.?	|>���?пc����2H?#���y)��+���>~�0?�cW?�>&����T�,:>;����j�5`>�+ ��l���)��%Q>vl?�ef>��t>*�3��^8���P�j����k|>a46?O㶾�9�G�u���H��hݾ;3M>W��>��D�^d������؟i���{=�v:?{?���ư�]�u��1��HtR>�\>_�=r�= �M>��c��fƽ*H�O`-=�p�=��^>8Q?��+>�Z�=O'�>�D����O��v�>�A>�[,>N@?%?(}�-^������d�-��v>��>���>�Q>vQJ��ԯ=�u�>�a>��s���'C���?�TCW>�{��=_�Aiv��x=@�����=u>�=Q �G�<���$=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�%�>���ř��K��vw�I�<=t��>��E?�����Q���@�	?��?��(2���mɿ�"w�)��>� �?��?��m��U��&�?�o�>B��?4�W?EMi>a0ݾS�W�L��>�=A?yO?�#�>�9���(�?3�?o��?ܰ@>�k�?�p_?js�>߶�=TI:� ����y�|�>d�ƼL�>J�7>zvҾԂS�Xԉ�w���q���E_�>b�=)��>p ��B��	x��&a�LD����ȼ� �>K�C>�^~>jp�>�{?���>�~>�t�����*����G��K?��?Gn���m���<�U�=� ]�1?�R4?\�e���ξ�b�>�\?�ހ?�9[?oʔ>��@>��J���]���9�<��K>���>���>Ɉ���J>JyԾW�D��b�>QR�>�	����پ�끾��t�Й�>�f!?���>��=S,?S�?jV>�*�>�N��k��P�3��=
?K��>ÂC?�.p?h	?�>��������葿�:��a�>#sh?=h0?#��>"�/8���]&������x
�}k�?�{�?�S��'?Ն?5DA?�2?�λ=Ɔ9��9���G=zCn>0�!?����A�L<&���)x?�V?��>�В�}ֽ�XԼ���L��-?�/\?�A&?����0a�vþ��<��"�t�P�Ɨ�;��E�3�>��>���d�=>�}�=�=m��6���g<l�=���>�6�=�7�o�����?�m����5�v=�����{����>��d> �����l?p	��8g��Ѹ��獿�����ޗ?���?:�?��>���m��w4??ވ?�R?�P?�A������m��jO����n�k5<�]�>_O9����?֪�D������I/�C�o�6i�>�	�>a~?�z�>>�>�L�>�6��� �{}о������k�c��%�3�P�-�����╾d�<��m���Ծy$r��a�>�s��$��>�?b�M>�ă>#[�>"���X�>4�=���>0W�>�w~>�&#>8�Y=�ۼ���g�R?tW����'����@=����B?��c?���>�_��Å�z��?�?���?���?e�v>�lh�o>+���?J7�>�̀�m�	?"ZB=�m�����<�������r��

����>�~ԽyK:���L���e��
??~�����̾7�ؽ�ᦾ�x�<LG�?H�?#j��T�T>y���I�:yO��u������"��[�+�vOg��4���]y�$b}�1����G=J0?ԓ?<Y������A�i�Z<k���b����>�U�>��q>d�>��k>��W <��0U��$�Oю����>ʆ{?-��>��C?u.G?�|R?�H?��>�+�>���B��>ꃽ���>Y�>4 H?�E?wH?4A+?�*?X�3>d~������E߾$�?q�?�?}��>c�>B����Ġ���<T �<��N�@ �$��<���;UȽ�b���=��[>ĜR?�>��I�L}��(�>��n?ט>���>�1�������?��/?�1>����0,l���k��>҇�?�qM�W�5<k�4>�I�>y�[�Q��=�/>����n~�=ܙ��Є���@ =ڼU>j>���=��K�ZT=N�ݽ[�#>���>��&?*x�>��>on��\�(/�-�=�p>6�+>P��;� ��揋��0���HZ��ۊ>j�~?v�?8��=P�>��>>�_����;m� �;����&=t��>AV1?B�@?/��?:�<?P,?�9�=��k������M���% ?7!,?���> ��Z�ʾ��m�3�=�?�Z?3<a�t��<)�m�¾��Խ׮>8[/��/~���qD�ƅ����_���%��?��?9A���6�Xw�񿘿\���C?u �>�X�>��>"�)�V�g�>%�Q3;>Q��>�R?��>J�O?DG{?:?\?��M>�6�Ԉ��@Ҙ��@�9��>T�B?ޤ|?�͎?�l{?���>��>8�&��o�������ś｛.}���-=NL>ɽ�>
�>^�>C�=�˽�Ķ��6�:{�=�l>���>8�>���>o>�o6;dH?��>�L��ӵ��<�������Q?�iv?���?� ,?��=V���E�(������>�@�?���?�T*?X�R��n�=�Lɼ������s��K�>��>�B�>��=SP=��> -�>]�>I�����mv8�JJ�&[?b�E?Dv�=@�ѿ�}�����t�1<>�m���R��c�=ꐌ���==�ӽ����h������%��8�򪁾��¾~>˾&��>�,*���l=L�=iU�=p�Z>4�<	�<���<�����ڽY��>c�?�֖�<r`�=�n�<�="9�=g=��Ǿ��{?��H?4J-?��C?�8|>b�>(yV��s�>�"���?R>|�2�2ٻ��4�"���m���ھUkվ7kd�G���X�>o?�V�>��,>���=|�*<�(�=Zʐ=(��=�-7��p�<rq�=<�=w�=M�=NV>s[>�6w?X�������4Q��Z罤�:?�8�>f{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?Ati��d�>M���㎽�q�=K����=2>q��=w�2�T��>��J>���K��D����4�?��@��??�ዿТϿ6a/>
@8>F�>d�R��1���[�E@b�M[�ؚ!?�;�il̾p�>Q��=�޾��ƾK.=8E6>�_=��\�l:�=A�y�VG;=n!l=�>�UD>RF�=諰��'�=.�G=�Q�=��O>���8�7�#g+���1=�u�=Ppb>�I&>Nb�>�A?7�0?/`?��>-�u��׾9���z�>���=��>�T�=Zy->O6�>��5?�=A?�H?���>sD�={*�>��>"�/��[q���ݾ�y����_<lW�?/��?�׳>d}�<u�5�z�<�:��=ܽoz?'�+?�
? Ԟ>������M�"��G*���;��[�<�=X=/�V���G�Yü��������=���>�H�>���>�#�>n2>�6>�`�>>��=A�=f�o=J��Z��;�! �z�.=���eX[=��u�D�=�I���۴��+����~�?f<���<���<�ü�ů>0\�=�K�>�d_=�N�<�N>�%o�]P���&>�����aF�Mo���n�D9������>�a/>5��Pz���?J�}>��>G��?��?Ef�=(E��9v������_�6�V�ھR��>o]�=񑽇�L�x��c��r��-��>���>�[�>�>Đ+�"�:�yp="���E2��\�>xh���ۻC��u�u��g��g矿�d����?rB?[ㅿ@0P=��?s�S?� �?b��>]���L���>�g3��=>��H���v�쩤��$?ɝ?� ?e��V�>��ʾ�˽|��>�J>�]YO��]���	0���c�^���K��>}��o�̾��2�d���G����B���j�W��>�sO?>��?��W� ����9Q��]�*�?@j?� >�?�d	?䪽7��a�l�Q��=��m?��?��?��>9��=L'���V�>�9	?޷�?벑?�ts?��?��l�>� �;u� >ڮ��d��=v�>��=�&�=fp?�{
?޿
?PO����	������e�]�<T�<��=���>�i�>��r>D�=�~g=u��=�g\>�>��>d�d>�>A�>W���a���-?	�O>��h>D�'? $P>ߞ�g�ͽ?�=��$��?�hQL�@�N0��T�"��;*�}�v-<�!�>T8ſ� �?�-�>'�?�Zɾ�ڽ�(;>[<�>S"2�:Q�>m�!>�|u>�Y�>�Q�>>{U>��O>$�<>���e�=����d+�ePb��h3�,���O$%>k~���B4��w�[�2�����j�����u�:6����0�=�=f6W?�F��݂��7�8�^�Հ??��>�l?�̾�ݑ�ε|9�@�>F�P>��˾0����������?���?Y^@>L��>ҤS?�?��8�oq���r�k\��7�NW�Uuo������������O�[?@�b?f�@?��&=ܕ�>�n�?<�'�4��E"�>�i*�} P���=Uq�>�ټ����p��+ǾqQ��|�>��k?d�m?I�?�h�=��<0:a>�S7? �S?ng`?�
"?�)?�|ɾ�;'?���=8�&?�>c9?��?��?ۦ*>���;�	��Z�j𚽔���X~�	�{��S���l���o>~��s��2>>>%4	�J���dI>nR���<��=�`�=�r�z��>@�]?!�>�>�D8?r2���8�r���/?�7=%����|���!��Dp�#�>��j?(��?�<Z?�d>��@�n�A��>���>��%>��[>�H�>b;ｔ�C���=�>��>��=6�P��まH�	����O�<�h >��>�0|>�����'>|���.z�~�d>��Q�a˺���S���G���1�E�v��Y�>�K?O�?蛙=1_�-��Jf�/)?�\<?�MM?y�?��=��۾��9���J��<���>�H�<��������#����:��z�:X�s>�0�����kb>��pE߾U�n��J�2�O=ȑ�?P=2!��,־��g��=�I
> ���+!�C4�������8J?�pn=&���cXT��ݺ�5�>�&�>�>896�L�|�U@��G��@ޖ=nj�>�:>I�����kG�?�d��>*@?��Z?���?���)*f�0�B���R󪾻<��?�b�>?Et->	��=꾾�'���e��!A��?�>.��>���e�H��=��\>��?,&�Xʓ>��?��>�a?�mI?�?��]?� ?�j?w�>AX^��Ÿ���'?��?A}=��׽dd��R:�n�I�H~�>��+?�&����>M�?
v?m!?
�L?S�?3L>���(l;��͗>Z��>q`[���|�h>NXD?�P�>R�`?(G�?$�%>E2�����4-��>�=r�">��4?eq!?i�?f[�>���>(�c�a=>�/�>�qN?��d?~.l?ٹr>��6?�zf>�P)?ؖ�<5,?�t?݉A?Մd?�|Y?�**?Fj�>�~=�tӼ�6�h��0�1<!�.�μ��P��=��W�����9|�9���=����9$a�R-=���<�{�<o�E��ĺ���>�u>1'��(p2>	�¾a/����?>k�ݼ����X����<����=�~>� ?Ty�>_"��Q�= ��>]��>����'?��?��?��D:vb��
ھ�M��װ>�H@?�%�=�vl�A�����u���X=�sm?2]?��[�x���b?�]?g�=�l�þ�b�>����O?F�
?�G�7�>L�~?T�q?��>�e�:n�?���Cb�j�j�Fж=r�>�W���d��>�>�7?�N�>��b>?$�=u۾�w�wr��X?��?>�?���?X**>��n�W4�U��E���l�W?��>rI��P$?BQ��T���[�ړR�R�Ծ�圾ڈ���r������7���Gk�Ч=l?��p?�n?A?����(�h��1���f�~�[��X���)�,���M��I�ɘo�#���d�#PQ�氍>�P�qAA��?֝&?0��a�>𨕾RL�S=ɾ�$G>���.����=�e��@�G=��C="d���1�ܯ���
 ?���>�&�>n\:?@�Y��=�<�2�FI7�Џ����3>�L�>��>�D�>��뺱�1����+ʾq�Ÿ���W>��i?9�Z?�_?	h�%2��J�~��(~D=xdȾ�9�>>�=�ǲ>�"��}��t��o]��qy� ���A������>f�4?�>f�<>�E�?�y�>n� ��+m�jء�s:A�̘m=4?R��?:��>�>�f���I�f�>J�S?��>���>��Ͻ��2�^ؓ�(x�\u>�/�>��=� :>����,R�~���+�k���3��4=��p?��$������"�=��s?y#���k�=۽?�}���<�夾��8>�g=hC?�<�2>���������g��ҾS?&?n.
?�~�1��.U�>O?5��>aO�>�;�?�]�>∙�6�;k�?2sc?J+S?�nF?�><')=m�Ͻ1\�����B=��>;:P>�bK=��=@����Q��N��2=BĽ=��Ӽ�(��x��<�\�6w�<X�<�(9>}�f�s��G󾣇3�|�\�ᅈ���Ҽ򛨾jr�Z⥾�⽾P���>�_�0�����Q�I��:ɨ�S�^����?�@�w�����ک���w��$��CQ�>gi������q ���������þDG����<���h�Bρ��OH�u��>J�D��=ɿ
���(/F����>k�?�X?�;��f��:'��S�=U�ٽ% ������͐��uտ"��N?p(�>�A���F�&84?ȫ>�A�>I/'������t*�?n"<n�?2�4?��'?#�ܿɻ���\C=�(�?��@�A?ς(����֩V=���>�	?;F?>J2�o;��ư�}��>�=�?
͊?:�I=��W����ge?cQ<�F��=���=�ץ=�Z=? �6�J>M�>��@�ܪ۽�?5>6��>� �\���f^��Y�<ν]>t�Խ����5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=~%���ѿ�g%�&�!��
=q��mɼ�o��ѽ��<y���>r����ܬ=j��=wD\>�`>bG>��D>�Oc?�Wv?��>�D�=�J�@��Y엾���=�a��Z�����yT�'�Ǿ�6��	꾌u�����'�T���*C��qG=�JX��;��Z~3��$g�
�@)-?T�=nq���M���w�cM�Ɣ��O�m�G	����H��d��v�?��^?������U�,'����ҽo3J?򓲽�Y.�ں���=�ǽ_�Z=��>�ן���cBC�8�G���;?�m ?�[žх���X}>����	s=-\�>�p�>沤�� ">�"K?��?�N��H)>��>�ȧ>ԋ?b�^>_þ˫�۠9?��f?��R����0X>�>ܾ�>�*ϊ�߶K>��@�#T���8>�9�k�"��ʜ�nd<��r'�f?Bx�>Ɣ4����^��f�i��ț�^\n?�\�>7�/>��-?pq?�86��� ��+�.�뾡!O>�Y?�e?j2�=���|
�Jd��h�_?f��?mO�>v�޾Ng���8������?G�s?��?�L�=ir�A�r��Q���W2?-�h?��p�A��X��c���ք�=�9�>Y~,?�r�ꧦ>�M?��{-��.����\����?ڏ@�h�?v���I����{�=�-?u��>���.�RzZ��Ѿ�"=l ?��ξ!I���8;��N}��@?G��?M?����+�=�=�ϕ��K�?���?OK��/�j<D����k��;��K:�<��=�G�#����7�7��ƾ,�
� ����A��Uކ>SI@�J����>��6�<'���Ͽ녿xyоy�q��K?���>6ʽY�����j�zu�A�G��H�q����u�>�>�����<�{�3y;��>��8�>��/R�>(�S�b赾f����f0<�Ē>i��>��>"o��깽�O��?���a?οE���Xy���X?�T�?d��?s�?0&0<%�v��rz���� �F?�us?$Z?A�$��\�sh6���j?C[���T`���4�dEE�_U>�!3?x<�>�-�&�|==>c��>�c>�"/��Ŀdض�����Y��? ��?jo����>��?	t+?�h��7��\����*��:(�f9A?G2>�����!��.=��Ӓ��
?r{0?Y}��.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�]�>���?p@	>� ?��>�Р��J�Z�'=�>O��U��>YUV?W��>�<=�I�?��8��^D�.g�EC��>�	w?=�O?��<>RK���vļ�D���COH��\^=N�^�Q�~���(���=@{F>���=2Z}��&;V-?��&���߿ޠ��㨝���Z?;�8> 0?k����ק��,�e?<�l>k��>��[����x��y�?!�?_p?b��X.m=����x?��>Pz�����=���<I�>R�(?cf�D옿job����>-��?�W@׳?;F��{�
?|0����=-�����A=⽿��=�J?0h�7N>�w�>��>��x����H���K}�>�?3�?���>��`?e�i�ۏ���<��>k�7?��?�N�<�����az>(�?��پ���]�\?��@�@�Pc?�Ǭ��F��
���񨾕0Ⱦ[2�=��S<L��=�Bh�y��=	 �==|�=�%��X>ޞ�>(�>ҟ>!�9>���=_ے=�j���'��ܪ��ّ�9�3�������>����#�$S#�}^�j���-r�����S��]F{��w���[��m����&='�F?ۿ?拈?W?��epl>�&�rC=`K����>�f���-H?p�|?�5H?��I>@����gj�7؜��"������R+�>ۛ�>��>�Y�>2ό>����Y=P�>(%0>=�b�<��=�ҹ=�ު��U>n��>Y* ?���>��>H�&>�鵿�ϼ�ȁ}�������";�̞?�կ��Aa�;��� -��Y׾@d	>�&*?"�:=*����ؿ�H����K?�D�ٲ�s$��]�<P�$?�4?���=�bq�2(0��M$>�5��̊i�k��=�����H�+��G3>�?�Pf>Wu>ҧ3��z8���P�=���t�|>�$6?Զ�H:��u�o�H�g�ݾMdM>���>QN���������~�Ii��%|=dU:?J�?'!��h����uv��d��;�R>��[>��=��=}�M>��e��%ȽQkH��.= ��=�_>��?��->�n�=ٽ�>�����F:�z��>D>�<>F#=?�'?��Y��5���E1���\>��>ij>�>)cL�̆�=vF�>"�b>�A.���o���R`H���U>܁��SL�'pv�`�}=l����Z�=���=��꽩0:���<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿg�>��$�R˦���w�p{��YC>A��>�|;?{\��^���6G�-��>:V�>O/�����5uڿge�����>�2�?���?-�s�V����:���?��?�5?�t�>�B#�QE���'>��[?�\T?b�>�,�Q�۽<�&?7�?@��?�P>�l�?K[p?�a�>a�>������"��\�2>�Uҽ��=�a>�[���?�ř��R�f�c5l����?-�>�8=J_�>�eU�;�þf��=�~.�[���_eD�3_�>[��>�y?>eH�=���>Y�>���>��̘����{�͡�Z�K?���?����2n�?P�<���=|�^��&?�I4?�n[���ϾIը>�\?n?�[?8d�>G��U>��B迿'~��৖<��K>K4�>xH�>�$���FK>��Ծ5D��p�>)З>� ���?ھW,��d5��xB�>�e!?F��>�Ю=˭!?�a#?=�f>��>��E������H����>���>E?�?z?D�?`缾�2����Ψ���FU��S>t�v?C!?��>W=���3��.û]t�+���Q�?�(i?NB��cT?"q�?�e;?(�9?f>�� ��DӾ�i��3��>[�!?�	�h�A���%�W����?�2?Pi�>Cᓽ�0Խ�ټ����V����?�\?��%?0�� +a���¾ ��<N�!�%O���;��F���>k>V���ش=3>N�=w4m��6�6Hi<q��=.J�>��=$(7�~����?���i�����ۼ��|�`�s�~Z>ĝ�>�]�H�n?sT��Jd{�_G��53���ޘ�a��?(��?
6�?p�ɽ$$x��E?Z'�?$?�C?p����r��s�F�bOY�%��8l�~��>�1��!��{���Ѐ������o���.�_8�>��>�h?h��>X�?>0>�ߒ���3�����a�g�D��X�bN���/�"��ĉ�_�x�C�_����2�W�V�i>�n��P�>�W?�{>�P�=,z�>JQ�<�-b>��^>���>��>"[�>KO�<X^<>�[��L�$�JMR?E�����'���~���S5B?�nd?�#�>xi���������?�?<p�?_8v>�|h��'+��q?MB�>���m
?��:=�J�|�<\�����aJ�����A��>�I׽�:��M��jf��e
?�/?m{��O�̾Q׽��Z�=p��?_�?�>�6�B�MȈ�F�4��?�ca��*��?5����%��>a������r��gt��\�B�%>P�(?��?PI��{a�� ��k��4�@FU>��>S0h>W/�<}�q>�K�~�9��#c����Z���B�?��?.��>�H?��:?�JP?�0H?A6�>^�>C�оG3�>��c��b�>���>��/?u�?��"?��?��#?L=R>�A���� �������)?p�?O}
?_�>R�>�����Ϳ�b���^�=�B��μ��z2<l;��|霽����;�Ó6>��9?�D�=��@�pz�c�>��o?Ɍ�>x-
>�_�����`���;?K��>�T�=;����b�l�@�1?˿�?DkH��1���"�>���=�ͮ����=J����u=X,�<6��oD��Dھ��RE>�n���<<􈄽;�<ȟ���P�>��?��>4H�>�Ă�n��=����=�"Z>��R>0�>:�׾Tq���㗿-�g�'�w>-z�?1�?�,�='��=@)�=I�������)��yx�����<LA?*�"?�HT?���?��<?9�"?�Q>v��Ғ�,�����-+?;�+?���>���˾�����3�٧?.W?� a�����5)��¾�"ֽk�>�B/�E=~���ID��}��2��-��~w�?�ڝ?�[C�D�6�)��'����ȫ��_C?mC�>W}�>45�>�)�Ah��7�*;>��>R?|�>��O?�z{?#�[?�4U>*8��M������u;��>L,@?q-�??ox?�H�>r�>55,�t�A�����!�������7_W=�aY>��>LH�>�ة>w��=��Ľ�X����A����=�\f>���>q��>I��>aCv>�<��L?b�>4���� �3��)v���6	�}W~?揑?�1?�ȭ<F��N"G��F�{i�>"�?�}�?�,?<,$��O>�4�<a徴V����>�|�>Lߞ>��>^�e=�=�\�>T)�>����%��i&��)�4?F9D?�>݆��@�p��g]�������;)~o��H��a���:�Y��=b���+���?��twH�sV���(���'���]������#?�"�=t >^ �=�Oe<K�K����NF<�R~��[O=5����0=V+��S,!�̼��]�8�p7i��.:=]��<�����{?�"N?X11?�<?5>~�#>) �hӔ>,
��x?�Ʉ>_#��վM�b�rg��������ھ�	��3�o�\ǋ��,0>�z��V:	>�!>���=��i=�=(O�=�l�==�7����=�C�=��d=D�=CAF=4w�=O��=�6w?X�������4Q��Z罝�:?�8�>�{�=��ƾq@?v�>>�2������{b��-?���?�T�?B�?Ati��d�>I��j㎽�q�=R����=2>l��=�2�S��>��J>���K��E����4�?��@��??�ዿϢϿ4a/>H01>3�>��Q�7�0��Y�h�e�(rX�5z"?c�:���ʾR�>�Y�=��߾��Ⱦ_)&=��4>�ad=}/�9m\����==��+6=�r=��>c?I>���=��o�=]>=)��=%T>��Q;�|����e�3=���=q�`>_$>Ɛ�>�?[0!?�Z?�s>z�N�� ��GȾ��y>��y>�%�>�
�=�C�=��>,2?��?��H?v�>º�=�|�>�i�>Jk'��_�����q�ް����?_?�?�ۘ>��= )��+b�ST5���L�&?e�,?�)?_��>x��m����'��1����� �4���Y=iI��j����<���ý� >��>iH�>��>�y^>L,>/&'>�X�>�k�=R6Ǽ�3�<��e��T�<�u�=��>2���,�=C�4m#�G����,҈�V��=��д�<�@=��<O�>�"�=Ψ�>~�,=��$p�=G�]�Z��z>�^����X��fi�J.���w0�أ �mII>��l>{���@��p?�>�ko>���?6<p?.	>���F�1�Cߘ���J�d��$G>c�=�ݽ��T�l�{�&�M��x��>�ʎ>�Ǣ>M{n>.�+���>�os=nQ��5����>��������1q�O���П�a�h�e��	�D?o(��\��=��}?�I?��?+�>�)��IhپZ�.>H0��$
	=���5q�@œ�\?B�&?%�>$쾞�D�g�ɾ�黽�}�>sME��O���Uu1�j"M��C����>�_��c|Ͼ��2����������B���m�Z��>4O?�n�?�9^�X��P�#t��q����?�<i?L��>�?��?�h����~��a�=w5o?N�?5�?{�>�S�=+_�����>a	?Ȁ�?j��?��r?M�@���>�2�;h >�����/�=�
>cq�=�H�=�/?�
?6s
?�$�� ^	�����v�]��<sc�=&Б>y�>�Ns>J^�=ϥf=��=��]>���>�Ǝ>>d>_��>@�>Z4׾����7?�W�=���>A�0?�|�>��S>�;�<��ϻ����d��$ȶ��������oX&�*7�=�=Pb"����>�k���׊?X;>R��ֹ-?X�Ⱦ��n�GP�>e�M>�{��?�r>�m�> ��>�y>2��=�X$>CK>�־UL>���g'��L��T�T�ƾ�|>.���
�Z�>M����yR`�$��[��sm�ڄ�z|D�%$�<`}�?����j� �
��n�	?Ȍ>�7-?/�m��
��`v>u|�>X�>��\��!䍿��ܾ��?���?��c>\ߞ>_kW?$�?;�,�I�2�y\��;t�b@��kc��Ra��㌿�_��y~
�� ŽE�]?�Xw?��@?4��<Ƥ{>�\�?0\%����!`�>�u/��B=�{�A=��>'=���Qi��&Ѿeľ�i���?>ͽn?�A�?�?w�N���a<3J�=�aQ?�<?�K?�?�X?�蕽�K?Ϧ�>�*e?��=���?�w?��Q?�?��%>�\�_¾} {:W(G�;k��Lj�Y�x��>�=> �=^C9>b�/>1�
>���=$�>>r=�4��z�=���=�@�=�.n=�'L>�3�>3�]?���>��>��7?�����7�W����D.?��=�?��mU���̡�~���P]�=ifi?�?�?wLX?�<i>AlC�h�>�?s#>)�>��#>�Y>�O�>���/C�H~�=��>&�>wȮ=0�V�<d��������*�<��>���>��|>✌���(>ɢ�m�y�dDd>`IT��&��8lU�ֽG��1�}rv�Q��>�tK?�?`ؙ=�����):f��)?K�<?�pM?DO?<`�=�l۾	�9�i�J�/��ؠ>d�<���������]:��4:$�q>r���Π�[mb>�Z�{޾�qn�~�I�t��{J=E�K�Q=����Y־G~���=�	>���6!!�y
��U����J?Fl=�N���V�es����>�ޘ>�Ϯ>�^9�[|�ND@�>����=P��>Ū;>����/�qG�av��,s>B?H�h?��r?$��a�Q���[��}�~���z6?v�@>�?�/6>ܠB=r�˾"�V�i��	]�M��>���>�\��مV��1}�ިþ[����>�l?A-�=�8�>	qI?��
?�l?�"<?�*?&�>'� �a��A&?���?�=��Խ[�T�99� F�<�>
�)?�B�.��>��?��?��&?�~Q?�?��>� ��<@����>�a�>�W�Yb��3`>O�J?%��>?;Y?�Ճ?y�=>�}5��ࢾ�ҩ�@t�=�
>��2?�2#?M�?b��>��?��]�R���>�]?L2�?��o?���=V�>���=�G�>�ic>Z�>���>L�?G7,? �w?�S?sy�>f$<)�Ž�~��$.�C��<4����5=�'�<NZL�Dh�]s����=^&,=K@��=����/��ק�O� ��ɧ<�W�>�w>�2��\�8>"��J�����>>�,
�"z��-f��$#9�Nt�=�g�>�< ?6�>5)��e�=�<�>D�>Z��#�&?n$?^F?з+���`���۾N[��{�>�;C?�G�=@xp�����:�r��9=!j?�9[?B8X�������b?��]?+�P=���þr�b�]S�~�O?�
?]	H���>��~?��q?M��>��e��6n�/��:Gb�>Jk����=u�>�E���d��@�>ɘ7?�;�>��b>!l�=P{۾״w��Q���?0��?��?k��?�)*>��n��4�����ao��]?M��>95��T�%?���J���w��
s���ž���D)���d�������b(��!����G�y=�?T�f?T�k?��I?�<���g��F_�� m�X�L�f�̾=�1�*-:�L�Y�YT��s������{�K~x�w
>q�����=��в?ϋ:?��c��>}叾��	���־�!|>�uɾ�J�*��=������<ga;=�g]�A�����d�?���>U׽>S�8?�<X��8��N&���7��8�d�d>p4}>3h>\x�>�<h�3�=�Ö���H��+o���e.�k�c>�nY?8�R?��{?��O�$��CV��3�ެ���ym)>���<�>�\D���P�A7�VA���k��S
�ڞ���H����=�z?h{9>q�E>>��?��?qm�14���wh��a ���<�[�>��V?���>�&>�YH� 6����>�h?��>�>�ܽ�q,�>��ȱc�G�?�e{>���=�|>.hM���A����NS��}jL�=�">� k?��v�~|�)p�>��h?�B*������>q�<yFE�\sھA!Q�Y�>��>��f�-\�>�΋��@��X���\v~��-?�x?�k����*���>�~%?��>�2�>8�?�c�>G���,�=:f?�W?��I?@�9?���>p�=�_��E�ǽH�%��Y'=U��>-�d>���=���=G�)�"�a��.��=�=>�s����)UP<d	�B�;Ϛ�<�$/>����k��v��u='���۾B�ξ�Mӽ5���ǘ����n�|յ�����]#=�Q&=RX����M牾=�L�1��?���?=���;ݾ�p��gD�� �Z��>m +�[�G���������?���Z���'��n3��O}��X\���E�F��>�m��˿	����m6���7?��[?��b?{}ؾ�yL��i�>yk<�=�Ex>�ʾ)�����Ͽ�.���3l?R��>e�˾l�)�vI?1?'�ۢ�>�"�<3��d�o�v���I��>� ??,M��G�ֿ����5U>Bz�?
�@u}A?��(�'���U=�p�>V�	?�?>1�0�r��찾da�>�>�?��?�N=�W�z��S�e?'5<Q�F���ڻ��=k�=*�={u�n�I>SZ�>����A��&ڽ4�4>��>��#� ���2^����<�]>��Խ���5Մ?,{\��f���/��T��U>��T?�*�>O:�=��,?X7H�a}Ͽ�\��*a?�0�?���?%�(?8ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�߅�=h6�ˉ��z���&V�z��=Z��>c�>��,������O��I��W��= ��7ȿbE$��4��C=9*����X�v���|���cH��
��(u��,��T�=�a�=3X>B!�>� R>��X>[R\?��l?���>���=9������L��)�;�����0!��̋��o����ut达i⾍�
��k�>�,Ǿ�]=�!�=2^R�Đ�� ��a��DE�[�.?�p#>
.˾�(M��/<!�ʾ������t��¥�.;d�1�1�m���?�cB?���{W�"�����o����W?�����a���L��=�̴���=��>�9�=���P@3�R�R���G?��?h_Ҿqjl���>v)�=�w >�?��>��l�$��>��T?]Q���~��>�~`=<��>�_�>-/U>8t̾"�Խw	8?��O?�$	�eS~�y��=����o�&�j���W�=c���к9|j>���3`������X��;{Bd?���>!�1���IPz���=v�'=4�?�I?��>��^?j9[?��H�������,����m�T>C�_?n�\??��= q�R`�A���nA?(z?���>p�ǾLr��;��5쾾h?Dys?�M?���<�W������ƾޤ?��k?c\���ם��$��Ӿ��>�(�>�j�>3����b?�U?�Qv�"����g���C;���?�P�?b�?�!�H�̽ڄi>�-?͍>�����;���r=}$��� N>��?�܁�d닿apI�wӾ�VG?���?d�>��A���뾃��=:ؕ��R�?W�?	;���
j<���Ll�Ρ���-�<jl�=@��R�"�x���7��ƾ�
�⮜����q׆>�N@>�T��>2�7�c8��VϿ�慿о��p��Q?�H�>%�˽��x�j��u�e�G�4�H����z��>��>Tm���s��L�z���;� 0ؼ�1�>��Լ�>-%X�e.��%-��U�';?��>6�>�@�>n*��z~����?F����ο�,��e�� Y?�&�?A�?^� ?7_<j�^�S�l��{��l�G?,�r?�Y?;��vG��7K�ݾj?Jc��ZV`�Ӎ4�IE�U>!3?�C�>�-�K�|=�>���>e>6"/�O�ĿIض�o���U��?���? n�l��>[��?^r+?�g��8��Z����*��0�?A?/2>,���n�!��/=��В�.�
?�~0?&u�0�]�_?+�a�N�p���-���ƽ�ۡ>��0��e\�N�����Xe����@y����?N^�?i�?׵�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�j�>K�?���=�� ?]�>� �������=�->�/���>��F?Z��>�b�=�>=��v0��y:�]�C��1���	G��~�>/o?��N?��
>��ʽ����.�]����KǽS%μ����y���ɧ�m~�=o(>˵�=�E���ܾ��?�F� sܿhq����V�u?�>�r?� �i?��IB�=�w[?i�e>�HӾ����1!���D�S�?��?_
?M��D��M�=*�?�o|=�گ���I��l$�K{�>�8?�>������d��
>���?��@$��?}��O%?'��ދ�Z(u�E ��U	��S�=�;?Ȱ��yq>E��>Ef>��p��֡�͓y��> V�?:;�?���>�+g?�k�v�1���<Zӱ>ɅJ?!+
?TѮ��l�����>
n
? �	��׍�u7��bc?�v@c	@��`? ~��zRҿ:���w��������=�=1�#>�̽��=d�Q=��4;�@ü�->��>�w>�̃>��8>u#(>�>�I����#�{��������[8�g���<�N;����Q��=��m��,�Ѿw���PԳ���O��&I�}+�C5���=�k??��{?��g?��?-3�iHC>F}�zt�>c�E�R��>�����t?ƃ? �|?��{>������s�ĵ��hkc���Ⱦ�BY>x�>=�?w��>��'>rY�=�qN>Q�>U�>��=�/�=Τ>���>=��>6��>�ѳ> ��>�@ >���=@o��Τ���k�Y :�`H`=��?���MsN�ͦ��!�������,>�0?���=�[����ʿHq����Y?�TY���#�#��e�;�,?�[?��%>Њ�������u>�����^G�{�>X�l��(�8���>�T!?�f>�$u>{�3��c8���P����Dj|>^36?�趾�K9���u�B�H�Zݾ�<M>ľ>�HC�)h��������zi��k{='v:?΄?0���Ѱ���u�4A��cPR>&\>�=/��=�M>=�b�f�ƽ�H�8%.=���=��^>��?��2>�E�=�
�>���m�C�,R�>��>H#3>�/<?O�"?i�=��%���\����3�ٓc>Ғ�>��>˔>�'R���=�T�>n�h>�K?�9t���*yA�R O>[;��I^�Y)��*��=f������=���=�b
� !B��6=�~?���(䈿��#e���lD?S+?_ �=�F<��"�D ���H��G�?r�@m�?��	��V�?�?�@�?��H��=}�>
׫>�ξ�L��?��Ž6Ǣ�ɔ	�/)#�jS�?��?��/�Zʋ�<l��6>�^%?��Ӿ���>/`��������}�z��k=���>D�F?���G����;�0�?�9?�龓t���ɿ��v�(�>�@�?+��?Q�l��ę��9;����>,�?�Q? g>zܾ;�Z��,�>B?�P?�>�>C\���&�͘?�?�?�?'�9>��?�uW?�=(G>�}5�껾��Fc����>��'>������<�{��<�"�Z?����{�i�d����?*�>5W=�o�>��H�eh۾��W�}Y�����/I�Û?-�C>��4>��(>=5�>�|�>�>+��h�������	�^�K?=��?���3.n�7A�<Q��=/�^�k ?uJ4?�c\�O�ϾϨ>U�\?�?x[?b�>���>���鿿�|���ʖ<��K>y7�>qK�>����0K>>�Ծ:$D�Ws�>�֗>涣�:ھo��Q��$K�>�d!?2��>�֮=� ?��#?|�j>���>�=E�c6���F����>���>~T?ۍ~?��?)��M]3������͡�Wb[��1N>��x?2[?���>����:���x�C�t&H��?��ू?�g?��彂#?w.�?�X??աA?,f>z}�n�׾+����ڀ>��!?����A��M&����~?Q?R��>{4��H�սDּ-���}����?�(\?�@&?v��b+a��¾$6�<�"���U����;�iD���>@�>Ԍ����=>�հ=GNm��D6���f<Im�=��>'�=B.7��v��q?���f҃������i���x�0g>@֢>�	�j��?���Cۀ���ÿPz��,_�C#�?�R�?��?��zw���V?K�?�X�>�?\���n�ھi���y�N�۱��)�y�9K�>D�D���ƾo���mm��y[��+�S�N�|�͝�>�s�>��?L�>�w=K�>�@��Ѱ�?wξk�۾�=p���澺+2��f�^����L���S�;�r˾�N~�
> ڄ����>x|?Q�i>+�V>f�>������>��y>A��>��>n]�>`��=ٜ���iý�	�LR?������'�;�辠����4B?Lmd?D�>
�h����������?Ԅ�?Pn�?u5v>8}h��&+��l?>�>{#���m
?�;=�q��B�<fR����������\��>}9׽�):��M�8_f�#^
?�'?�{��+�̾V׽������+=N�?�"?����E��k���C��J����=7]Ծ�cH�F�!���p�s�� QN�\�q�,���>��'?;�?�	� �5QH�����d�S)�>�?j�>�Ҽ<v�:=��0��}5���h��u��G@S��|?�Wu?�l�>��G?�Z8?�mU?��D?v�>Ա�>q��^��>G�� ��>�g�>(9?�##?u"?Ic�>}� ?�"b>0��5��ֱ;��#?�?�\�>3#�>��>���"Ľ@_~=f���d���^�S�w��=�AԼ�	��%ƽ]�=_�'>�Q:?�ĺ+A�oK �fP�>�L?S1	?�>��9�$7��ɼ�<nA$?��?$>�`���Rc�CǑ��
?IXi?ش;�~����&>�>ta=���3�=��`��^�<�B�����c�p=`>9�o=�p���?<�Ͳ���\��C=���>X�? j�>j}�>��~�������lB�=�|[>�U>w�>�M׾󫊿�^���Th�|dw>���?>��?�U|=�R�=���=-Т��/¾���0������<��?3�%?�]S?�ݐ?Z�:?�"?3�	>��S���2��������?�,?I}�>�����ʾ��Fy3�X�?:T?3a�����9)���¾��Խ��>|]/��4~�	���D�(}�\��<������?���?��A���6�͇�!���`��K�C?��>�X�>��>��)���g���ik;>̇�>IR?�o�>^�M?�%|?��\?g�^>��6�{1��Lᘿ^&�9I3$>��@?��~?��?u�{?f��>�!>��1���p����(��b�k��0�E=)�]>#/�>��> �>��=���諬���>�|��=��l>�s�>�C�>�c�>ɭw>R�<@T?{��>0/���'�������/� �A�?_��?��4?��5=���K�N��u	��S�>6R�?W@�?a�'?M&�d(>��<X������r��>�F�>�ޯ>��#>P�=�R�=?�?b�Ž�
ᾙn��W�~�?�b?<1�=J�ſ�%q��m�����5|<�{��Fld�����sK\�u��=T���c������*\�MN���ْ��o��H���.�z�l��>ϭ�=���=<^�=
��<2�¼r]�<��C=xɋ<�=�;y�-�<��A�����̊�)!��L`<�H=����4Ǿ��{?�SJ?�Q0?9�??�5x>�n>%����>/6}���?�B>ߎ�l����kB��
��<闾�C׾�@Ծ��g��\>7�T�Ň>B�>k��=�g�<��=#Ol=�[�=��� � =#B�=�A�=�Z�=���=�P�=��>j6w?\���߲���4Q��_��:?�8�>E|�=тƾ@?��>>�2��旹��b�-?���?�T�?��?qui�Fc�>_���ێ�Vr�=�����92>���=��2�'��>�J>8���J������4�?^�@E�??�ዿW�Ͽ�b/>w3>�V>��Q��31��RZ�c���X��!?��:�ޘ̾�8�>��=�OݾvlƾȞ4=��7><�e=L���x\�m��=����+G?=�r=`ĉ>�H>Y�=6��a
�=�O>=�_�=�1T>�";����>�)=�B�=~�_>"}$>�`�>w�?q0?�gc?U��>�p��Ѿ���j��>~X�=?\�>6��=W<=>�r�>�K6?aD?��J?���>ڥ�=�>�ө>	-��Sn�R�⾏����e_<@��?�#�?�>���;��B����U�=���̽��?��0?H	?AΟ>Q��4d��v�"��~�;5{�1_K�=��DV���T� ^��q��̨=6��> ��>���>8o>!��=/�9>���>�)�=����
7b<)i���cP=�=��=箎�8�=�K;�!M�����8��/A��u!��=�!=��F=�8��6��>��>O��>��=�(�r-
>��T�ּZ�^*>��v���b�liu�uŃ��	(�m������>%/U>�h.�`ᒿ:�?Tx>�1 >��?�h?&j>�P���S�KR���A��6{�^��>���=W���I��Xm��R�@�1�>Q�Z>`�>�g�>�/�OwC�Şm�Q�辇2�R%�>��9\	=8#��={��ޘ�T���1�X�����=I?�ȃ�ӥμ�w�?l,o?R|t?���>�;�=��F�mY@��ܽ�"����>����?R4,?`�?��!��Z����텠�V��>�*w��A�2f��n3��\ �����!#�>C
��ؾ�%�R쎿%fv����S���m>��Q?#)�?Ѩ�:����:w��H��S�7��>߻�?�~�>p(�>"�I?�r�<DQ��Η��n6>/XS?^��?�??����=쬴�S�>e?	?���?*��?�ss?��?�9��>��;f
!>G7�����=l>fÝ=e��=hM?[q
?m�
?i���+�	�������c�]�|g�<���=ҍ�>�<�>��r>��=,7g=⪢=�1\>y��>�Ï>��d>ڣ>C�>w�q�߾�?o>��>��#?KId>VVS=i��L��K5>��/��=L�0;��=�~O=�AS�#3���j����>�����?3f�>^{ɾ�+?�߾.�$���=�8�>���l/?�3>и�>6��>j!->s7�=��4>wZ>�7Ӿ��>D��0�!���B�+R�w�о�k{>�M���&��y�����GJ�Ob������i��B��W.=��.�<B�? ���N�k���)�i ��k?�
�>�5?����'Ί�7�>�2�>�Ս>�����y��sލ�'��%��?���?�sa>��>%�W?�?�K)�qH8�i�[��r��U@�мb��a������܁���
�
̽��^?��v?&?@?C��<�!|>�&�?��&�\����S�> 0�ۼ<�f3K=:.�>�u�� ak���Ծ=�ž��5�=>ylm?��?B?��L�bAG�*p>?�@?�;9?�}?��5?M@?�Aٽ�N-?�<Q>��?���>5�G?BK?�$$?��m>a{=!G�Ĕż�����Q��w��xjѽ�� ^�=��=��=�}�;�HM=�Js<T����m���m�<�WS�Fn�<~��=}��=0%>
��>��]?�)�>_-�>p�7?d$��~8�ퟮ�\/?/�:=�悾���Kբ��4>5�j?˫?�GZ?'hd>S�A�]B���>��>�%&>�\>;�>Ć��tD��؇=y>�> ��=�dI����3�	��ӑ����<jD>��>��|>\��(�(>,
��� y��ed>pHS�;��r�T���G���1�ŕu���>��K?h�?擙=�龒k���Pf��)?צ<?�]M?�;?�m�=��۾"4:��J�����>�N�<���剢������:��r4:UNs>�g�������_>������M���9����d
��g���Q4>����9m�ñʾ�j�>tJ
>Ε���x�삗�J����c?���=^.ھD^�K���$Q>��>=�>^��W��[�D����I�S=˖?Bf`>�_��"��G�����ӆ><F?6�^?�;�?�_���=t���A�D���ޢ�:��m�?T�>��?�:>�=�����h�r,e�E���>���>P����D��3��c����"��3�>�Q?<�(>.?�P?K?@"^?#Z)?��?4Ï>�f��yR��B&?)��?D�=��Խ��T�Z 9�AF�A �>v�)?E�B���>q�?��?�&?��Q?��?u�>�� ��C@����>iY�>��W��b����_>��J?͚�>_=Y?�ԃ?��=>I�5��颾�թ��V�=@>��2?�5#?E�?���>7��>A���i�=*��>X�b?k;�?.�o?a��=z�?�2>;�>~�=�n�>�l�>�?IO?��s?��J?j\�>^:�<��,O��@�r���P��x;�A<;fx=C��z�s�!I���<�u�;~巼n����－]D�i?��=7�;Ϫ�>k$t>WS��4W/>�?ľ�ڈ���?> �������5���8��u�=���>�	?�'�>��#�p��=uļ>q2�>���(?7'?�?Vc<;��b�s�ھ��M�hʰ>�aB?Dd�=��l��T����u�k= n?e^?�Y������g?�K?x���G��՝���+�Z����v�?��?�s�����>���?q�l?u�	?��G�+ք��E���$�����U�=<ji> �Ͼ��u��6�>I�J?���>�>����̾�j�Xd��[?���?���?�ۇ?h�=��.��Tؿ�+���Y�b?���>o꠾FA-?6%<5bھ�霾�<v�Jݾ噣�����>͕��s������jn��?���"�=a�?Mo?�lr?[	[?����Pd���c��L~��X�u������-C�;E��@��h���>i�/�~���=�r�ɹ>�{��?=�$?G�)��0?���N����ؾs�X>�盾�a
���_=䘽=��X=�9T�h���2���l?SU�>��>XA9?K�W���=�	6��9�( �G�9>��>�;�>�'�>�3���S-�;ܻ�������\�"���/m>��h?KJ?n�w?���b7��U|�r�$�|��Hž��a>y�=���>:z�^4<��s&���>�u�/=�	q��	~�x"�<�;?�_L>��e>��?= ?�����@QL�w�2�PQ=�.�>�b?5I�>r�d>�Oͽ��
�!`�>٪v?i��>p��>Y4�U$��x�g�:���>$�A>v��>��>b� ��^�����N"���~(�֠l=�tH?4t�OD�`�N>�R?/�=-\x����>Ldؽy�3������^<��>u�?4^�=��/>�ԾC�.��.}���T�_T)?�H?�˒�,�*��>~> "?�c�>�r�>,�?��>�Kþ���?��^?�@J?:A?d�>��=ȋ��XKȽF�&�U%-=���> �Z>)*m=}��=N��O~\��1���D=O�=��ͼ�X���/<������J<<��<�3>��ҿ��B�%�־�"��������~l��y������]���7���p�u�o�B���}����!�6LN�m~��N��_X�?R��?������Z���! d��fp�̺>k��N=�<\'��R�W��߾뒹��������z9�(Qh��Fg��{)?Tר��Hǿ������3?��D?V�k?�z��A4�S'E�Z��>T��=�<S>3������Xd¿aC��W$h?-��>����K���j>��>�K�>�{Ѽ��>�X��n�ֽҎ?j��>	�?�����%̿9���M?=,�?�@�|A?��(�(��nV=��>��	?X�?>�T1��I������S�>�;�?��?�|M=��W�|�	�e?د<��F��ݻ��=�E�=�F=^���J>�Q�>���WA��8ܽ�4>dم><�"����O�^�-��<��]>�ս"5�����?Go[��*I���<�p�����=�wW?�؟>��&>��J?BV�;{ǿ�zV�^�h?џ@���?��)?��TG�>�澙�T?SQ;?6��>���]��V�=t]	��U�����ºf��C�=Gi�>OmN>��սɋ��R��������>�8���Ŀ��"�F�;�y<��)���y�j����x��ݦB����q�h��ҽ�Ռ=���=<U>�o�>�Y>UmQ>�Y?z
m?\��>F�>��=��Y��q]��ig�F,�����>e
�����i龆�߾	�7�~��� ˾��<��\�=�Q��'��h�'�1`�2�<�ݶ'?y@>�ֿ���K��c�<Ѿ�\����������$Ǿ�0��n�cL�?�D?�Æ�+�O�=�b�Ӽ��μT?B������{��~�>�q���o=QP�>���=>��:$6��V�J�0?I?ـ���/���	+>� �2"=�,?�g?0
;<���>Ώ%?=w(�h��	]>��1>���>G��>��>d/��6(ڽS�?%dT?;� ����]��>CԿ�Oaz���n=�>?16�����IY>�֜<t���>IK�H���7�<�(W?X��>Y�)����b��}���^==Z�x?v�?d*�>�zk?��B?�ݤ<�d����S�� ��Gw=��W?�(i?��>����оȄ����5?��e?��N>rZh������.�?U��$?(�n?�_?rx���u}�������m6?�yx?59a��b��P4
�^���T�>��>,�>}x%��E�>#RA?��Ž\J��'���ϼ0��ϝ?;� @.��?0	<=T����=�k?Tκ>ӡ��1r�gqx����x�=�?t���ۿ����G�Z��<�^?-�?��?�������"��=�֕�y[�?;�?�}����i<���nl�b~���4�<л�=��"�D���7���ƾݵ
�o����A�����>�X@�I轾+�> ;8�'6��UϿ����eоTq�<�?�h�>��Ƚq���|�j��Du��G�"�H�����n�>�>Rڞ��Q��+�}���:��j'�U)�>i���נ�>�V�X
���Ģ�X�<�4�>���>��>\"��?����P�?Y(��U�Ϳc��W��u�W?�?1��?|?�K{<��{�~�q�wE����G?�r?�W?�/���d�?Z�H�j?9l��\`�(�4��;E�#JU><"3?�<�>_�-��|=�4>M��>�h>�&/�F�Ŀ�Ѷ������ �?���?�f�7��>���?.k+?�f��5���Q����*�dr �>A? 2>������!�n4=�5����
?׎0?0}�V9���_?��a�~�p�B�-�� ǽQ١>��0�a\������z�0We�5���Ry�{�?p_�?o�?n���#�a5%?��>?����&Ǿ�C�<�l�>��>�,N>f__�7�u>s���:� V	>v��?O~�?Pn?����6���U=>u�}?`��>�wr?aԯ>-�>WST>�:���﫽^��>h�>#M;<�C?�S?��?��=An=6 ��a�ޙF���3�s�;��%_>Μz?SiK?�/>)AJ��n=}fJ��u��Q8�=E޽I�p��ݺ=�xQ�')>Țv>��>YU��������,?z]7�`8߿Kۍ�[��hiX?	��> 2�>l��_g�*O�<�8f?|��>����������(Q*�6~�?C�?� ?Nƾ5 i����=���>騋>]��.��d��V�>��V?E�$��Æ�����u�>ɛ�?m!@	��?Z�/K?��
��W���{�H�ﾪ�ҽ�
>}�0?��>���>H��=�k��z���v����>P`�? �?gF�>�Ad?ղa�ۼ0��^�<���>>r[?��?D�~����/_>hc?WB�đ��8�	�-Os?�r@�@�S?�L��)l˿�Ĕ����zо�ʈ=��={�>��Խ���=�f>�=��v=�d>ڤ�>z�J> ��>�Z(>諊=ê>�x����#[��wv��wA�k'��d��`7��%���+��%����P�ؾ�|����`B�+���b����<=>�M?��i?�lZ?I��>giֽ<>n�Ҿ�
=r沽��=��>;RQ?��=?��3?�1=/Ѷ��Te��݆�f���t'�����>�f>ֽ>@˯>���>
`� >�4>0�Q>O��=�4�=6��;K��<��4>?��>���>�>/>B>gm>�
��ے���H|��`�jY=�?}3N�pT/�l����)�lľ�@U>��)?� �=�����ο+�����M?M�����j�7��&4>�7?�iI?�IC>�T��{���x�=}����[����=n]��T��w<.�	�Y>�{+?T�f>pu>c�3�X8���P��s��x�|>�*6?�ö�v9���u�z�H��lݾE�M>=ƾ>ID��l����l�7i��+{=�h:?m|?�벽���� �u��,��'AR>�\>�=lū=.�M>%<c���ƽ�#H���-=i��=��^>:<?a+>�7�=3��>�����L�Sթ>��@>s�)>�2@?"�$?���9������#.���v>8j�>LL�>(�>
�I�1�=H(�>=�a>������Q��((A�ikU>k�z�X}`�eu���s=����<��=*W�=����{R:��>)=�~?���+䈿���e���lD?m+?� �=V�F<��"�E ��DH��8�?o�@m�?��	��V�%�?�@�?�
�����=�|�>�֫>�ξ��L�ñ?t�ŽHǢ�ܔ	��(#�XS�?��?��/�]ʋ�Cl�f6> _%?��Ӿ̯�>�l��6�������0t��DW=���>&�G?Y��9�t���@���?q�?q��f:��� ɿ�@v�JD�>[}�?��?kn��Κ���>�:a�>'y�?�mT?m�a>XW޾�\P�Ϥ�>%]=?m�Q?�K�>j��	(��?w�?ﺅ?��<>}��?Bo?��>2�P=52��&��������?<��� 2�>&��=*���[H��{���p����d�nV���A>�-=_
�>�?�h���[�?=�]�o�d��jZ���>�Jq>���>��>�1?F(�>vқ>�&�;gA�S銾 �M��L?aa�?Y��Xoo�Yw*=N9�=��h�	p?��0??�����^�>��^? �~?	H]?�z�>U���ו�%m��U\����<'q>���>���>����\J>�M�7h>�Vء>��>b��Ҿ6����@<0�>� ?(�>j��=�?��1?r6>-?3?$�(��`��[�'��y�>�?��>���?u�>tQ�}�\��m�����E�d�C�=��?/�)?�Ո=��a�ȥ���:�'�>"�j���?�Cj?Y�����>+R�?vY�>�_?�ma>��y�<�ھ�	�=OX�=��!?,���A��N&���_~?�O?���>�4����ս�$ּ}���{��� ?�(\?2?&??���)a�� þ2�<��"��U�R��;:RD���>~�>����䉴=�>�ذ=�Om��C6�[�f<7s�=���>� �=�/7��y��)=,?�G�eۃ���=s�r�:xD�P�>�IL>����^?�l=��{�����x��4	U�� �?���?Wk�?���8�h��$=?�?U	?g"�>�J���}޾=�ྙPw�~x�sw�d�>���>�l���L���ۙ���F��f�Ž�v��K	?���>��?��
?Ì[>x��>�o��?7�)���@۾~�j�.�� �9� |(�����^����h�*H��gc���戾�Q�>K����>M�?Orw>n�>Q��>Gb��( �>O=F>�}�>dǟ>	_>��>�Q�=A'<��ٽ��U?	����1��������<?�I?{c$?=b������fӾ��-?
��?<�?��>��k���=�%{?��>�9���?�d�=?E9;L�H=_h�����/��lg��t�>K7����4���;���y��?�E?!����9ھ��D�����->|�y?�S?�g��gp�vNV��W�F�J��K2�CdȽl��p� � �}������,�������.����=es'?�fs?U�,]��*�̾��v�Y�!���c>��>H��>���>c�>Gc�N9��sJ��P-���x��~�>)P�?Ċ�>)�I?�
<?IqP?$jL?���>�]�>�'���h�>ԍ�;��>��>ө9?��-?S:0?�u?�j+?�c>���������ؾ~?٦?�E?6?e�?�ㅾ��ýf/����g�`�y�L����=��<$�׽u���T=+T>��?[��z18�l��~7k>d7?ާ�>x��>#���԰��F@�<��>��
?@��>JA��=�r�!�����>�.�?�d���=�!*>��=�z�z�g����=�6ļ��=�oo�A:�, <���=�|�=�w��u�:�j�: ��;&��<dw�>�4?�|�>���>&ݽ����_5�x&=�ԕ>>Y>�(���$��l����F��93k��.�>V\�?���?/�d�ȹ=���=u"���	Y��ﾜ�ƾڻ>k��>��?t�,?��?xw8?]�?�>�2���y���Pھ��	?�!,?p��>��3�ʾ�𨿻�3���?)]?b;a�ܻ��9)���¾�Խ��>�Y/� /~����D�������}��$��?���?�A��6��w�M���[��ŕC?� �>�V�>��>��)���g��#��2;>���>.R?2�>��O?,�{?�s[?�KU>�8�d�2�����8���!>�@?l��?:�?[�x?��>��>|�*��z�}��� ����r���NN[=4?Y>Rґ>7Z�>8l�>N��=aǽ�௽'�>��ɧ=�,b>4<�>�,�>��>�w>���<p�G?��>
Q��ԓ�ܤ�{���=�̚u?ɖ�?%�+?��=K����E�MN��C�>Gp�?���?27*?��S����= �ּ�߶���q��&�>�չ>�*�>~��=�#G=�]>��>M��>|$�<_�s8��EM���?F?�x�=}fſ�q�(�m�U��Tw�+씾��j�Ӫ����F�N�={����n�EР��PG�3��}
���沾�Õ�|�{�<�?�"�=ȿ�=>�=0�9�ɼԈG=�Ud=�Q9=��Y=/�y��o�<\��@��s\���3�W��<�R4=�m����¾�'?�3>?b�)?��G?aB~>I�>��k��U>o���Y�?��	>|*p��	ƾ�BJ�/N��Ë��6#龃�۾h[������(>R׼�6�=�n>��>��'=~��=M=�s�=�DT<�b=���=�(�=��=�Q�=�>�H>�y?ؼ������ �\�
[�I�3?�@�>z��=���s�X?
|U>*�w�-?���>�^_�?O �?M^�?�m?�S�L�>�҉����=�0�<����LJ<�{�=�Z%�v�>
"�>
�4�@��ֽش�?#|@�5?����6ݿh�&>H�7>,�>R�R��r1�u\��]b�jUZ���!?�Z;�S̾V�>�й=�$߾�ƾ�8.=�F6>��b=Z���R\�xf�=�{�p<=@�l=��><{D>���=_���=5hI=.I�=�O> ����7��e-�r:3=1��=މb>��%>���>��?�a0?5`d?;�>�*n��Ͼ�E���0�>L�=�G�>���=�pB>zq�>L�7?T�D?��K?|�>��=��>7�>��,���m�jm��ߧ��A�<P��?y̆?j�>AR<��A�ȗ�mh>��/Ž)o?cO1?�k?��>?��	�п̺���������3CԽ|��� ��?���q~�����B�t��>>/��>H��>��>p	(>���=E��>ӑ�>�qJ>W�=��>�Kk�(��<n�9��E��%�=��������#5=��b�{ϔ�8����:��\<��>��)<R�=�>�>�r�>���=���2>�0���W����=�ǒ�"0G���d���z�6�"�,,��/[>��>(�ǽ�=��u�?�#;>L!b>��?��r?N��=H����ᾜ[����4�|�Uu�=�Q�=�"���@���U�|eG�j۾a��>iߎ>%�>��l>�,�T#?�d�w=��Zb5�g�>�|��+��)��9q� @������si�qҺ�D?�F��_��=^"~?	�I?V�?���>���Նؾ?;0>�H��J�=o�\*q�Bi����?'?���>�쾔�D�dG̾�	��8޷>�4I���O�MÕ�H�0�?��Pͷ�Q��>����X�о�"3��g������*�B�HOr��>��O?A�?�:b��W��kSO�5���/��rq?V|g?�>�K?/A?�%���x��s��^u�=�n?���?�<�?�>з�=�$��`O�>�'	?���?���?��s?>�?��T�>՞�;�� >ī�����=��>�d�=�"�=�s?��
?��
?�P��'�	�e����^�n��<�]�=�i�>9R�>��r>{��=��g=95�=�\>KϞ>��>y�d>��>�U�>�tr�%?�
>`�>ouU?8��>ض!<��a��+�=*��`}u��Xc��� ��# ����;Xօ=��D��r��>�kƿ&t�? .>�����)?�ҾCa ���->�:�>Q<�N?���=hӂ>aW�>�J�>g>��>�>�g��r>Hq�����$N���E�}4���w>!\p�=��������O��2��`����kd�"�����B���5Q�?�!�fbf�#�*�v╽�\?먔>z7?�>���
�o�>?��>�ʧ>�,��R������y�k �?���?b�S>���>`�o?Z�?�v6<�W��Mh�l1I�ƈ����"�&#c�j+��xN��t���/��Chf?xQ�?"�[?���=M�><��?� �i�V��]�>-DB�At�'>Nů>gcӾ�ɾq����Mab�D�>nhp?1?��?�̝�Q�l�I6'>��:?~�1?�Ct?��1?�{;?�W���$?��3>HC?Cz?@y5?-�.?��
?��1>�6�=�A���t%=qm��<犾5jѽ�ʽ,F�3=��{=�}���<�e=  �<U�+׼j�!;%r��݌�<��:=���=�-�=��>@�j?�?���>7M?���8Fb��,��B�?b�X��f��ξEξ�{�Ęm<�|?��?�qi?E��=�*2�22�?�=��>�>��>B�>�@S��a�=�/=S>�R>���=�;+�����Q��K����8���Zb={*�>��r>L���<
�=����FDi��>R���SwϾ�1ӽ��N��3�E���J��>�Eg?�^%?�>����3X	��m�Y?s?&T?�F�?0�=d��S3��q���q�i��>��������_���ʮ���M��j�<�-J>�Ѿ΄��xx�>N��.�����=B��z�:m�=|���]�=��Ȁ���LU��>L�o>�h��_�/���۹�@�L?[�/>��y�3�ٽ�-.�=A�?r�I>��3��\�=�/P��|��n�G>b��>&�N>n���)_��^�����>�D?��a?7��?�s���u��=�L(�;N��q�I;Q?R��>k�?g8(>t�j=E���u����^��ZD����>34�>;����F�HX��j���,���~�>�W?i�
>�r?�T?l�?c�a?��'?���>k��>�ˡ��#��#A&?~��?��=7�ԽܺT� 9��F����>|)?+�B�x��>1�?��?(�&?M�Q?��?}�>A� ��A@�1��>�S�>��W�,a��� `>�J?���>�8Y?KՃ?0�=>�5�+ࢾ�ʩ�I�=�>�2?�2#?��?	��>`��>ޭ��l�='��>c?M1�?��o?7l�=��?�=2>	��>���=V��>w��>�?|UO?��s?��J?���>؍<5�� ���"s��P��u�;�qG<�y=<���9t����u�<z;�;���M���?񼅙D�����e�;E��>�x`>����W��=Q����t�ߣY>+����H�����X�K��� >��>b�?h	�>"�?��=���>T��>)�'�5�@?���>{$?�>��f�b*���D��~>�yM?�j>�ف��W��%̄��R�=� c?4W?��X���0�b?G�Y?V���Q�W��p����f����N�?�� ?c���P1?o�?�s?���>�\���������k�6�b�e�x�"=�Ah>fԾ�Pg�̨>i�??�y�>��9>T0�=>���Q�r��롾�?fj?W��?�%t?/��=`�`�zٿG��7E���"_?���>������$?Q�(��_Ҿe���T����h�V���v��+����;��f^%�����bͽ$�=�r?�q?^�q?r_?X{�F1d�Д_�����S��|�����E���D�h�B� �i����y��\����V=Dyy�s@����?�&?�Q)�\t�>-2���~��ξ��F>Q�tu��K�=}Ћ��k?=�QS=٥c� �)�)̪�9?):�>�i�>��<?8�[�!�>�6X2���7�����&3>h�>ɬ�>�h�>ď���$��%ӽ�=ž�s�e{˽8v>�zc?��K?��n?s"��11�}����!���0�������B>h�
>W��>�>X�7��,&��E>���r�����d���	�xZ~=��2?/�>y�>X�?�?aZ	�gU���
x�j1�� �<�<�>��h?Q	�>�܆>��ϽN� ��g�>��l?�� ?J^�>�:d�*n#���w��J��E�>ۍ�>���>ց>;�6�P�k�`Z���{��)	,�\/�=b\Z?.ℾz�8�� >��S?�+8=he��x��>���[�̣��k����9>Hp?��=%��=�)ʾ���q�iS��~I)?�F?З��ԟ*�kU~>�"?j�>,�>��?��>V�þA�Q���?��^?�[J?�~A?�U�>��=�����Ƚ�'�L�,=��>��Z>S�m=\`�=�����[�G:��;E=�?�=ndмщ���G<���&�L<��<b�3>Կ��A�.^�ս��$�����s����+i�[�R]%�����}D���H��S�a�]���c��)�d=x��l���?u	�?(s��q=���Y����s�XZ����>�M��yT;����W���?��U���y#�����F���^�}�q��6%?ԅ��ƿ����?r��?��$?r?U��=	��8�N�/>u�=)�����	$����Ͽ0ۢ�X�a?׭�>g/�$H꽺��>�ڎ>]RN>�[>+����^��T��<��?�$,?�?�>�u����ɿ�غ�>I�< �?e�@#}A?I�(�{���V=l��>�	?��?>�V1��I������Q�>�<�?7��?��M=$�W�u�	��~e?��<:�F���ݻX!�=VG�=%F=����J>'S�>����VA�c:ܽ;�4>�م>>�"����4^�ɬ�<ˊ]>5�ս�6���ք?�}\��f��/�H����>��T?KG�>)��=Ь,?�H�yϿ�\�k.a?5-�?Z��?��(?H濾�ɚ>�ܾ�yM?}A6?m��>lj&�Ͽt����=�#��[������CV�jB�=���>4B>�5,�&����O��h��-*�=�) �p�ÿ��$�L��@�*<|���<��������f��K���f��*gf��� �SkI=X��=7�E>踉>��N>��]> �Z?��s?Is�>|�=ʽ�A���=F��=�<�>�}i �~����.�����`�,�׾4��|���Q�о�4<��0�=��T����O'���Y���/��23?C2�>S꿾S�=���<.�ھ�����ܱ<�l⽾/����)�	Cv��O�?��X?�����J����hT�"��=��P?]g�|�Ѿ�tľk@�=��=/Ɯ=���>[�=S���x�<��e��u0?a\?偿��`��5+*>�� �x�=��+?��?�Z<�%�>zL%?Q�*��6佫c[>:�3>�ԣ>Ӷ�>�7	>���X۽t�?ֈT?��O����ڐ>/c��2�z�t.a=0>#?5��أ[>W[�<	���U�|P��j6�<�/W?V�>�j)�i��'����!��R<=>y?4�?�؟>C�k?�PC?V��<����r�S��u��#l=ӟW?"i?��>�W���о�Y����5?�e?�lN>}Fe����^/�/O�WF?�n?�]?�꘼C&}�$$��q��,6?
>x?��]��٠�������R�>z�>^;?!-���>�N?ݺ��l����w¿�O6� ��?�>@�U�?Y|�<L�d;#���W�
?�#�>/��)G��z�	��ݙ��j�=)��>c�v����������ܽ�H?R�?_c�>�ư�J
�y��=о���Z�?F�?Hs���.e<����l�Ql�� x�<羫=�����"���f�7�"�ƾ~�
�횜�=Ͽ�ύ�>�U@`<�	=�>98��-⿂DϿm��+cо��p���?�u�>4Ƚܢ����j�Ku��G���H�2���w?�>Z�>���}�{�jo;��L��J�>�%���>Z�S�s��U����?6<�>?��>ȱ�>�N��-���Qř??��(:ο򥞿���X?2m�?j�?�r?O�;<�w�9{�!0��,G?��s?�Z?��%�Eh]��8�%�j?�_��vU`���4�tHE��U>�"3?�B�>T�-�'�|=�>���>2g>�#/�w�Ŀ�ٶ�=���Y��?��?�o���>r��?qs+?�i�8���[����*���+��<A?�2>���K�!�C0=�RҒ�ü
?V~0?{�c.�L�h?m5f��Zq�;9*�$�	�|H?̺���A��*��={����7��Y����)��[�?��??��?w����"�qN?a��>�R���A��+32=O{5>T�v>�4�>ފ뽠��=�[/��n��Xu>���?�� @�;?]���ꬿ+G�=�'s?� �>M�?�v`>�ؓ>�W>Kʐ�w�)�ܝ�>��Z>����f?�P?� ?���=;{��x8��&f�}EL��&���7��Vr>�r]?�>?�HX>��ɽ�̌�ݙ*��pڽ�4h�H�*p�	�T�"���c>�:i>>e�{���.�?Bb���ܿ�5����a���?�<�>*�>�E澄���=�$a?,j�>�-$�N���4���!��o�?���?�?K���$���ey=?$�>�H�Dg�<���,�>�Q?ۗ��A��ҋf��!�>�<�?��@uX�?qe��S?'��W`��nd��Tܾ{㱽�2>�7?1����>N�?b�>)1s��V�����o��>�@�?�Z�?r�?l�n?�����<J���g�>9��?k�>���=��پ�3=��"?8���������U�t?�-@f�@��[?~"��4ӿ�噿�u������W;S>���=�8׻�#��|�<?���+s"=�߼I��=�,h>�@>�pn>k�>'�j���>S���JD�5婿����B�*�?N��" ��_������O��������'�ƾ����\x5�k�>��A�'�{zu����=ƫU?�R?�p?܏ ?��x���>���n,=��#�ƽ�=�-�>,g2?r�L?�*?I�=	�����d�`��s@���ʇ����>�tI>�}�>�J�>u$�>�&A9*�I>�3?>���>�� >�V'=`��M=*�N>�M�>P��>z�>0p7>&�&> ��4����k���z� ��s��?�����F� ��v��G������=�/?
�=S���W�п�쯿��G?��Ԕ�&j"����=��-?��Z?Q>xԳ��V&��D>�w���]��$>y
��`k��)���?>��?0�E>HΨ>�T2��1�Ts��¾��>!%?�[�,Ž�W{���3�o9��յq>���>�&��i%�\��:��;�$G�=ؼ9?��	?�QB�d^���M���Ͼ&)�=v��>xM<-ߵ=�ci>���$���W�����A=ꞃ>�B?��+>�\�=U"�>?��,N�*{�>4@>��)>4@?��$?2E�f����ȃ�.�^?v>�9�>�6�>s�>ѦI�"��=���>�Zc>��
�R������+A�WW>��y�ѷ_�%�x�0wx=�}�����=��=d���g�:��`(="y�?<ŧ��E����羹�߽,�Y?�-?�m>yl1�>�-�	��8E�*e�?.�@&U�?�����J�g�?Iy�?Е�t?�=�;?�g�>�����Ә��??v����� ����xȤ��N�?�T�?WH�=�׉��g��� >�%%?���cR�>L;�Aڝ�1g��`��T+ս	��>D .?4P���_�==y:��W?V?���Y�����̿Ƃ���>7e�?�
�?
g�5���S�,�ɺ??I�?G�7?�&�>����r����>	�1?5?��>�"�XQ�g�,?/��?���?�uK>ۄ�?�6y?�m?\�ļ$3��Ѭ�l���_^�<�=���>���=����0R���;��G^�x�x�U>��0=�¬>9&潚֣���=�z�+Zc���ڽ���>��l>��g>��>E�?��>~��>2��R���
kl��:����K?�?��	�ARp����<��=�T[���	?	�5?�o����þ#$�>7]?��}?{Y?�>���(��x���y���P0�<\!S>��>@��>@|���jC>B�پJQD�)��>�3�>�o�vؾ�Ӂ�]��;^��>�u?��>*J�=��#?�T(?�r�>��?���!������W�>G??Y/?	�?�?�C��;]�u���-̟��hT�Ƞ�>aW?��?�0�>�M���Ŀ+�ý.Z>��A�?�GW?�ɾ=�?�n�?܎-?�pM?���>ͻ}����Ʌ����>��!?��
�A��L&� ��Yv?I??���>oO���Hֽ|ؼ4��Cx����?�/\?�M&?����$a���¾�W�<{�$�	T��< <A�D�!�>��>�������=}>��=�Om��R6��f<�'�=|�>��=7:7�|��0�+?�C��Jw�;#�='6p�Q�C�@�r>�O>�����\?#D���{�r������d~U�,��?���?L��?����Vh�2>?ߘ�?�?ɏ�>K��}ܾ�߾u�{�xea�@��>�N�>d뼙y�8���(N��z��H������
?�k�>��	?�F?��@>I��>̃����N���ľ��ľ,�p�����6�6<�T�����F,�^��ľz�����>a[μ���>N?�S�>;G>>�>��;1y�>>HG>|�j>�t�>�W�<� >��=�,���g�V?Y��T��/ �Υ���7E?b�f?)�>�%�������PJ?���?�'�?�h�>p�V�M��>��>���8�&?E<
>�޿����=����A���\��=���>�刽�b2��'g�h%��bo?�u?]w�=�پ<c��g��QRp=FQ�?;5)?�)���Q�ؗo���W��S�_��$�g��}��S�$���p���nV������(��N*=�*?��?ώ����G���#k���>��^f>�K�>X�>���>��I>��	�Q�1�:�]�.W'�˱���W�>#B{?s��>	vI?�<?6<P?�^L?���>ְ�>]��a�>'6�;B�>��>�r9?��-?�e0?�?\u+?�c>�g��`���q�ؾ��?�?�(?�?�?\䅾X����O���d�b�y�2.���~�=�S�<x׽�?t��;S=��S>oX?�����8�g���H
k>Ѐ7?e~�>	��>6���.��5�<�
�>e�
?E�>8 ��}r�d��S�>j��?���r=��)>��=�����κM]�=������=�1��Ć;�ts<��=-��=�Wu��}��D�:��;�6�<�6�>�+?��>��	?�E�R��R[�A&�=��#>�2z>1	=/F��Ǐ�����[�X���|>�k�?P3�?�=`=�W�<5�^>&s��r�0���Ⱦ�<˾�X�=���>�0?f-h?3�?8�&?��-?	��6J��h��0S��������	?�L ?�k�>@����¾�[��K38��-?�W�>�aG�g��*�/�<���.�T��+>$�; x�~����]�-"�����`��1��?ϙ�?�צ���6��1׾T���޾e�A?O8�>���>���>��)�>Gr�#��=�>w��>ŉd?�"�> �O?^G{?�[?�T>�8�%���̙��]<�L�!>��??���?�؎?c�x?"m�>R}>�O)�x�߾�5���_���߂��W=Z>�\�>�A�>���>T��=�ZȽ�̯��d>��p�=�b>�a�>�v�>��>�1w>�p�< �G?^C�>Vp����ME�������I��t?�W�?ܩ*?�=���2F����"�>��?�?;�)?��T�s�=���O��Q�m��>,��>M~�>���=^�J=o>f��>�@�>��)�d�8�7�S�P?P�E?<��=i�ſV�q�F�r�z����!I<#p��@�f�ϗ���W��f�=�ʗ�3��Щ�t[��^���꒾P)������Gy����>|(�=�!�=���=�~�<28ؼ���<�oS=�N�<\�=��v���B<	oD�t���������k[<p�G=J#�E:˾��}?��H?�o+?��C?D�y>�>��5�<L�>򘂽�<?[ET>�Q�7����<�hǨ�cC����ؾ�H׾�d�������	>N�H�\F>�X4>��=`��<��=��t=�:�= �.�v�=#	�=l�=T�=���=!->!�>�=}?ѐ���P���G����dh?�q�>&Ta>r���B?���>,�x�&J���j���f?��?�s�?�S?=$s�%��>:������;��H=�ж�� M>���=����x�>~s�=Ah�p�	�=���?�=@A0$?����`xݿ�5�=g�7>�F>��R�t�1��i\���b�}�Z���!?�S;�M̾.2�>���=�*߾��ƾce.=?�6>?Nb=�d��M\�b��=��z���;=�#l=?Չ>%	D>�v�=�.����=ԏI=���=�O>6#��r�7�4�,�$�3=N��=��b>W�%> ��>�??�C1?Fyb?b��>�m�d�ҾSþ<P�>��=K^�>d}=�	=>�(�>�8?��F?_�K?��>�ׄ=cq�>�ע>s�*�Dj��!�'t��4
�<��?�?�J�>Ur<��C���u%=���ս-?��0?6\?��>.��2Ͽ���=��Q�|<�rB�0�\���\���/=���]�Jx�4� >�eZ>]�>���>���>J��<�Y>'�>�T�=$%0����=m�����<WA�=940=�Y=P�=������K=j=����;�eu������6=���=I� =���=R��>�M>�Q�> Z�=�G��8�>�g���1R���=�=����E��`a���|���*���7�6�=>XPT>��Y�+���l?��B>f�S>{�?`�o?�>y��F׾�����=��n����=-��=k
k��':�eg^���J���Ѿ���>}�>��>��l>�	,��"?�װw={��a5�
�>�z��7���-�K<q�K?��0����i��RѺ�D?�E��Ҭ�= ~?ֱI?��?��>� ����ؾ�20>{=��f!=��]q�ao��B�?'?���> ���D���˾����{!�>��G�EP��ᕿ��/�[�#������>����x�Ͼ��2��j���<��6�B���s�b#�>`P?�ۮ?c�?p��yO���?���_�?J�g?D��>�2?��?�`���������ȶ=��n?���?�l�?�
>r��=ܵ��y�>`?7��?�ԑ?P�r?d�A�\��>�8�;��>1ږ�C�=v,>���=�C�=�R?~
?x�
?-���q	���a�J a����<�^�==^�>��>(Yq>�5�=��^=�=�Z>#�>ў�>�f>�L�>R��>]gd��Hʾ>%?��<sT�>hR?T�d>�.������S��=�$r��N��KO�iڻ�i�ɸ,��r��3Y��k���>f��|p�?E>m���A?=n��
T�G4�>b�i>�ތ����>&"�=	��>G��>���>HY�>1��>f�Y>����A�>�������ۄ�Bh�geJ�S�R=1����e�==��u-<T0;��㫾��Yp�����lj���R=�#�?��-��k����X�y=s��>�c�=�?W��Ɉ�;� n>t8�>-]>���ۡ��썿�k�1Ԕ?�I@�>���>��n?��>fܽ/	ֽ��l���k�b|O�ԂF��~��!����y�ɷ��9�=�b?:�q?uG?�3��/>B�Z?vm	��ٽ��/>��E�J�?��E�=�RB>Ȝ��\���XNվ:���wൽs�~>���?��g?>�>iG��-�m��'>��:?Û1?�Ot?��1?\�;?�����$?8o3>}F?�q?2N5?��.?,�
?g2>
�=j����'=�6���M�ѽm~ʽ��q�3=�^{=%θ�<R�=��<���ټݪ;�%��H%�<!:=U�=�=U^�>��.?r*?���>k0?�G:��x`�9";���>�b�������\�x~����>Uj�?x�?��2?��=tm
� �}�S�>û�>�@�=��4>L�>ɞi��k=�5->��2>Ze�=����Ř��ʿ�����m���;r$>�I�>���>I���g��=@;+�-]x��2L>�l��@N��J$���5��A+��h�l�>O�L?ou?"V�=L.Ծx��;��r�7MB?��
? �M?	�?4t=���������I�ܚ���>*]b�r��ޒ��`����k6�B���
\>�N�������_>������M���9����d
��g���Q4>����9m�ñʾ�j�>tJ
>Ε���x�삗�J����c?���=^.ھD^�K���$Q>��>=�>^��W��[�D����I�S=˖?Bf`>�_��"��G�����ӆ><F?6�^?�;�?�_���=t���A�D���ޢ�:��m�?T�>��?�:>�=�����h�r,e�E���>���>P����D��3��c����"��3�>�Q?<�(>.?�P?K?@"^?#Z)?��?4Ï>�f��yR��B&?)��?D�=��Խ��T�Z 9�AF�A �>v�)?E�B���>q�?��?�&?��Q?��?u�>�� ��C@����>iY�>��W��b����_>��J?͚�>_=Y?�ԃ?��=>I�5��颾�թ��V�=@>��2?�5#?E�?���>7��>A���i�=*��>X�b?k;�?.�o?a��=z�?�2>;�>~�=�n�>�l�>�?IO?��s?��J?j\�>^:�<��,O��@�r���P��x;�A<;fx=C��z�s�!I���<�u�;~巼n����－]D�i?��=7�;Ϫ�>k$t>WS��4W/>�?ľ�ڈ���?> �������5���8��u�=���>�	?�'�>��#�p��=uļ>q2�>���(?7'?�?Vc<;��b�s�ھ��M�hʰ>�aB?Dd�=��l��T����u�k= n?e^?�Y������g?�K?x���G��՝���+�Z����v�?��?�s�����>���?q�l?u�	?��G�+ք��E���$�����U�=<ji> �Ͼ��u��6�>I�J?���>�>����̾�j�Xd��[?���?���?�ۇ?h�=��.��Tؿ�+���Y�b?���>o꠾FA-?6%<5bھ�霾�<v�Jݾ噣�����>͕��s������jn��?���"�=a�?Mo?�lr?[	[?����Pd���c��L~��X�u������-C�;E��@��h���>i�/�~���=�r�ɹ>�{��?=�$?G�)��0?���N����ؾs�X>�盾�a
���_=䘽=��X=�9T�h���2���l?SU�>��>XA9?K�W���=�	6��9�( �G�9>��>�;�>�'�>�3���S-�;ܻ�������\�"���/m>��h?KJ?n�w?���b7��U|�r�$�|��Hž��a>y�=���>:z�^4<��s&���>�u�/=�	q��	~�x"�<�;?�_L>��e>��?= ?�����@QL�w�2�PQ=�.�>�b?5I�>r�d>�Oͽ��
�!`�>٪v?i��>p��>Y4�U$��x�g�:���>$�A>v��>��>b� ��^�����N"���~(�֠l=�tH?4t�OD�`�N>�R?/�=-\x����>Ldؽy�3������^<��>u�?4^�=��/>�ԾC�.��.}���T�_T)?�H?�˒�,�*��>~> "?�c�>�r�>,�?��>�Kþ���?��^?�@J?:A?d�>��=ȋ��XKȽF�&�U%-=���> �Z>)*m=}��=N��O~\��1���D=O�=��ͼ�X���/<������J<<��<�3>��ҿ��B�%�־�"��������~l��y������]���7���p�u�o�B���}����!�6LN�m~��N��_X�?R��?������Z���! d��fp�̺>k��N=�<\'��R�W��߾뒹��������z9�(Qh��Fg��{)?Tר��Hǿ������3?��D?V�k?�z��A4�S'E�Z��>T��=�<S>3������Xd¿aC��W$h?-��>����K���j>��>�K�>�{Ѽ��>�X��n�ֽҎ?j��>	�?�����%̿9���M?=,�?�@�|A?��(�(��nV=��>��	?X�?>�T1��I������S�>�;�?��?�|M=��W�|�	�e?د<��F��ݻ��=�E�=�F=^���J>�Q�>���WA��8ܽ�4>dم><�"����O�^�-��<��]>�ս"5�����?Go[��*I���<�p�����=�wW?�؟>��&>��J?BV�;{ǿ�zV�^�h?џ@���?��)?��TG�>�澙�T?SQ;?6��>���]��V�=t]	��U�����ºf��C�=Gi�>OmN>��սɋ��R��������>�8���Ŀ��"�F�;�y<��)���y�j����x��ݦB����q�h��ҽ�Ռ=���=<U>�o�>�Y>UmQ>�Y?z
m?\��>F�>��=��Y��q]��ig�F,�����>e
�����i龆�߾	�7�~��� ˾��<��\�=�Q��'��h�'�1`�2�<�ݶ'?y@>�ֿ���K��c�<Ѿ�\����������$Ǿ�0��n�cL�?�D?�Æ�+�O�=�b�Ӽ��μT?B������{��~�>�q���o=QP�>���=>��:$6��V�J�0?I?ـ���/���	+>� �2"=�,?�g?0
;<���>Ώ%?=w(�h��	]>��1>���>G��>��>d/��6(ڽS�?%dT?;� ����]��>CԿ�Oaz���n=�>?16�����IY>�֜<t���>IK�H���7�<�(W?X��>Y�)����b��}���^==Z�x?v�?d*�>�zk?��B?�ݤ<�d����S�� ��Gw=��W?�(i?��>����оȄ����5?��e?��N>rZh������.�?U��$?(�n?�_?rx���u}�������m6?�yx?59a��b��P4
�^���T�>��>,�>}x%��E�>#RA?��Ž\J��'���ϼ0��ϝ?;� @.��?0	<=T����=�k?Tκ>ӡ��1r�gqx����x�=�?t���ۿ����G�Z��<�^?-�?��?�������"��=�֕�y[�?;�?�}����i<���nl�b~���4�<л�=��"�D���7���ƾݵ
�o����A�����>�X@�I轾+�> ;8�'6��UϿ����eоTq�<�?�h�>��Ƚq���|�j��Du��G�"�H�����n�>�>Rڞ��Q��+�}���:��j'�U)�>i���נ�>�V�X
���Ģ�X�<�4�>���>��>\"��?����P�?Y(��U�Ϳc��W��u�W?�?1��?|?�K{<��{�~�q�wE����G?�r?�W?�/���d�?Z�H�j?9l��\`�(�4��;E�#JU><"3?�<�>_�-��|=�4>M��>�h>�&/�F�Ŀ�Ѷ������ �?���?�f�7��>���?.k+?�f��5���Q����*�dr �>A? 2>������!�n4=�5����
?׎0?0}�V9���_?��a�~�p�B�-�� ǽQ١>��0�a\������z�0We�5���Ry�{�?p_�?o�?n���#�a5%?��>?����&Ǿ�C�<�l�>��>�,N>f__�7�u>s���:� V	>v��?O~�?Pn?����6���U=>u�}?`��>�wr?aԯ>-�>WST>�:���﫽^��>h�>#M;<�C?�S?��?��=An=6 ��a�ޙF���3�s�;��%_>Μz?SiK?�/>)AJ��n=}fJ��u��Q8�=E޽I�p��ݺ=�xQ�')>Țv>��>YU��������,?z]7�`8߿Kۍ�[��hiX?	��> 2�>l��_g�*O�<�8f?|��>����������(Q*�6~�?C�?� ?Nƾ5 i����=���>騋>]��.��d��V�>��V?E�$��Æ�����u�>ɛ�?m!@	��?Z�/K?��
��W���{�H�ﾪ�ҽ�
>}�0?��>���>H��=�k��z���v����>P`�? �?gF�>�Ad?ղa�ۼ0��^�<���>>r[?��?D�~����/_>hc?WB�đ��8�	�-Os?�r@�@�S?�L��)l˿�Ĕ����zо�ʈ=��={�>��Խ���=�f>�=��v=�d>ڤ�>z�J> ��>�Z(>諊=ê>�x����#[��wv��wA�k'��d��`7��%���+��%����P�ؾ�|����`B�+���b����<=>�M?��i?�lZ?I��>giֽ<>n�Ҿ�
=r沽��=��>;RQ?��=?��3?�1=/Ѷ��Te��݆�f���t'�����>�f>ֽ>@˯>���>
`� >�4>0�Q>O��=�4�=6��;K��<��4>?��>���>�>/>B>gm>�
��ے���H|��`�jY=�?}3N�pT/�l����)�lľ�@U>��)?� �=�����ο+�����M?M�����j�7��&4>�7?�iI?�IC>�T��{���x�=}����[����=n]��T��w<.�	�Y>�{+?T�f>pu>c�3�X8���P��s��x�|>�*6?�ö�v9���u�z�H��lݾE�M>=ƾ>ID��l����l�7i��+{=�h:?m|?�벽���� �u��,��'AR>�\>�=lū=.�M>%<c���ƽ�#H���-=i��=��^>:<?a+>�7�=3��>�����L�Sթ>��@>s�)>�2@?"�$?���9������#.���v>8j�>LL�>(�>
�I�1�=H(�>=�a>������Q��((A�ikU>k�z�X}`�eu���s=����<��=*W�=����{R:��>)=�~?���+䈿���e���lD?m+?� �=V�F<��"�E ��DH��8�?o�@m�?��	��V�%�?�@�?�
�����=�|�>�֫>�ξ��L�ñ?t�ŽHǢ�ܔ	��(#�XS�?��?��/�]ʋ�Cl�f6> _%?��Ӿ̯�>�l��6�������0t��DW=���>&�G?Y��9�t���@���?q�?q��f:��� ɿ�@v�JD�>[}�?��?kn��Κ���>�:a�>'y�?�mT?m�a>XW޾�\P�Ϥ�>%]=?m�Q?�K�>j��	(��?w�?ﺅ?��<>}��?Bo?��>2�P=52��&��������?<��� 2�>&��=*���[H��{���p����d�nV���A>�-=_
�>�?�h���[�?=�]�o�d��jZ���>�Jq>���>��>�1?F(�>vқ>�&�;gA�S銾 �M��L?aa�?Y��Xoo�Yw*=N9�=��h�	p?��0??�����^�>��^? �~?	H]?�z�>U���ו�%m��U\����<'q>���>���>����\J>�M�7h>�Vء>��>b��Ҿ6����@<0�>� ?(�>j��=�?��1?r6>-?3?$�(��`��[�'��y�>�?��>���?u�>tQ�}�\��m�����E�d�C�=��?/�)?�Ո=��a�ȥ���:�'�>"�j���?�Cj?Y�����>+R�?vY�>�_?�ma>��y�<�ھ�	�=OX�=��!?,���A��N&���_~?�O?���>�4����ս�$ּ}���{��� ?�(\?2?&??���)a�� þ2�<��"��U�R��;:RD���>~�>����䉴=�>�ذ=�Om��C6�[�f<7s�=���>� �=�/7��y��)=,?�G�eۃ���=s�r�:xD�P�>�IL>����^?�l=��{�����x��4	U�� �?���?Wk�?���8�h��$=?�?U	?g"�>�J���}޾=�ྙPw�~x�sw�d�>���>�l���L���ۙ���F��f�Ž�v��K	?���>��?��
?Ì[>x��>�o��?7�)���@۾~�j�.�� �9� |(�����^����h�*H��gc���戾�Q�>K����>M�?Orw>n�>Q��>Gb��( �>O=F>�}�>dǟ>	_>��>�Q�=A'<��ٽ��U?	����1��������<?�I?{c$?=b������fӾ��-?
��?<�?��>��k���=�%{?��>�9���?�d�=?E9;L�H=_h�����/��lg��t�>K7����4���;���y��?�E?!����9ھ��D�����->|�y?�S?�g��gp�vNV��W�F�J��K2�CdȽl��p� � �}������,�������.����=es'?�fs?U�,]��*�̾��v�Y�!���c>��>H��>���>c�>Gc�N9��sJ��P-���x��~�>)P�?Ċ�>)�I?�
<?IqP?$jL?���>�]�>�'���h�>ԍ�;��>��>ө9?��-?S:0?�u?�j+?�c>���������ؾ~?٦?�E?6?e�?�ㅾ��ýf/����g�`�y�L����=��<$�׽u���T=+T>��?[��z18�l��~7k>d7?ާ�>x��>#���԰��F@�<��>��
?@��>JA��=�r�!�����>�.�?�d���=�!*>��=�z�z�g����=�6ļ��=�oo�A:�, <���=�|�=�w��u�:�j�: ��;&��<dw�>�4?�|�>���>&ݽ����_5�x&=�ԕ>>Y>�(���$��l����F��93k��.�>V\�?���?/�d�ȹ=���=u"���	Y��ﾜ�ƾڻ>k��>��?t�,?��?xw8?]�?�>�2���y���Pھ��	?�!,?p��>��3�ʾ�𨿻�3���?)]?b;a�ܻ��9)���¾�Խ��>�Y/� /~����D�������}��$��?���?�A��6��w�M���[��ŕC?� �>�V�>��>��)���g��#��2;>���>.R?2�>��O?,�{?�s[?�KU>�8�d�2�����8���!>�@?l��?:�?[�x?��>��>|�*��z�}��� ����r���NN[=4?Y>Rґ>7Z�>8l�>N��=aǽ�௽'�>��ɧ=�,b>4<�>�,�>��>�w>���<p�G?��>
Q��ԓ�ܤ�{���=�̚u?ɖ�?%�+?��=K����E�MN��C�>Gp�?���?27*?��S����= �ּ�߶���q��&�>�չ>�*�>~��=�#G=�]>��>M��>|$�<_�s8��EM���?F?�x�=}fſ�q�(�m�U��Tw�+씾��j�Ӫ����F�N�={����n�EР��PG�3��}
���沾�Õ�|�{�<�?�"�=ȿ�=>�=0�9�ɼԈG=�Ud=�Q9=��Y=/�y��o�<\��@��s\���3�W��<�R4=�m����¾�'?�3>?b�)?��G?aB~>I�>��k��U>o���Y�?��	>|*p��	ƾ�BJ�/N��Ë��6#龃�۾h[������(>R׼�6�=�n>��>��'=~��=M=�s�=�DT<�b=���=�(�=��=�Q�=�>�H>�y?ؼ������ �\�
[�I�3?�@�>z��=���s�X?
|U>*�w�-?���>�^_�?O �?M^�?�m?�S�L�>�҉����=�0�<����LJ<�{�=�Z%�v�>
"�>
�4�@��ֽش�?#|@�5?����6ݿh�&>H�7>,�>R�R��r1�u\��]b�jUZ���!?�Z;�S̾V�>�й=�$߾�ƾ�8.=�F6>��b=Z���R\�xf�=�{�p<=@�l=��><{D>���=_���=5hI=.I�=�O> ����7��e-�r:3=1��=މb>��%>���>��?�a0?5`d?;�>�*n��Ͼ�E���0�>L�=�G�>���=�pB>zq�>L�7?T�D?��K?|�>��=��>7�>��,���m�jm��ߧ��A�<P��?y̆?j�>AR<��A�ȗ�mh>��/Ž)o?cO1?�k?��>?��	�п̺���������3CԽ|��� ��?���q~�����B�t��>>/��>H��>��>p	(>���=E��>ӑ�>�qJ>W�=��>�Kk�(��<n�9��E��%�=��������#5=��b�{ϔ�8����:��\<��>��)<R�=�>�>�r�>���=���2>�0���W����=�ǒ�"0G���d���z�6�"�,,��/[>��>(�ǽ�=��u�?�#;>L!b>��?��r?N��=H����ᾜ[����4�|�Uu�=�Q�=�"���@���U�|eG�j۾a��>iߎ>%�>��l>�,�T#?�d�w=��Zb5�g�>�|��+��)��9q� @������si�qҺ�D?�F��_��=^"~?	�I?V�?���>���Նؾ?;0>�H��J�=o�\*q�Bi����?'?���>�쾔�D�dG̾�	��8޷>�4I���O�MÕ�H�0�?��Pͷ�Q��>����X�о�"3��g������*�B�HOr��>��O?A�?�:b��W��kSO�5���/��rq?V|g?�>�K?/A?�%���x��s��^u�=�n?���?�<�?�>з�=�$��`O�>�'	?���?���?��s?>�?��T�>՞�;�� >ī�����=��>�d�=�"�=�s?��
?��
?�P��'�	�e����^�n��<�]�=�i�>9R�>��r>{��=��g=95�=�\>KϞ>��>y�d>��>�U�>�tr�%?�
>`�>ouU?8��>ض!<��a��+�=*��`}u��Xc��� ��# ����;Xօ=��D��r��>�kƿ&t�? .>�����)?�ҾCa ���->�:�>Q<�N?���=hӂ>aW�>�J�>g>��>�>�g��r>Hq�����$N���E�}4���w>!\p�=��������O��2��`����kd�"�����B���5Q�?�!�fbf�#�*�v╽�\?먔>z7?�>���
�o�>?��>�ʧ>�,��R������y�k �?���?b�S>���>`�o?Z�?�v6<�W��Mh�l1I�ƈ����"�&#c�j+��xN��t���/��Chf?xQ�?"�[?���=M�><��?� �i�V��]�>-DB�At�'>Nů>gcӾ�ɾq����Mab�D�>nhp?1?��?�̝�Q�l�I6'>��:?~�1?�Ct?��1?�{;?�W���$?��3>HC?Cz?@y5?-�.?��
?��1>�6�=�A���t%=qm��<犾5jѽ�ʽ,F�3=��{=�}���<�e=  �<U�+׼j�!;%r��݌�<��:=���=�-�=��>@�j?�?���>7M?���8Fb��,��B�?b�X��f��ξEξ�{�Ęm<�|?��?�qi?E��=�*2�22�?�=��>�>��>B�>�@S��a�=�/=S>�R>���=�;+�����Q��K����8���Zb={*�>��r>L���<
�=����FDi��>R���SwϾ�1ӽ��N��3�E���J��>�Eg?�^%?�>����3X	��m�Y?s?&T?�F�?0�=d��S3��q���q�i��>��������_���ʮ���M��j�<�-J>�Ѿ���fb>���-Y޾�n���I�����J=�����R=�K�վ􍀾h�=�	>�t���� �7������ӐJ?�o=��*NV�e@��H>6�>��>�p8���y��@�a���Ɩ=+�>c�:>�����mﾷfG�����Ԇ>y+G?�^?L��?�����Ms�k�@�r���/���/���3?���>P^ ?��>lpg=�쵾g�
���f��G�-��>���>\��UuE�����(�������>�?E2>K?P\T?��?�Kb?��#?��>��>�󊽠����?&?��?	�=��ԽX�T�N 9�� F� ��>�u)?��B����>@?��?��&?2�Q?�?�>� ��?@�Ꮥ>X�>W�W�`���`>��J?̏�>Y:Y?<у?z�=>m�5��ݢ�����)�=�>��2?�0#?�?Ѭ�>���>�a���?�<�`�>=a?ʥ�?RAq?)e�=	��>�/6>±�>μd=�|�>8��>+?�hM?MHr?�I?	�>�<�Y��?e��s����w;��Y<y��<ko�="R��e�$�
A�<�<�$�����-�����r2��M����>�le>Ѓ��-�>uv޾)�=�s��>��(��ƾ�v����L>
�>�z$?���>P��S>�Ɗ>��>S�*�uT?��>"�?�sC>�2W�X���-�k�W>(�2?-N*>Ԁ������}��ku=U�_?�\?�O۽	$þm�e??�S?{�ӾO�E��iU��(��r�Ծ	,s?!?����;��>5��??�c?��?>����{��]��Ʒ:�7"�bG=\�>շ���tY�Uu�>`7?�g�>l�U>�V�=%�����z�bt�
'�>zт?�x�?=�}?v!>��Z�R�ݿ����'��]?^?�6�>�Ҧ��L#?±��]hо���N���Y��;H�����č���#��O�#���r)ӽ;_�=R�?0�r?uxq?�_?����c�L�^�����WV����3��0F��D��XC�.�m��w��v���]���4J=��}��F@�cV�?��(?+(/��q�>E���
��̾"FB>�ȟ��"����=^����8=�X=�f��!0����?��>��>�<?�[��R>���0�%+8�~����4>aܢ>�ԓ>|�>���:��/�8��Eɾ�4���ҽEu>�Qd?zPK?Rqp? �Ȧ1��g��c%!�'J2�����?>"�>�>cc�۩ �s�%�G3=���s�0��p��<�	�ʃ=�?2?�d>N~�>�f�?Z?�G
� ��^(t���.��=y<i�>@`e?ĭ�>="�>p�ӽ�' ��>�.o?e��>�>S�����"�f�{�^�ǽ��>�X�>T��>VoT>��.��ga�]����Ќ���5�?��=�Kb?�8���d��}�>�P?��^�+����_�>J���tT$��)例��S�>�|?��=�>f�Ͼ�A���z������C)?�]?-���*��U~>�"?4��>E��>u�?G&�>?rþ��?d�^?v@J?�MA?cU�>rm=�4��"{ȽR�&���-=�g�>++[>'�m=c��=����u\��_��E=�M�=�7μ����� <�s����D<(d�<��3>x<ֿ��E�i߾Z�����̃�w�������>���8I��٣��X������a��@>��K��)��g,c����?EK�?����☾e����p��絾 ��>�������Ⱦ�"ܼԠ� ��EK��)��e8M���d��`�=�"?W���ǿ����y%��3?��C?_`n?f|���-��YD���>�2&� �J=3�����vϿ2Ĵ�*�j?T�?� �̽"��>/�D>EG^>��k>��=���˾|�=B�?�A?�?2�~�&^��N��0�c=�?J@(}A?o�(�k����U=0��>x�	?i�?>�O1�$I�x���O�>�<�?N��?j�M=�W���	�	{e?wX<-�F�o�޻�*�=pP�=�N=���J>pP�>��8UA��*ܽ��4>�م>�"������^�B��<��]>��ս�O��߄?v�\�g3f�(�/�6��a�>��T?(��>2��=�,?D�G�	XϿ�.\�7Za?��?o��?��(?*t�����>N�ܾ�M?�q6?���>d�&�~�t���=��⼨���@侂�V�ߔ�=�Y�>�S >O&*����R�N��
%�=r)���ĿU$�1��6�<?Uy��V|�	���e0��IYQ�GL���*{�h	�b�F=��=�P>Ƙ�>��P>�6V>�X?`j?�U�>�&>������p����F� 	g�{� �����?��zϪ�8��ha޾���~1�EI�ȮǾ�:���=өT�{Չ���(�&~P�]�,���?�N�>��о��J���<)_��ֳ��(o�����u¾W5�a�b���?�UJ?A"����\�B#�+Y����=��V?l�������о�J�>�Ӽd��=�̘>�ln<�9��Gp3��IF���0?X3? ��mȔ�h+4>���	=�/?��?)[;H��>٦'?��(��ս%�S>'>[ٙ>���>�t>�&����ڽ`�?ñS?,@�R�����>�о��Ez��}m=�� >'~9�K�ּf�U>v�<&�4�����7G<7�_?���>�`�����z.�@�4�S =��?f�?���>�H�?��N?G�>����i�0r"�#�$�W�U?�}?���=��Wξ�,ﾀg[?��y?���>����c����]���
�50?��N?��$?{#=�vm�A����w���?�[y?��`�X֣�G�
��~E�66 ?�g�>0�>�4 ���>w|K?:�½_������Oa9���?
�@Z��?�#O:��x`�<pE�>�#�>���ܼ�)��b����C�=��
?5L���C}�,a*��+���G?�*�?��>.ꤾ"�����=2Ǖ�gX�?��?����f<���l��d��Sȟ<���=ʥ��u"������7���ƾ�
�B����B��˞�>�W@�@�y0�>J8�76⿫LϿ����ZоW7q���?�>��Ƚ-���u�j��Wu���G�.�H�f���;q�>J�>s����?���R|���8�Y,����>���G&�>��X���E
��L�u<��>���>�`�>�Ný$u����?���(�ͿD���f#�!dW?켡?g'�?�?�?`;.���$�^�l��μG?y?q?D�T?��_�ڂb�X�3�&�j?=^��bT`�Q�4��FE��U>2"3?F�>,�-���|=�>��>g>�"/�/�Ŀ�ٶ�����3��?��?�o�L��>n��?+s+?�i��7���[��n�*�eb,�V<A?�2>U�����!��/=��В�ռ
?�}0?�|�/�Hj?��h��y�b�,�� �^��>*�O� �F�R��<=m��[Q�
,�����M�?!
�?��?~����<3�r�?y͖>�ܟ��dV���d=�M>]>(>'w�>�T��.|<֑"�(�`�k�2>���?a� @�#?�Q�����2c�=~��?���>�c?�]�>)��>B}C>������@���?JJJ>Щ��B�?�SU?���>��<��W�Jo@�uu}�rjV��%L���@�v��>R�E?�b}?W��S�<K:�<)�D�n��y���_?�����Kn��������>|�)>�`�>�E�����bJ*?�V���ֿ�������^�Y?s��>���>�nƾKy���c>>�i?�.�>����Ӱ�9��.�9=�?�?y3?�v�����=�L?�1?4��"Tнu/�2$W>p�o?��:��l��i����s>Lc�?:k@?��?�2����
?�+�]J���d~����0��*>�=w6?��k>m� ?���=n�p�?o��Ԝt�xڰ>x��?�Y�?s6�>l�j?�Go��d@�+=!=�6�>#|o?��?�;⻻��k�J>l	?������=P��De?�@�9@��^?=	���n׿o���m��6)���3>)�=7.>��
��L=/��=-6�;{�E<tW�=�p�>suL>4V�>�vf>*�4=�O>z�}k�U��䒐���6�R�E���i����v+���_����������ʽ>`�;��0������=<5-�=�^V?yS?�Sq?ˊ ?��n��^>@���}9=�	'��R�=���>~�0?Q�J?��)?W)�=Jߞ���d�����§�b�����>� H>z��>��>�&�>rK��M>�0>>�Ձ>�Y�=e =?'�:�J=��Q>%L�>��>���>�7>�
>wд��ݯ���m��i��΀��s�?1?���4K�v��8x�/[žve�=(?+�=�����Ͽ����T}N?�(�����9�9���=��.?��_?Vs3>�r�� 녽�">�Ľ�U���
>�r���ʅ�^z.�ӷG>�?*�f>�iu>s�3��U8�ʩP�W��2�|>@6?� ���9���u�a�H�.Fݾ -M>G��>��B��Z�^����~��^i���y=k�:?�r?m���������u�C2���bR>�]\>�="ƫ=okM>c��\ǽ
7H��m-=���=�P^>��?g�1>��x=�,�>T◾m�L��	�>��=>1�!>C�??�#? � ��^��ɂ�`*���w>ѫ�>��>)�	>��J�0G�=���>��^>��鼄�z��o
��<���U>��w�%�]�ԑs�zK{=~���N�=��=���V�B�4�=T��?�����߂�%g�󝈾{D?��0?`=�dj�A��R���h����?�`@
d�?�A���E��u�>��?� �#3>��?��>�n��c`�j�?$bp�%־� ߾i�u���?�#�?��:�酿e�a��5>m(?�=�����>pQ�ͥ��h͂�.��)�m=���>�[E?Z]߾i���P���?0�>ţվ�'���ʿ��w���>���?��?��o�뱓�=�0�{&�>���?7?L�^>��)����>e�.?�J[?DF�>�R�77/�4R+?�S�?�,�?��D>�~�?�q?m��>e�`���2�]����势G�8=M�L;?��>c �=*<���FP�\ܓ��t��b�d�&���H>@�S=��>�ǽ�ݴ�M��=������G��>�s�>$�W>��>���>�Z�>�σ>�:�/���z�>a��p�K?�?��A1n�z��<C��=&�^�W,?"I4?�[�9�Ͼkܨ>!�\?���?O�Z?�Z�>����<���翿������<g�K>E?�>N<�>�;���GK>�ԾV<D���>̗>�y��:9ھ�2��Z롻�G�>�f!?��>4��=q�-?:(?VW�>4�>��O�錄�?���?v�?#2?-��?6S�>}7��I�*�ꕙ�������2��Xf>�0a?O�-?�C�=c����ճ���n=����[׻��?!�q?�q��9?=1�?mr[?�c?��>�$��= �"c�="S�>�0!?����B���%��d!?]?�R�>gG��l�ս����1�����a�?R?\?<P&?��ɢ_�{���(��<�
'���9b��;��
�T�>�>&؀����=E�>�5�=b�k���5�Hv<�=*v�>���=��<�閽� ,?�1�����=ƃr�jJD��	~>dPL>����,^?Ի=��|�K���񊜿�?T�3��?W��?p<�?�鵽��h�u)=?[�?�B?y��>�対�ݾŕ��Ov�cw�q#��Q>;��>
�y�[�趤�S����A��5�ƽ�g��;?�V�>q�?�r?٨9>���>EѨ��15�q;:� �_\�u*��D:���#�>������V�1�ռ��
䝾i��>������>Dh?Q��>�NV>'g�>��f=3U�>敏>�Lp>�]�>n��=��=�ޚ=xm�������U?i;ǾLE�*���wؾ5^=?��m?���>�U��1r��d�,;?K$�?+ģ?�W�>�4V��#���>�n�>���� ?G��=���<k=�����(E��@�����'�>?����#���U�gz���C�>3�?�Fo=��¾w�j������= �?A	<?�"�(&T��j�_�Y��5P�!���zb�����F�&��w|��W���R��vax�Q�/�~��;A�.?~�u?�N���������Jh�"90��,k>���>��>ͬ�>avw>�
���uZ�7�)�6va���>�r?��>��I?��;?�oP?�jL?���>l�>d2���L�>y��;���>���>f�9?�-?�10?Xr?Lm+?�,c>`�������ؾ[?)�?�H??��?�΅�
qý�N���h�O�y�=H�����=6��<W�׽��u���S=��S>r�?4�ս˞,�:���ɛ>�&?+��>��>m�l��������=f�?��?[��>� �X�x���!�3<�>�Mx?
�P�2�!=ejM>g��=���X�<��=E��_�`=�!I����ju�;��=I�~=��=�C<}�t�'6��l�����>�?2�>X��>4���� � ��(?�=�Z>�+N>T�>�ܾ_��O���7�f�K#x>�;�?��?ӧU=��=��=�$��(��V]��`���=��?W�#?��T?q��?��<?��"?�V>z���œ�lք��z����?�!,?���>��p�ʾ��T�3��?a?�6a����<7)���¾�Խ��>`[/��/~�����D�a���3��4������?保?�MA���6��u�9����\��)�C?�>�O�> �>��)��g����7;>�z�>&R?�>��O?��z?�Z?��V>){8�I��L㙿�o{���>��>?� �?��?x.x?î�>��>��(���}��c����$҂���X=��Z>*=�>4�>qĪ>B�=K�ƽ�C���J=�ȴ�=�F`>Ŵ�> ۥ>ro�>�nu>��<��G?�'�>�����@��:���Q���E�=Yu?6X�?��*?�*=��:�E�������>��?��?!�)?��S�a%�=!�̼E䶾qo�br�>F��>�0�>��=X�P=��>�W�>��>���#s��8�8�R���?��E?+/�=�꽿��v��J��<����_{={���C6��Ο1���T��}�>%qa�aK��A��KC���0���+B� �!�Df=�5�����>��=o�#���>���< �w=��-<�����=��<Scp��M���&��f�<�=��w��}C�<TP�;�:=8������?��x?EAb?M@?oI>�@
<��=-"?�z�ѕ:?),>~�������&�z_��.�l���-�]d���=k���<�9Ͻ8&=>��#>Bk>=�ܻ��G>HJ=�3�=|9���
 >�>(���> 82>?tA>U�[>�}?�m��DS����O�Gߠ�Ǎc?)��>�g�=�Gi�??sP�>x�p�#��%�}b?���?\a�?"�?�S��@��>�ɠ�Ӳ�����=����H����%>r�R�
��>D�~>�Z4��l��?�	�g��?	Q@��C?؈���Uܿf#$>x7>Hh>>1S��)1���Z��Ya���W�_� ?_�;��i˾|s�>��=��޾{,ƾ��3=�(7>DVg=��[[���=a�z�#�A=��h=pN�>��D>w#�=��i��=��J=��=-&O> g����>�-�3�7�-=�A�=.C_>�#>	
�>��?��.?ߤU?���>y�Q�����#/ľ/>N�><C�>�^�<�>>���>u�G?�X?��E?��>��=̱>�X�>t '��G�v��)􃾩K<\E�?k��?���>��%=�M���%�,=�i��_0	?��0?Ƨ?_��>.����׿+�����tdͽ�Y�L���z��i���ġ�>�۽�B:��|O��p�>���>���>�&>�2>�#�=y�>Ư6>"��;U�F��@Q��:���t���=~KR<fU=h�z=�Ǚ<%�ý"��݇ѽ�hռ�ۼ���=��ؽ���=ֶ�>
&>�2�>
ޙ=�{����3>$\��ٷM�Yp�=1b��(5B��ic��}�gn-��f3��eE>�}Y>X>v�gّ�|�?�pY>��=>��?m�t?{�!>1L
���վR����b��xT��Ͷ=��>�D@��[;��>`�!�M�xӾL��>n��>	�>Ȳl>�,��"?�U�w=��_5�S�>ex������$�6q�=?�������i��Ѻ֜D?�E�����=-#~?��I?��?
��>���$�ؾ�60>"B��U�=��$q��s����?t'?4��>����D�g繾�e��¿>7�ǽL��%���w.�������>pR����ξq�9�,	���X����D��G����>???]\�?���}�y��/R�ޚ��߽p>�>�Vw?/��>y�?o?�n4�^���6��I�=
x_?��?��?�)*>!��=S�����>&	?��?p��?"�s?
�?�oL�>+�;� >0����3�=��>f��=�E�=�t?�
?;�
?d��r�	������]����<��=��>B`�>��r>��=^3g=�x�=�\>Cƞ>�ޏ>�d>��>W<�> �\�",پ�^?�ۓ=T��>	�B?�7�>j�b�J��	2C>�����,�?/何T%<�����9<R�-=PЭ����<R��>�e˿���?��.>�� ���?=������U�>`�*>�3�,�>�X�=�5�>���>���>ɢG>RR�>Ɔ`>������%>�j��L'�Փ[���;���w�n>�C�iBe��`�l��������<���+�ܽd�O냿�I��#<���?齳:k�p�&��b��u?��>n�>?L<���ǽ���=�	?���>R1۾Nw������N��ق?���?�>".�>Uyb?�p�>5��A�</ri�X�}�$�f�+�\��5��+���<���о/��>��?�g?��W?��>�>`{?���2񿽜��=��F��Q[���=ה�>@����R�����,U����r��>��]?�H?�/�>\����C�5C>�5=?7�1?�~r?�`-?PZ6?n��\@*?��+>]G
?�~?"V5?~+?#?X!!>���=MՋ<$=o���w��[�+0ͽ~��]�&=���=�0<�$�:�n�<���;֪��<�Q�y;�4��ɀ<#� =;�=�^�=
��>�6d?���>��>�<?�v�Gt��
���N\>�k�e���m���I�#��?V@�?�ˌ?���>�O>��?�^鷽�P�=9�>�VX>���=���>�R��&�P�>n[>�N>-�Żq!��oX���tݔ��y����=��>���>5�J��1@>4D�<��)�>����:�PFA�� -�Εc�E��>�~O?� ?:�<> ���%=�0d��=?��?�8@?,(~?P*=�߳�`T���?���2��>�K����C��a���ˏ5�o4��y�h>j���%W߾���>[-��9c�����3�� �@���=i����.=�A���;���˾�>4��>�4��gI�칠��c����5?ێ =(�g��m���7о��=U��>
ie>�\���ԃ<��/�⍱��	T>$
�>i�=lʼ�!��a)E�IƾQ�>A�D?t�_?��?����%ar�WmC��D���e���uۼ�B?�ݪ>�T	?$,E>!2�=��0��Kd���F��s�>ŋ�>��GG����ns��b�%�VA�>A�?s�>�?�R?F?��`?��)?\{?Sp�>�b���.���A&?4��? �=��Խ�T� 9�OF�x��>q�)?9�B�׹�>N�?�?�&?�Q?�?n�>� ��C@����>�Y�>��W��b��?�_>��J?К�>l=Y?�ԃ?w�=>[�5��颾�֩��U�=�>��2? 6#?L�?���>c��>!������=<��>c?�/�?[�o?a�=��?:2>���>�ܖ=ޕ�>V��>�?�WO?"�s?��J?ܒ�>~h�<>���%��@s���O�H�;O�G<��y=��|Xt��*����<���;��������:�d�D�1��j��;9�>�BH>ڙ>���>J����Z�.�@==nϾ&�'7��Z��� `�=���>w�?*[�>�D�s!�=���>D�>-AO�3V?�>?��>�{=��Q��:X��2"�׼�=J�?j"�2a���>������7���k?u�o?LV��}�r�O�b?��]?=h��=��þz�b����g�O?<�
?(�G���>��~?d�q?P��>�e�-:n�*��Db���j�Ѷ=^r�>IX�O�d��?�>m�7?�N�>-�b>%%�=eu۾�w��q��h?��?�?���?�**>��n�X4�g~��'K���^?J��>�?��' #?� ���Ͼ�P��_(����S��>��sC���w��z�$�G݃�V׽��=��?�s?;\q?��_?{� �]d��1^�
���kV�Q(��%���E��'E��C��n�"b��.��>���G=�:%�e4/�3o�?h��>��C��>?��Ӿ}�0����<k@��;\&�kޖ>I��=�N>�f>���;ٽE���7�?�Y�>?�>@�6?�.���M�%�]���8�%��cI=n1[>1�>�B!?i[O>��5�9aѽXK�+}I��2��v>�xc?ݏK?K�n?WZ��1��x����!�_43�
��;B>K
>��>U1X�F�G&�e>���r���o~��	�	����=֭2?�A�>�t�>�<�?��?��	�?ͮ�[�x�ފ1���<a��>�h?P�>�_�>�|н�� ��r�>
�c?#M�>=��>�Nu�{��3C|�rw��,��>�#�>�U ?��n>��)��R^�h����ɑ�I�6��B>�`?�ș�C;����>�(T?��<D�Y��"�>�%b�i�!�kNϾ��H�*�=��	?���=$�L>��Ծ�����w�r��FO)?[K?�璾��*�h5~>Z$"?�}�>"*�>/�?�(�>�qþ��H��?��^?)BJ?�TA? I�>��=����(AȽ��&���,=<��>��Z>jm=ep�=E��qt\�,{���D=<v�=�yμ�L��)�<P����J<���<��3>F��<R��)���X�}:�Y ��5'��
8�\�G������˾�?���Ǿm���P�R��[3�bd��M��QU��^�?���?���7/ƾCٞ�Oe�,�~�l#�>���n޽NQ̾�3�{߼�T\Ծ���s�#���5�әD��U{�:�&?�現l_ǿ�9��� ���?�"?C[y?+����!�c�8��Z)>ã�<4ق����۟��+*Ͽ�)��1�^?��>�7�����>�1�>Dpd>�i>%N��K����S~<��?�/?FZ�>ۺu� ɿsn��|��<(��?o@�zA?��(�=����U=��>��	?�?>�j1�zQ�	��K�>�8�?��?�N=�W��	�ste?�<Y�F��޻�!�=���=��=����nJ>TC�>���fEA��Uܽѻ4>~��>vB"�����z^�j��<4�]>u�ս�*��HՄ?�{\��f���/�T���\>��T?�+�>�:�=ױ,?W6H�}Ͽ0�\��*a?�0�?���?��(?sܿ��ٚ>G�ܾ��M?�C6?���>�d&���t����=�Cἃ"����㾟(V�$��=	��>��>�|,�I��R�O�.I�����=#��3�ǿO�"������< *����Z����(�Ľ��Z�9��س\����m��='?�=CO_>uNg>�/>BZP>�a?3�m?�	�>U, >���ᇾ-溾х���]��{+�>藾����Ա��ྼ㾜-�>���m��~Ӿ�BF��]�=n�\�ߜ���1��$^�k�$���?m/6>��˾èN��Ɨ=���R���$��0��־��1�4z���?FAM?@����?�
��������.Z?�����������+>�M,���n<��>$�N=N�Ѿ��"��
e���1?��?�ּ��ڕ���/>0F���6�<h�+?f��>��<g̬>�#?h*������>>{/>>��>���>�p>`��Sƽ�?�4U?���&���3�>�i������[�=���=��3�Z����f>�R�<}������Ξ��ܷ<m�f?��>�\���"�[�d��晽QR0�c�|?`~$?�k�>۲�?Q�?	��7�#����㾪q?>)qW?��G?��$=��=�N �w��΁>?��^?��(=_�Ͼ�G;��q���'��8?�ID?�?�|����eW���/ ��>?��w?F<j�y졿���v�����>�d�>�d�>w1+�K��>f
I?F.���R���񹿦G5�ҷ�?�@��?Is�=GH����<Ŭ�>}�>�(�ɾ>���C妾��=�� ?�]��pф�ó$�L�V�L?OD�?��> �¾���=����_�?�҆?�]��3dn<)D�l�( �t�<5��=J��X��"���t7� ƾ�
��_�� ����e�>�;@'-��:�>�l6��2�fdϿ
���о��q�n�?i��>�Ľ�ۢ��~j��<u�¦G��vH�rT��r��>��=1]=s���:|��_7��S=r?�>�I=���>�z,�!�d��iK��-��>��	?f��>�X����N��?#�����B��Z6�w@?g��?)��?��M?37R>�S0�@��G4���?�I?�W?�Hb��B��T���j?MO���B`��4��,E�2U>. 3?�N�>��-��~=#?>�~�>�U>+/���Ŀ.ݶ������?�y�?ޒ�S��>h��?�{+?FS��2��!3����*�?�Z��FA?�1>����F�!�y=�������
?�V0?.��7"�f5d?k�j��>u�ox4��1K�)��>��-�o�)��ۼ�� �k�T��꘿@�_��~�?�~�?>��?s����T(��R'?*��>19��M����M$=�V�>CF�>X�2>X&��S�>t����W�k3>���?��?J�?>Ö�3P��@T>6cu?0Ӳ>�z�?�^>��>	GS>�����A��W�`>�.I>�Ar=j��>�8?q:�>�؈��l��hNC��H�G�6�bI�zNb�y<�> �V?��d?��J>��ļ�mD=���p%<io���4��Alc��N��K򽢨�>TV�>�E/>��W����"?͵(��lֿ�����`1�kY?Z��>y?��澙)�����=_�?��>*U�fI���:���Ƨ��}�?���?O�?ە��΀���==�� ?���>�����ϯ���6�B�>g@]? ň������p�Z&6>`��?*@���?lb��j?���<����������D���L��=��6?��6W>�k?�	>��o������u� �>^j�?�.�?�L ?�Wj?�s��t8�U�G=���>9}f?x��>�oW;�Nݾ�TQ>�?q��/A��u����Mf?��@�@�+J?���yhֿ����xN��\���c��=���=҆2>��ٽ^�=.�7=��8�&?�����=c�>��d>Bq>W(O>�a;>�)>���F�!�r��R���B�C�������Z�B��*Xv�Iz��3�������?��G4ý6y���Q�2&��>`����=��U?$R?g7p?# ?
>y�=>>߾��\ =��"�dۃ=���>�O2?�kL?L�*?�x�=�>����d��@���4���͇���>�I>S��>Q�>��>+ �9#~I>$�?>hW�>�� >_t&=���R�=�O>��>��>[^�>��'>=&>f����+���jr����o�d��?b=��=C����1��
%�����=��)?�T�=V���Կ_���vH?�[���?�ET�'�=G::?t�W?�(>`
��-���22->�Jͽ�`���
>|I�3Dg��"'�KpU>��!?��=�C�>��?��-��^�&H��ì>�c2?��t���Z��u������+hG>�
�>]�ν��0��I��m���C��� �=��1?k�?['(����mӍ�J�;��Vm>�W>S��:��;��>���:O�Z=��:�1G���A=�R>D�?B�1>�7�=�W�>����KQ��أ>j;>'�>�@?1�!?E�K��c��eч��2/�Ds>�-�>Rx>�i>�N���=^r�>�Hh>�ۼ����3���;��9P>r)I�8!c�o����<p=@���e#�=ด=�k�#+@�C�!=���?�ٮ��l����� Th���a?f��>�=ڠ��Q�2�������g���?l�@�f�?b���R<�T?�?R�$��:�=|��>�b�>3�wž�?�m���;?�����f�?(�?04y=S���Bi�D�S=�<?3�徵��>~���&������:�~� ��=~� ?�oH?��䦽��e�w:?���>��ž%����?οq
��1�>��?'��?f���S�����I� �!?���?M�?��H>�ۺ�/�{���>�fE?K�K?�WK>0�(����*?`��?�ٔ?bI>���?"�s?�k�>�/x��Z/��6�������k=̀[;�d�>W>����MgF��ד�kh��D�j�}���a>q�$=��>;E�4���:�=��I��ۻf�2��>�,q>�I> W�>h� ?�a�>v��>�w=�m��$ှq���}�K?���?���2n�O�<o��=��^��&?cI4?o[��Ͼ�ը>��\?o?�[?&d�>C��E>��>迿3~����<<�K>-4�>�H�>�%��/FK>��Ծ�4D�Gp�>�ϗ>�����?ھ�,��9S��&B�>�e!?���>�Ү=� ?��#?�j>�(�>1aE��9��\�E�ɲ�>բ�>�H?�~?��?�Թ��Z3�����桿��[��;N>��x?�U?�ʕ>V���僝�iE�[BI����U��?}tg?�R�?62�?�??a�A?�)f>#��Fؾ������>]�!?B�H�A��M&��W~?�P?r��>T:����ս�Pּ��������?�(\?pA&?Ŝ��+a���¾k4�<��"���U����;�D�f�>��>�����=>gװ=�Om��E6��f<1i�=c�>n�=/7�\u����,?j�p�P\����=�sr�yD�OI~>�R>#���_?��5��|�'����w��:Z�'�?���?+Y�?�<���h���<?S&�?�~?Ʃ�>����J�ᾃ��v_x��}�G��_�>˪�>٭W���澲���MS���ك��ƽ]+��Q?=N�>�O?<?<�A>���>� ��>m(�9P��'u��yb�`u��D9����� �
�d�I���WM:��Ӿ�b}��ܰ>���֞>QA?�S*>�>
�>��2�.��>�)>/`>��>��>~77> >4>�5e���T?xB⾜�&��7��,��`�@?��\?�_�>^��(3������L.?�?Ş?Hƀ>�ca���!�,�?#y�>����!?�W�=�߼e0p�bE۾ww��z�T�ΌB�_��>#N����+���X�@����>.�?ϼ�<Ʒ�Ѩ����=�n=N�?��(?�)���Q���o�θW�S�0���6h�Mj��P�$� �p��쏿�^��%����(��r*=��*?j�?Ќ����!���&k��?��df>_�>a$�>,�>"uI>��	�r�1�g^�M'�K���gR�>~[{?ZN�>:�I?�<?Q?��K?��>~o�>�ʰ��-�>=D	<��>,Z�>J59?D-?�0?�|?�+?�`>� ������Xؾ�\?|�?�=?+�?��?�k���'ƽ�}��w�7�z�����av=eq�<J�Խ�|f�(xP=R�S>�X?����8������k>R�7?��>���>e���,��� �<��>ŵ
?�F�>! ��}r��b��V�>���?-�	�=M�)>���=4�����Һ�X�=�����=;��>x;��g<)��=W��=-�t��-��P��:劇;�m�<��>�?r��>*2�>�V��� �1�����=-�Z>8T>��>H�پ�e���$���%h�ZRz>��?�n�?2�f=N��=���=����ݿ�T������99�<:?��"?��S?�q�?��=?E,#?p�>�N��R���Y��������?�!,?2��>���!�ʾ"憎T�3���?�[?�9a�Y��o8)��¾�Խ̥>�^/��1~����rD�r	������m��}��?ݿ�? A�Z�6��r�𽘿�[��4�C?��>�V�>��>��)���g�=&�,";>��>

R?�n�>(P?6u?X-/?���>�1�C	ɿ�k����ξ�㾅�!?WR`?d�?�?�?��5?������<<'<�G��B"���ͽ�&���.�>�3E>�Ap>�d�>-@>{p�>%�[�� <ʾ��ۏŽ��l>���>E�d=���>��E>�N�=�X?j;:>�����1������̫�A�>2=�?kS�?)nz?P��>OGg��t%���.���>���?�?fY/? ;��yo�=l̽�2��#���}�>$Y�>����C�>c$7>U�S��g?Xg�>��Ͻ���‿lD�N��>�EI?SHl�̨ſ�zo�.x�����eT�;�o��`�[��a���W�n�=y����P�t���d+Z�Mu��&+��0y���Y"�����>�*�=3��=Kq�=e �<��
�X�<�b=r �<2�=�eu�׋�<��1��@��]u�9<c�3,&<*�F=��Q�!�꾠��?FK?�)?�g?#�g>�]�=XO>(�?���=�~>?�w����E�n���=�9.�����d��A�Y˾Ϩ����=�P��"�=�4�=� >�������<�kh<AS6>ᘟ<�z�=�c�=٢�=���=~�1>r{S=�jZ>Fo}?$w��!���T�{��;�e\?y,�>¡>ͯ��gw-?��>7�}��)�������i?���?�)�?{s�>���;��>(����6�i3�=�y~��}�=���=�^'��>��B>2����
r=�}�?I!@9&?�|��]�ֿ�>�h5>�>�S��41�S\��d�F�X� � ?�#;��˾h�>9]�=��߾�8ƾ��4=�5>�^=����$\�mi�=��{�Y�A=�Dr=�x�>s<B>L�=6D�����=ٵF=Xj�=�ON>!B�9�G�.�z�-=���=aV`>R�%>M��>{V?�$D?�d�?(}�>p�u�<�;�ؾY+>#}>��U>�����$>U�>�<?2�J?c?7V7>[�)>�>Y��=���Hj���6N��RV(> ��?b�?���>�=�� �uM�~&&�C���ݿ?I�?��>�&�>���`俞D#���(�1��������@<�a��宽�6v<Á�H�^��]�=��>U��>�}�>V8@>�m�=���>Ն�>A>���q
>��������&��<i�Ѻ#�Խ�Y������*Y���@<Q�V�/=G`ӽr2_�U�p��=�d�>]�=}ȴ>��=���.>�	��4wQ�7>�=���+�D�ݖb��Dw��Z$�[��HV>V�l>�c�[=���?�C>�PE>�S�?�mn?�
>�9ٽ�ؾ�ꚿ�HN�L^k�|��=��=�W� �8��[��JI��tľ{��>��>Z��>!$;>��xr4�/�޻�נ���$F?C(d���2�c��m�i�>������lDh��d�;\05?�_��iXG>�`�?߄b?~�?[�>��=$S˾��f>{��;���$.��x�#�㼌_'?�:?�!�>`	��6�]F̾���=�>+<I�q�O�b�
�0�Yu��ʷ���>�����о*$3��g��#����B��Fr���>K�O?t�?�>b�yW��QVO�$���(���r?�~g?��>FL?�A?�+��?y�=t��o�=��n?	��?H=�?�>J��=.���q9�>;-	?侖?J��?�~s?�?�1l�>�G�;� >*瘽$=�=;�>���=><�=�u?��
?i�
?il��L�	������H^���<4ɡ=��>dn�>�r>���=��g=�v�=Z)\>՞>�>!�d>h��>�N�>���������?��F �>�0?��>��������P�.��Si���P����?ܔ�Iӽ���=��;��=`��=��>=�ſI��?ި=i-�ݠ?9��L��=�(W>$�==+�꼚��>Q�>pH�>���>���>1�9=�aP>�M=(�ȾB�H>Q��SN�0u���V��5��x��>�ɍ�)���������PL���Q�,龘*c�Fي��l�Y��z��?Y�<�\�YL�^�^��X@?-g�>�O5?̓��s����>
�'?G.�>6澭���&���������?2�@�`>���>�UY?g�?�Z*��A8���W��u��E���Z�b�`��я�NG}�������:_?�|?L#7?8F=�z>L	w?��������Ӊ>h(,�&5�J`P=�٨>Ds��6�`��ξ�sþ����I>Klm?5l�?F�?#lR���m�j4'>��:?�1?Pt?��1?�;?L����$?Un3>�H?�n?�J5?��.?��
?�2>��=Ep����'=�E�����ѽ8�ʽh-�\�3=Dj{=����-)<ܝ=�ޥ<��|ټ�;�����<:=ޢ=�,�=>�>�]?R��>��>@�/?&�&�I4��콾Ӓ? �=C���f�����#���K�>��g?��?�4D?��>� ;�-�Q�r�M>ڐ�>�0>: C>��>)�νޟC�w3�=n��=L�>ial=z����@q�����lU��E�;Q�>�3�>���>!��̚�=p��=U\���X>,Z���پ	T'��H�Td3�,O��@��>sH?�!?Y
�=��ľ�μ�q�]?2?�2"?�8E?�m?�K�=N۾%�#��K����5�>s������GN���ٛ�J�.�魜<�U>����0D��G[b>�����޾��n�%J�U8�`GM=�?���R=1X���վ��~�An�=f�
>�b���!�� ���ת���I?+&j=����aU������G>�ޘ>��>��;�1�x���@�ǽ��͖=�n�>z�:>\���9ﾬ�G��%���>O�D?_?���?kJ��Gr�V�A�Zr���a����S�?�;�>��	?��E>/�=�E��N��kd��cH�E��>���>����F�1Ǡ�����f"��u�>]�?o�$>��?�S?1?qm_?�*?"_?�=�>�c��M'��S�'??�?�S�=	QͽNt�>p=���A�l?1+?�樽>H�>ϳ?h ?��(?��N?�?�T>y�ξ�;����>ɿ�>K�T��갿õ�>��B?�h�>��T?B�?[d>)�Oe���_4���>�O">�|3?�&?��?I�>˔K?6�y�+�f��Yt>mA]?Ws�?��s?���>��?�h��
5?Х�>�HY>�=?_!?g�n?M��?."w?�'*?���=�փ���ҽ��A�	ck��*�=���=W@�=H�<yYR��K	>���=���<m��������=.��<6�=��W=&_�>��s>�	��C�0>��ľ)P����@>�v��Q���ي���:��׷=���>��?���>|X#����= ��>�G�>��X6(?�??P";��b�0�ھ�K�Y�>z	B?+��=��l�(���U�u��h=��m?��^?�W��&��O�b?��]??h��=��þz�b����f�O?<�
?4�G���>��~?f�q?T��>	�e�+:n�*��Db���j�&Ѷ=[r�>LX�R�d��?�>o�7?�N�>4�b>$%�=gu۾�w��q��i?��?�?���?+*>��n�Z4࿍P��%Ӥ��Bd?�t�>M���8?�����侳�������=ƾ"$S��ᚾ@þ_.G�m��m�����L>Â?�W�?��f?8�k?ĬӾp5p�k\H���x��:K��'��4� �<�:�^��L�{=l��$�	������ؗt<�}���lF��?��&?:�1��/�>{���X��BʾD�O>r�����	����=���N�c=��^=�zb�4�&�hb���j ?dx�>���>o�=?a�Y���:���-�
8�����,>%f�>��>e7�>��W�6g)�vi콗�˾�Q���\Ͻ-�g>!�X?��??7�N?���<	�������_�� �ӱ���2�==A��V.�>�<h�����~;�ת-�?f�5�)�Y�]��u����<�L?�:�=�x�>�	�?7�B?l����.��R���+�Y��>�L$?�j�?�?X��>�w��t?����>��l?��>�Ϡ>nE��5M!���{��*̽�>��>���>�co>!-�� \��w��م��W9����=�h?ji���a��ȅ>yR?Bc:;EJ<�v�>(u�N�!��򾨼'�
�>�?�ݪ=�(<>u3ž
!��{��x��Di)?)8?P��F�*�be~>;"?v��>�?�>},�?	�>�þQż�Ҧ?��^?r2J?�aA?��>� =������ǽ5�&���,=�|�>��Z>N�l=���=��=\�i:�<�D=�d�=%�μ`���?�<�����%H<�E�<4>@mۿ�BK�s�پ�S�v?
��爾c����c��ݲ��a��6��ZXx� ��J'�kV�k7c������l�Ї�?�=�?"���p0�� ���=����������>{�q���������j)����n���ed!���O��&i���e���&?#���ǿ񶡿�Oݾ'T?+� ?�y?�7���"���8���>��<�u��2��󔚿fϿ����}^?���>������R��>Q�>(&Y>�o>h���ɑ��佥<�%?e�,?��>m$s��Wɿ����;o�<s��?��@�|A?��(����*OV=���>�	?`�?>�X1�`J�����bU�>�:�?y��?��M=��W�I�	�xe?�z<��F��Iݻ��=�;�=f<=`��l�J>V�>o���NA��6ܽL�4>��>�i"���~^�P��<o�]>��ս�#��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=W��3�ƿ��$�L�	=��ZC]�,G�H���R�O��ܟ�EQn�*����e=��=oQ>�r�><�W>�
[>�`W?r�k?5��>RS>�㽤����;4
��j���K��������1��B��T]߾pr	��������ɾQ�K�W�=;bm�,g���?���i��q���?�ؐ>�d���)j��3�<���i��OO�=\c=O���B�C<{��bR?W"?�����(W�X82�ON����<�OA?�䶽��|N� �T=�q/������>��X5�_e��V��r0?�Y?�y��
J��0*>)� �!�=:�+? �?�t[<�(�>M<%?��*�g��&S[>��3>�٣>!��>	>��`۽߉?��T?������j�>d^��T�z���a=�O>�<5��v���[>fY�<�匾W�S��@���{�<�(W?n��>��)��na������Y==��x?��?.�>v{k?��B?�դ<h��u�S����bw=�W?4*i?��>�����	оX���?�5?٣e?��N>�bh���1�.�]U��$?�n?(_?=~��"w}���d���n6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������*�l=M��F�?��?������uO���s�{�E���a=*�Z=ڠL�Í��N"����'���x�� �=�~�>��@8Z˽��>44�<	��п�~�ߚ��XS˾��?�9@>P-���ߒ�ٌ��g��SyL��SN�D���M�>�>�������+�{��q;�k#��s�>�	�A�>�S��%��옟�L�5<�>��>S��>�%��d轾bę?pb���?οJ������;�X?�g�?�n�?�q?t9<��v��{�v��.G?d�s?3Z?Bl%�3=]�P�7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?]$�>��?o�=�a�> d�=P��-��k#>y"�=��>��?��M?	L�>nW�=��8��/�B[F��GR�`$�@�C��>��a?�L?Kb>*���2��!��uͽ�c1��P鼩W@�G�,���߽C(5>��=>�>_�D��Ӿ��?Mp�9�ؿ j��p'��54?/��>�?����t�����;_?Oz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>B�Խ����\�����7>1�B?Y��D��u�o�y�>���?
�@�ծ?ii��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?pQo���i�B>��?"������L��f?�
@u@a�^?*
?��[N��L���~z��*�=��=�4~>�y�'�%>E�j���R��	=��>��>��>��>S'N>�bu>\��=���������cn����i�R9��]Ҿ�"��g�վ���IqK�W⸾���:
�k��\�0�C8þ�uǾJ�u�MB>�<?"�L?��?���>�p��Q��=a�p8��I=��>��ӫK?��_?�]?8�>�T+��nQ�ύ��o�Q���|��,�>3.�>_��>���>>z�>�PK��U>2��>��>P�~>[�	>gz��>�	>�u>�۴>���>�H�>$�6�reN>U���r��%I���پp�>�?�H� Bg��������u����,<�}.?�t=U����ο8���Od9?n�]�u��k"ཇH>�{?!:8?���>rB��2��A�H>hJ_�pd���{ϻ��r�aq	��u3�y�>�s3?`��\>ɍ6��7�3�b�K���Ch�>�HG?5�1��w���{��\�Z��6ȾЄ;���>��e���I�ʏ�3aO�j�b��Oؽ)�y?)?�yU>7�����E@��Ƴ�<�>�w#>����|>_�e�)�E����<E>�o�=��{>�U?E�+>��=��>Q���UP�$q�>��B><�+>E@?�'%?T������U����-�.w>�[�>t �>w�>�3J��=�b�>u�a>������0r��?��zW>v}�0J_��yt���x=G��:&�=Oh�=�W �A�<��O&=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾOh�>zx��Z�������u�m�#=S��>�8H?�V����O�i>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?roi>�g۾8`Z����>ѻ@?�R?�>�9���'���?�޶?֯�?�d�=�8�?�~g?�#�=&��>oX������M����=ȼ��q�0>�Վ��6��Y\�`����B��P�C�a� ��O>X��={��>Z�^�b�Ծ1�A>5F�=9\2��kB�>��w=�=��V=�G?[�>�V>27�=iͼC�����쾰�K?��?���80n�^�<��=/�^��'?�G4?�=[���ϾKШ>M�\?�?M[?d�>����=���迿�|�����<��K>�6�>G�>G(��>NK>.�Ծ'6D��s�>`җ>z��%=ھ`'�����4C�>Ff!?���>oǮ=Й ?��#?��j>�(�>2aE��9��c�E����>̢�>�H?�~?��?�Թ��Z3�����桿��[�V;N>��x?V?�ʕ>^�������gE��AI�k���U��?�tg?HS�'?/2�?߉??Z�A?)f>ه�ؾĩ����>��!?��A��F&����+{?M?=��>�N����ս�ּ���Zr��C?]$\?@&?)���*a�i
þPN�<#��5T�Y <��D��>-�>�����}�=&>���=Om��:6���h<>��=��> %�=+*7�c���0=,?��G�~ۃ���=��r�?xD���>�IL>����^?kl=��{�����x��	U� �? ��?Zk�?b��@�h��$=?�?S	?m"�>�J���}޾6�྿Pw�~x��w�Z�>���>$�l���K���ڙ���F��_�Ž��9�|g�>���>/�?xn�>S�/>5w�>f���u2�@�����be��d�7�r$$�N����2[=��Z�Eƾum�� W�>3
R�4[�>V�?�/>!>u��>�㙼Zђ>�6>N�~>��>��]>p4A>�c>�O�<�}���KR?����$�'���辿���g3B?�qd?U1�>ii�<��������?���?Ts�?=v>
h��,+��n?�>�>G��Vq
?uT:=�8�;�<V��w��3���1��>E׽� :��M�Enf�wj
?�/?�����̾�;׽{�����=?N�?� .?���,3T� �x�j1_�ZI������M�H����98�"`v��ܐ� ���̲��	'#�~��=�y$?�я?h6 �����{��Z��D��jA>���>�	�>�̷>� >/�
��$�P�r�Dn%�*�^�^]�>�f?���>�qI?p�;?ՒP?�XL?kz�>�(�>�˯���>N��;��>|>�>�9?o.?�0?�n?�k+?��b>�J��i���8rؾ�?G�?:'?��?��?9 ���ý�����]\�YJy�����P�=�g�<��ֽ`�r�edU=X�S>Z?m��ڬ8�a���k>E�7?���>���>k���,���;�<��>e�
?�I�>(  �H{r�q`�QZ�>���?�����=~�)>���=������Ӻ�Y�=(���D�=V$���;�eP<��=��=Tt���z�i��:9�;(��< u�>6�?���>�C�>�@��/� �c��f�=�Y>=S>|>�Eپ�}���$��v�g��]y>�w�?�z�?ѻf=��=��=}���U�����H������<�??J#?)XT?`��?{�=?_j#?е>+�jM���^�������?%�%?U�>�U�a�Ͼ�W��T5�V|?��?�f���+���ƾ~�߽>K�=��*��F�u����C��Մ��������g��?'�?�4Ҽ�I1����Ֆ�����-F?��>��>��>�='��c����@>��>*�O?�5�>5dO?� {?�\?��T>|98�@���Tv��l��P%>��??@р?B�?��x?տ�>~�>��'�F�߾9T�����������?Z=�"V>�.�>Y��>g��>�i�=���y��5�9�	��=B`>��>@��>�><�y>�s�<8�G?�\�>���|e�Nת�PŐ�n?t�H�z?�ː?�6?`
g=�;���;���A��>C�?���?f�2?�5U�� �=��&��h��������>�$�>���>��=g9�=)e�=ѵ�>�ɿ> {O�9U� �2����[<?8�F?�?�=��ſ��q�0�b�i������<k�����d�Ch��ZH��~�=�֑���&����j3N�	$��Մ������.f���fo�'A�>S�==E4�=���=S$�<��(�G��<�U�<�M=q�=|//�Ӭu=�W����o����T�:�x�<��B=�J:1�˾�}?�;I?ܕ+?��C?�y>;>��3�M��>�����@?OV>/�P�������;�J���� ��S�ؾ%x׾��c�ʟ��H>c`I�#�>�83>�G�=K�<D�=�s=�=<�Q��=$�=�O�=wg�=��=��>HU>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>`�7>�+>��R�3�1�ɾ\��b��YZ�W�!?&M;��K̾��>*��=�&߾n�ƾ	�.=�e6>u�a=Az�GR\�]�=�{���<=�\l=݉>q�C>�R�=�1��q~�==^J=;�=3�O>�ŕ���7�� ,��}3=n��=Y�b>j&>�t�>�U?�7?i�w?��P>KW���뫾�n���>��>���>�k�=�|�>F�>�g%?�I?�yP?:0�>:k��K;�>� �>�	�Z��$���!��چ�?�?��?C�>���<��u=;�����,? �B^?��B?lR0?��>�B��k���%�Em.�_ח�4io:�r)=ׂp���N����`���P�=��>���>n�>?�x>E�9>H�N>�>��	>N~�<"Ʉ=IӔ�ƾ<}���n`~=p�k�p��<S	���f;�S����(�҄���ߘ;(�;̨Z<���;S��=���>�<>���>���=���B/>v���b�L�[��=&H���,B��4d��I~�/��W6�صB>�9X>�|��4����?��Y>�l?>���?SAu?��>\ ��վ�Q��!Ce�FWS��˸=ֶ>��<��z;�bZ`�:�M��{ҾP+�>IR�>Pf�>[xk>,�UH?�HAy= r�ts6�MD�>�b��F+�e���)q�"���p⟿�Ci�~ʑ�&D?t����=��~?%�I?}�?,��>`=����׾	0>�u����=j]�J�n������?�'?k	�>2�뾇D��H̾C���޷>�@I�-�O���W�0�(��:ͷ�2��>������оn$3��g�������B��Lr�N��>$�O?��?M:b��W��IUO����,(���q?�|g?0�>�J?�@?5&��	z�}r���v�=�n?ɳ�?N=�?t>�5�=�I��x��>�?�?>��?�fs?�B;�>k�>�T`;\}!>Vї��=Ci>�=��=:�?��
?�6?����0�	�K񾫜��#]�?��<Į�=���> ��>�r>�s�=�qj=���=JPY>���>'��>�eh>WK�>Lˉ>���"�N��}?(f=�P>�V.?���=g\=��=�!>	>"=�2L���ۼ7eO��l<}w���<z�=N%>�v ?_���W��?�0~>N����3?#ξ�^���M0>&Y�>o׬���)?$�C>�I��G�>���>�pR>��>��>eؾ��>S��X$�PG�ƊT�Rľ���>0q���g7�G\��* ���L�����&6j��m��	>� Ē<&&�?|���d��>&����l?0ݣ>U5?[�+�Q���>���>=��>�����e��7䎿S����?P��?�;c>��>O�W?!�?��1�e3�vZ�4�u�b(A�'e�A�`�}፿���	�
�M����_?��x?yA?+T�<+:z>Y��?��%��ӏ��)�>�/�'';��?<=o+�>
*��"�`���Ӿ��þ�7�=HF>{�o?7%�?ZY?_TV���m��'>��:?J�1?XOt?��1?ʌ;?s����$?�m3>lF?[p?�M5?��.?��
?�2>c�=n৻o�'=-3��u����ѽm}ʽ���J�3=S_{=���uG<L�=E�<�`�"�ټ/�;�(���.�<�:=��=� �=���>;�]?@O�>٠�>��7?:��Ov8�׺���&/?|0:=!���F��9������>��j?���?�aZ?�Cd>�A��C��>xY�>pu&>\>i�>ϔ���E����=�U>}]>���=pBM�=ȁ�'�	�����1�<i)>���>M0|>���!�'>�|���0z�R�d>�Q��̺���S���G���1���v��Y�>1�K?��?���=g_龏-��eIf�-0)?�]<?�NM?��?�=��۾��9���J�>>���>)Y�<�������#����:��K�:��s>2��{���7d>@����4�n�A�I�~�ʍ`=�v�r"B=+X���׾�������=o>>�=����!�����媿�J?��}=b���>X�2ػ�$�>;�>㩮>~?��tq�~@�_��@��=��>��=>1���zﾧ�G�ߺ�葈>�cS?�w?}i�?s��5g��-Y]�e�B�+�g���>N��>n �>�.?��>X`'>�Ww��޾�k�j�R�+|�>�!�>��I9������ξ��T�Xj�>�V&?�+:;�x.?�Z_?v?L�b?�8?5�?��>"w�l@���0(?���?�l�=����'L�s�X�ކ]�5ɽ>o04?/�ٽG��>�!?�=?8a6?�}B?��?]Tk>�+�(�c�)��>f׀>,􃿩G���N>��2?���>�G^?I�i?x�=�4d��4
�dy�=9�	>��4?��4?��A?�h�>� ;?�� �G<ž�́>��9?�s�?ǯJ?4��>kK}?�P�=�O�>5l>�$�;��?MK?-)t?��?�`?��>b�L����.����������0�=l��=��K=ob�,���#_�=�q\�8�-6���+�=LS�;2\��/�=�_�>��s>���7�0>u�ľcO����@>p����N���؊���:�n۷=G��>��?���>cW#�纒=���>wH�>h��v5(?t�??4";�b���ھB�K���>�B?^��=��l�*���1�u�Lh=N�m?ы^?��W�Z%��O�b?��]?@h��=��þz�b����g�O?=�
?3�G���>��~?f�q?U��>�e�+:n�*��Db���j�&Ѷ=\r�>LX�S�d��?�>o�7?�N�>/�b>'%�=iu۾�w��q��h?��?�?���?+*>��n�Z4�d����Pc?���>��?+ ?Ǣ��ѽ��ޒ���y�"��-���/��꠾�ן�*v"�N�v�6�����=�?�_q?WFm?��c?=��6<b���^�	���\�Ů��b%�V�=�{3A���L��em�����W����>=	pw���E�i$�?�B(?�����>D����j¾�:վb�o>v���X�s��=4L��bs=��E=�;��d����Sg ?��>oG�>�8J?'�D�Y�:��f2�J�@��2���l>��z>���>��>��mu2��n�y/��_������c:t>�.c?�N?pn?[R꽮�/�x��s�"��RV�2�����>>Zg>�Ñ>�L�`��7%���9��Rq�{���K��H��,jz=y�1?58u>��>�h�?��?^u�������v��1��[�<��>e�g?���>�>֮ҽ���0��>��l?ª�>��>�����Z!�;�{�ܮʽ�$�>�>���>��o>ì,�U#\��j��>����9�8r�=4�h?!����`��>R?�:�G<�{�>��v�D�!�����'�4�>�|?���=��;>�~ž$�¦{��7���q4?��>��o-'�@�`>�'?�$?'I�>���?�6�>�V���&8�w�?0"V?ցG?7G?(�?���=��#����3'���<��]>���>�ƹ=�T�=HB8��p�;d׽2'�=�	>�(��/b�1�S�I.��m\~=R�̼(�>�Lٿ@I��E��%�o�޾�o��{����0��C67��/�$k˾�e��@����^��+��8��}����t�}��?�r�?��/�� ��ʥ�앃�Pvؾg�>��h���<�͑Ͼrj��|����a���6����x��̌�*�|�S� ?��J=��������P��?1?* >?��ؾ��l�C�t�qV��Wm0<�A�����|)���߿ox�E&X?g~�>7��%�=�<?��d����>V?w��)轿Jľ�Cϻ0�8?��:?�.?�mǾ�.���ѿ�V>E+�?��@_�A?Q�(����dW=��>z=	?qu?>lb1�U�����/w�>�:�?(��?��O=d�W��e��e?v�<�"G��ܻ���=b��=�k=�m��K>���>���+<B��Nܽ[�5>*ޅ>s�$�@����]�߻�<��\>��ӽ� ��aՄ?Fz\�hf���/��T���U>X�T?/�>SU�=�,?�6H�x|Ͽܮ\��)a?�/�?���?��(?�Կ�{ښ>��ܾ�M?YC6?3�>Ee&�7�t����=^2�@�����o%V����=o��>/�>S�,���ҀO��g��7��=�����ƿ$�'��	��3=�ş<�c0��ؽ�d���S��֫��蹀�I� ��=r��=Q�S>�~>��@>��_>�.X?6�t?�;�>Ur�=�c�5Z��e#վ�H�<�zp���G�7�����V�Ś���>ݾ�~پ*�� �"�$���ؾ�D��7�=��H��ǚ��(���`��*���;?���=����se�����x�$a��6�A;��Q����S�Q�g�u�N �?��e?�vo�X�z�l7�>_)����<}�^?~�4�l�
���о�	�=�z�p�.�^��>��=Ȃ�)lX�O�]�F�0?\?�����3��
*>�*��=@�+?8�?�]<gG�>�H%?ɀ*�])�'�[>�(4>�>���>��>a����۽Vj? mT?ӎ�#���:�>�a���y{�)�a=�>�#5�x�꼂~[>�|�<�㌾�A[�]����ſ<�+W?���>��)�n��^���z�B�==V�x?e�?~4�> vk?��B?���<2Y��^�S���_x=��W?Y&i?�>����#о݀��8�5?٢e?i�N>�sh����-�.��J�A'?�n?9_?쳝��n}�r������f6?��v?s^�ws�����R�V�h=�>�[�>���>��9��k�>�>?�#��G������tY4�%Þ?��@���?�;<  �Z��=�;?`\�>��O��>ƾ�z��������q=�"�>����}ev����R,�b�8?ڠ�?���>������|�=툆�Q�?�?�^�0�����`T�9�� i>���sV�X�W��H#�\�+�V"߾�-��Ҙ��K=�_>\�@�F��T�>w��kϿmÿ�B��Z	�Q����?�ʬ>�~ɾY���t�� ���U;v�F�n�ਾ���>γ
>q���1���8�x�f�9�3������>�����>ϸK��P������{�<c�>��>nu�>a����1��ՙ?���.�ο���nS��FW?���?"��?�
!?h�;��w����� Z��aE?ǘr?b�Y?-r���U��2�
�[?N>���H�R.D��`z�+֎>���>�? zH�������>��>��>n&l��qԿ�ſ����ٖ?���?��۾K+�>Ew�?]J1??�Ӿ�繿��`��: ��1?<\�Q?w��>C乾ݘ@���8��K�z?|(Y?���=�8L�]�_?+�a�N�p���-�~�ƽ�ۡ> �0��e\��M�����Xe����@y����?M^�?h�?ѵ�� #�f6%? �>f����8Ǿ��<���>�(�>*N>RH_���u>����:�i	>���?�~�?Qj?���������U>	�}?#!�>M�?��=n�>�o�=�����-�?E#>0��=��=�ɘ?
�M?R\�>�{�=��8� /�TF��GR�$�Q�C�c�>�a?K�L?�1b>HV����1�!�UOͽ~P1�p�|]@�P�,���߽'/5>��=>x�>H�D��Ӿ��?�/�Reؿ\n���>*�(�4?,��>�p?�#���u��	_?)��>���vZ��6]����Uc�?���?��?��׾�Y��=c>_�>���>�Aս�U���Ň�c�8>.�B?7��@���p����>���?r�@�?9�h��	?���P��Va~����7�_��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>!�l?��o�O�B���1=9M�>̜k?�s?�Qo���k�B>��?"������L��f?�
@u@a�^?*XZҿR���p��24��m_�=��=H� >�3꽹D�=	��<���<�Ϊ<�ݐ=Y�>5Nb>�p>��R>��R>�P&>+���A$��ש�SH����=���T"�0�R�C� �s�]�%�����adξjn���.Խ*݆��ES���+��8��0��=I�Q?�Z[?�{v?/ �>���ey><
���2�ν	=�j�<��p>�.B?leI?`8&?�`=6ʋ�=�b��x��욾�2~�/��>lb�>��>&֗>4��>������c>�P>�^>�\�=?<+<��q��F�=�ރ>�2x>~��>��>�K=o�>/���"�п"ł�[4���>u��?e����[����R��}ʾ����g6?v#*>b���Z��m����kB?�ky���B�o����~�i?VN?"Ѫ�ip7�h����*R=v	����s�����ռNo�x+���w>��#?��f>P�u>��3��8���P��e��)}>)6?BҶ��9���u���H�imݾ��L>�߾>�sF�������a ��@i�ţ{= ]:?R�?�޳������u�󁞾nR>ۘ[>�=�ӫ=�	M>A�d���ǽI��+-=��=d�^>m^?v+>�,�=Ɉ�>�U��R�O��M�> �A>�b->�Y@?��$?��0[��ZɁ�\+��w>�V�>v�>�[>-I��U�=�y�>��a>�o�h�s*��3@��>X>g{��k_���y��u=ޘ�h�=9%�=j �?=��'=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿf��>�ѽ㙿#���ȇ��Q->�ژ>�G?�
��7����G�{#�>�c?��
�\j��q�ο�
��ɻ>a��?9�?��s�͛���I6�� �>I��?��#?7j�>��>���H�>�'C?4;d?��k>��.�� u�'�?|9�?�&�?�L2>��? �?���>,�>�N�c��>��1T��-rb�Lh>B��<Ȭ���K���T���fc��4$�~��=.T<cʾ>���>���2�<��Ͻ�O��#����\�>l�H>�3�>��?Z,?SI"?N��>�ז=r�=Up �.v����K?���?�����m�z@�<~k�=��^��?�L4?RsV�D`Ͼd�>��\?���?��Z?���>΋����=�u[���A�<k�J>q5�>KP�>~����L>��Ծ*E�oM�>N�>/��8fھ-��z펻CQ�>�$!?���>��=ڙ ?��#?��j>�(�>AaE��9��Y�E����>բ�>�H?�~?��?�Թ��Z3�����桿��[�p;N>��x?V?qʕ>a�������_kE�)BI�B���]��?�tg?^S�2?=2�?�??a�A?�)f>ч�$ؾg�����>�!?SA��A�=&��3��x?�f?�%�>�됽��ս��ּ1��.n����?	(\?�T&?`���`�0�¾�9�<I���V�4��;yH���>��>�������=!�>Fܰ=i�m��6��b<N7�=H�>���=?m7�=-��.=,?�G�oۃ���=��r�8xD���>�IL>����^?ql=��{�����x��	U�� �?���?Yk�?;��8�h��$=?�?U	?q"�>�J���}޾A���Pw��}x��w�\�>���>�l���I���ٙ���F��X�Ž��C����>���>���>!x�>S��;~>2dj�FI�M�2�5�ܾN7`�T[�_��G������n���<��=7��	�c��k�>���N�>��+?�=�`�>�o?�<{��>��@>�P�>v.�>�]�>+Ҹ>0�~>z|�<{�ǽLLR?6���d�'�5��)����2B?�qd?@3�>t�h�����I��~?ޅ�?s�?@v>�|h�0++��o?�>�>���p
?O:=)q�5�<�U��ҹ��+��V����>:I׽H!:��M�Nof��j
?/?B ��ފ̾�5׽�朾��=�Ɇ?vg&?*y!�K�Q���p��Z�QRW�I��^�m��¦�o9*�s�p�������!��6b*�J�=��%?nÊ?Z��R��������j���;���E>�|�>wچ>!�>'�?>�-���)�7�`�K�(�g�����>�[s?��>��9?G�?��k?p�4?�q>�	d>t&���	>I�>C�>?~�=?�]??Q3R?�?1?�""?��?�i�>�k������P�?]?��?��,?���>���T|��[v���z<z�I���%���="z%=Lr��d���=^��>lY?���ͬ8�]���gk>K�7?���>���>|���,��
�<=�>J�
?�G�>�����{r�ga�mX�>L��?���l�=h�)>H��=����;-Ӻ1\�=�����=����};��%<$��=i�=�:t�ҫ��c��:\�;v�<�t�>5�?���>�C�>�@��/� �b��f�=�Y>9S>|>�Eپ�}���$��v�g��]y>�w�?�z�?׻f=��=��=}���U�����F������<�??J#?)XT?`��?z�=?_j#?е>+�iM���^�������?��(?�(�>���\p�����h	�T�>U�?�.g�9H���$�\���0*�<� <ȵH��>������?��=<>����<��T��?/��?¦���=��+���Q��ްʾH�A?���>s��>:��>JX8�r�^����7z>��?�-P?Q١>�7T?~��? MZ?Hv�>���Я����N+��[�?v�4?�s�?��?9�W?��>!�I=�s=96۾2:)���f���\�t�j��h+>�0�=Uj�>��?Z��>�o3:r��=�!=�0����n>my>��?K�>��>�08>�{�=��O?5��>GѾ&���W����O�B�=3|?u�?OZ#?�=���~j<��g־���>�R�? �?�5?���L�=�T󼪫��}���7�>cS�>%�>��&=�ݑ;0X>Ġ�>���>vO������-�Ӂ��
?&7,?D"�=B9ƿ�Qr���r��ߗ�O?\<3U����`��⓽k�[�ý�=�7�����⪾�{\�-���_̒�+���>��_�z�N�>ij�=3��=���=B<�<�ѵ��<{�D=�Q�<�=�w��!@<�7� 尻�@��Q�_�eiR<@uI=q��~k˾�}?KI?ݣ+?)�C?TYy>x>9�4��m�>�Ā�O#?.�U>bN�:P��RK;�ݥ�����K�ؾSx׾��c�^���n>��G��p>2�2>��=�\�<�S�=/�s=�}�=#�d��j=;�=,��=��=F�=��>[b>�6w?W���
����4Q�]Z罢�:?�8�>�{�=f�ƾk@?��>>�2������jb��-?���?�T�?D�?:ti��d�>X���㎽�q�=<����=2>���=U�2�Y��>��J>���K��H���~4�?��@��??�ዿɢϿ;a/>�7>�">��R���1�R�\�țb��xZ��!?�C;�FF̾:�>��=J*߾Ԍƾ�.=��6>��b=�]��U\���=�
{�n�;=/l=�ى>h�C>��=�,����=��I=o��=��O>C�����7�D,�>�3=5��=��b> &>���>���>,�?�mP?p��>{J"�^�ʾ(�����>y��=7h�>*��<r�=���>%�3?�p9?g;@?dj�>ټ�<36�>2Y]>^CZ��sF�ҿ�=��R�=�]�?�J�?�N>�A&�A:���V$��)��ች��?8F%?�?&�>���P���(H�����sm�pj��O�>q�0��ll�䕛<T��0D��,�.8$>Pw�>,��>�!>U�>�a>�E�>	e>?��<�Uw=P[���=�Y���5��"���N�=��^��;��n;t��<�����YM�q?��>W*�}0��M�=�9�>(>���>Y��=+Ƹ�9�1>\��PM��ۮ=���%�B�Me�;/}��1�� =���=>��\>vix�l'��p?_m_>��=>���?��t?�B>L�DҾ�N���`f��FY��G�=nr>��2���6���]��_M�Ѿ��>�Tg>k,�>�H!>�YE�Kp�3��<.ŀ�F�C�]Ǫ>��O�5hѽ�0<�W��� ���۪�TA��)_>��G?�C��ۃ�<�]t?>�k?���?f� >��8>Q���)M>�㱾����p���>&� ?�
Q?���>氭���b�zH̾*���޷>�@I�,�O���Q�0�4��)ͷ�>������оu$3��g�������B��Lr�p��>(�O?��?i:b��W��3UO����q(���q?�|g?U�>�J?�@?&��z�cr���w�=�n?ĳ�?H=�?>�-�=�*ֽ~��>��?l��?�Y�?��f?ګG�0A�>5�<9�R>������=@@>�U�=��> A?�?. ?�i���������w5��k�<�z�=���>���>S>�(=a/=N#�=oqD>���>��>"�a>$D�>X�>�ҫ�?��ӟ@?J��=���>�}#?��m>A r>q�����+�\�.�R����6���ĽÓ�\�;A�=��>>�&=`J�>TRĿ�?���>7����N
?�HǾS$�=r7��bl�>�|���}>�g�>fNr<tW�>8��>5�3>�XB>1�0>�@Ӿ�>o���j!��6C��yR�g�Ѿ7tz>�����;&�]�������:I��y��"k�@j�!2���>=���<F�?����r�k�o�)����˜?�6�>�6?/⌾>���>���>mݍ>�P��閕��ˍ��Wᾟ�?���?)9c>��>��W?f�?��1��3��tZ�B�u�(A�l	e�Z�`��፿����2�
������_?E�x?yA?Ik�<�2z>r��?��%��ԏ��+�>$/�<';�G<=?0�>�,��M�`��Ӿ\�þ+3�SOF>A�o?%�?X?RV���:�Ķ=�,!?�+?�C}?��1?�@?�փ��?.2v>	?��?�I?�<?L?��\>�0>��==u6��"7\�#'X�D�D������Q�/8
=4�=Ȯ=�l�=�p=j�ɽ�ǭ� ]�X��J�����"=��<���>�]?�u�>���>%E7?����:8�����C/?iG?=ɀ��߈�C�������P>�j?H�?AZ?�O^>�YA�<E�U�>�֊>T�'>�^>���>���qJ� ��=�>�>B�=Z{N�O���	��ɒ�w6�<	�!>���>�.|>	����'>�{��20z�A�d>a�Q��̺��S��G��1���v��X�>�K?��?V��=�^��*���Hf�0)?�]<?OM?��?��=��۾��9�E�J��<�	�>B\�<���0����#����:��<�:��s>�1��%u����b>1���߾=�n�6J��:羬�W=�@���N=s_�K־>����=\�
>W"���!��,���Ȫ�d2J?�"l=���}(V�*���>}V�>w�>�:�Het�@����݇�={��>";;>J吼��ZG�c$��֖>�d0?��\?��??$��[���G�'�����t��>��?LU�>�\-?֔�>!��=��t�������Q�
=F�'��>�S�>����6�=)ܾ���O9���=�4?p$�>�r?&�Q?U?e??3?1,?"Z>$��H��`�*?p��?Ʊ�=�et��A$��M6�:b���>��+?��<d�>ý(?T^2?�'?DZ?��?D0>���_�;�_�>�d�>�,>��%�����>��G?z�>��M?!�?G��r�#���+��3?�&0�<�&">��,? �&?�E6?
�>%a?�̾y����_�>�c�?l<�?K�6?І4>��L?���>*�G?YG�>���>yW?>J?�i@?rWa?��]?(A�>���:��*£��"�=Dv�nл���=�x�=+E���iy=v7����Wê�Q�/�����x?���i��VG�E!�=-_�>T�s>r	����0>{�ľP��*�@>E���Q��sي�f�:��ݷ=�>��?S��>�Y#�n��=���>|H�>����6(?��?@?�|!;]�b�m�ھ��K���>�	B?���=��l����|�u��h=E�m?H�^?S�W��&��N�b?��]?<h��=��þ|�b����d�O?<�
?0�G���>��~?f�q?T��>�e�*:n�)��Db� �j�&Ѷ=Zr�>LX�Q�d��?�>n�7?�N�>.�b>0%�=gu۾�w��q��h?��?�?���?+*>��n�Y4࿹�þݖ����e?W��>�ƾd�?��=�E������S����þ�kA�?�ɾ(U-�W"�%���{���o=��?�p?��g?� h?]gj��R��6t��O��=�d�ɫ�����Z��W���9���r���]x��㫾1һZ�w��C�K��?Y'?��4�X�>j������)о��I>�4���b��[�=␽((a=�[=��_�Bf+��z���<?�|�>���>G^>?��X�
g;��s0�ƛ8�ϑ��~A>궢>D�>X*�>�����'�%j���ɾ���u�Խvy�>%�j?y�U?��Z?EZ��+�/����.�3�;Z���{��p=�ϐ=:b�>E&��$f�N:���'�&�^�8�����/��@1���F:?�M�><��>�(�?�?��ܾ�����4N�����m	=56�>e�r?8*?�~�>����0������>��l?���>��>�����Z!��{���ʽ	$�>�߭>���>��o>S�,��#\��j��E���V9��t�=�h?���0�`����>R?�[�:+�G<E~�>��v���!�b���'���>}?Q��=%�;>�|ž�#���{��7��QN)?+?��a�)�Z=�>*C"?z�>���>!'�?mߛ>J����F;��?*�^?aJ?�gA?�J�>uX%=���@ȽR1'��(=��>�g[>��r=���=S�+*\��� ��H=Г�=R�ͼ)���jT<�Ƹ���;<���<��3>ڧ쿼�[�J�辝�.�#V征:��@��c&�=����0B��|Ծ_��%��+��5<��5�ãM��	����m��1�?�I�?�|���
ܾgѝ��~����#V�>iw2�:������A��놾r6��r��c�������Ɣ��.z� ��>��㽇	ֿKe��h�1�u`�>EL)?�i?5k��$c��E���Q��*�����Qb"���ڸֿe5�spS?k�>;��6�<=��?c�<QOt>��#=9���{Q¾,�>��P?Z�2?į&?oyf��fݿ������=L��?��@|A?��(���쾳?V=���>��	?��?>�Q1�J�6����S�>E;�?m��?S�M=��W���	�de?�<��F�$�ݻ��=;�=�W=���ǑJ>�Q�>���:OA��ܽ��4>�܅>�W"�����~^�8g�<��]>��ս9;��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=@��1ο�1"�D%�6�<�/˻X��U�\�����%����Yހ�Jj1���=��>�Gc>7��>�"e>�	d>!!M?1�n?��>��d=���Q���;i<显r�\�����1�Nl��V���v̾�����)��#(��hξڛa��=�2X��y����&��b�=�@��P?�"6>�9��eq��f�?k���oھ�+=�Y��u��D�^�� v��&�?z�[?u�����]��95��$_�>�=�W?�/�����־�A>��/=%+���Ֆ>1�i>���mpl��w`��q0?�V?�[��}5���T*>j� ��=ѿ+?ny?��\<!"�>�J%?¹*���㽇][>��3>+�>���>��>��/e۽�?Q�T?H���眾�А>5V����z��Yb=3�>5�p����[>9~�<Q���Q�R��P���@�<�(W?s��>��)��va��]��,Y==��x?��?$.�>o{k?��B?�դ< h��|�S���bw=�W?2*i?��>����	о^���D�5?�e?��N>�bh���=�.�]U��$?�n?5_?\~��(w}����n���n6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>�������>������?ܣ�?b|����������[�k�����x�<�I8������b	�f�$�y�پ[��/����*a�0�C>O@y��_��>j7m�D�ٿY��u������eu��a?�Cl>?����"���+����w��N�$�;�3]�����>�>m?�� ����v��:��L��m�>գR�s�>�\��㾾���^�;�	�>���>6�~>\ݶ�?4���ɕ?�%�n+˿Ƌ��1���Y_?� �?~t�?r�+?�;	�[&Q�\�����U�I?�_t?��Z?���I�F�����l#`?�����W����t�S��w�=�_6?��>��>���%<F�>�P?�R>>�8�v4п������ٝ?_�?}Z����>���?LQ5?��Al��4Z��B'��z���S8?+�e=Bݘ��#��@������� ?h3?Y:߽W+�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?C$�>��?��=�e�>�q�=ﰾ�_-�Wk#>��=
�>�[�?�M?lM�>*g�=��8�~/�gWF��ER�m%�,�C���>,�a?��L?.;b>�!���=2��!��iͽ�E1���TM@�g,�t�߽�(5>��=>>8�D��	Ӿ��?Lp�8�ؿ�i��.p'��54?0��>�?����t�����;_?Uz�>�6�,���%���B�_��?�G�?=�?��׾�Q̼�><�>�I�>9�Խ}���^�����7>/�B?J��D��s�o�v�>���?
�@�ծ?gi��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?mQo���i�B>��?"������L��f?�
@u@a�^?*��Dh���4���־��=��=F��=/��=��(>�ف={�;%R���ˆ�Q��>�)Z>t!�>3��>FF�>�>�^��������Bx��}�9�4� �~��������^�� ��J���Tܾq��[�=6���I��Ѓ>�⣐�R�>>�N?�:R?��n?Wp?ȼ�����=��Q<9�	�TF	=i�>��/?_�H?AV!?�+�=�����zZ��7�_���ƒ�&�>�j>�Q�>6b�>�m�>�*0=�
>wh[>�A�>�>�_=uP&=��=a"D>��>���>s:�>tܽ�ڷ>K�¿�~Ͽg:u��vݾ��>g��?mS���������mϿ�(� ��c%�̏+?� �>쯣�f��H׫�:�B?���:1��T>��=�?��Z?!�h�0��������=�l����g��-�=FU�)n�j�"�*K�>&�	?�b>~y>6%5�i9��Q��l��7��>�,5?K�����@�z�v�X�I�ݙ߾yG>�>�>��[�� �1K����r?f�6Br=ɯ9?.�?P��{(���s�sV����O>r�Z>IK=K�=uML>�w�I�ѽXJQ�6%(=^��=Jc>�"?1�+>�q�=?��>�L��"�O��ħ>S8B>�&>7@?&�$?˱�v��T���>-�J+v>$��>>+�>i>�I��8�=��>��b>�-����`
��A�иX>��T�V�W���h�`#�=�����=�ϑ=]���B�>�ϗ#=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ��>���̕���k����v�=�=���>��F?G����]�� <�_f	?�e?i��;H��X9ɿ�w���>t�?Å�?7cm�Yt���>����>@��?��X?	�o>6�ܾ��R��>��A?c�R?�:�>~��'�*���?���?�K�?�Z>�8�?� �?�R�>k?��r(��[ο:A����;�=�9D=$�:�y��n_b�����N}��l�Q�8��"��q�=��>^���|��v�=!ؽ�}������S�>�Y9>������>�
6?V�?���=�=�=f� >��2�����|�K?���?$��G1n��f�<���=�^��$?�I4?[���Ͼ٨>ۺ\??�[?:f�>=���<��~翿d}��E��<�K>n1�>�J�>����HK>o�Ծ5.D�ti�>gЗ>ǣ�Bھ-��u���GB�>g!?>��>Dծ=�� ?��#?z�j>�(�>4aE��9��;�E����>���>�H?��~?��?�Թ�Z3�����桿��[�`;N>��x?V?sʕ>Z��������lE�7@I�e���f��?�tg?�S�:?02�?܉??`�A?�)f>w��ؾ����>[�!?q���A�;N&����|?DP?���>$0��v�ս"Fּ���8�����?l'\?�>&?x���)a���¾�F�<�#�y�V�,��;vE���>�>^r��[��=L>Iݰ=�Hm�T96���f<p�=��>w�=V*7�&w��0=,?̿G�~ۃ���=��r�?xD���>�IL>����^?kl=��{�����x��	U� �? ��?Zk�?b��@�h��$=?�?S	?m"�>�J���}޾6�྿Pw�~x��w�Y�>���>(�l���K���ڙ���F��_�Ž`ZM�0��>s��>L�>�]�>�i	>�>���z�fԾ���?�g�f�/�>�$�߯����QJ����:z����M�1�g�J>A!��\�>W�!?��%>J�>!,#?�f\����>d�?>�Rk>�ý>L�>͑�>��>;�=�=��KR?����"�'���辽���g3B?�qd?S1�>gi�;��������?���?Ts�?=v>h��,+��n?�>�>G��Uq
?kT:=�8�';�<V��{��3���1��>E׽� :��M�Cnf�vj
?�/?����̾�;׽�<����=\0�?%-)?��#�M�M��w�Y�Q��rZ����gY�0���
">��t������U������*D#�-/�<{�?z4�?p�پA���#y����g�,\��.>�+�>Y=�>���>��4>#���b/��+a��$��4���H�>��f?ݫ�>p�L?��<?`j=?�O?uS�>a(o=�W�l5?[D�=��>8z0?kC&?�+?��?U�2?�X?��>���u�Ѿ B���>��?2�?Z^?�E*?�m_�=�C�,����L=��M�#͟���3>-
������=���=��b>�X?T��j�8�e���lk>��7?��>���>;���,��g�<7�>ϵ
?�G�>�  �)}r�Qb�W�>M��?)��܁=:�)>���=9�����Һ)Z�=���g�=�.�� v;��p<���=��=�Lt�����`�:���;�w�<�t�>6�?���>�C�>�@��.� �_��f�=�Y><S>w>�Eپ�}���$��p�g��]y>�w�?�z�?��f=��=ܖ�=}���U�����>�����<��?DJ#?&XT?^��?z�=?dj#?Ե>+�dM���^�������?U�? �c>;�%�NP���/����+�@"?�`�>J�u���K�y�!�����=|bE�>�z�Q���U��C!$�k��>m�e�ܽ��?�}�?Y�>�|�R�g@���B�0BԾ�8D?:�>�?���>"��"Z�|h�彫>c?�qU?Yr�>��V?�;y?�'P?&�[>�4������:��ߨ�<9�N>w�4?�E?�2�?��o?���>�]7>�� ��o̾L ����]��?�|�VB=�}�>Xˠ>r��>f}�>��>�#���������=��d>G6�>܋�>@�>U��>��)=o�G?�H�>�达�|�������c�B��Gu?��?��+?6-=�d�E�����Y��>qg�?��?�:*?6�S�[�=�ռ�n���q��x�>�:�>�i�>�k�=ʚI=t�>��>[��>\!�aT�{8�qQL�K>?�?F?��=s�ſHq��p�����`<���
wd������rZ����=�������A����[�Wz�����������]����{�۸�>D��=-��=�[�=e��<��ļށ�<�Q=��<�=GJn�y~u<��2���ɻ~������ŋh<��J=P|���:˾�d}?9:I?��+?i�C?�ly>`�>T}2�u)�>H�-?GV>�5O��$��+W;�m���Ҕ��ؾ�׾��c��ן��>�"G���>�t3>'<�=�2�<�0�=bDv=���=XS/�9x=.c�=���=ca�=c��=��>`>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>	�3>/�>>�Q�2�1���\��"c��SW�x!?Ѷ9�c�ʾ�T�>�E�=	hᾱ�ž�1=)�1>��W=���[��ӛ=~���M�1=�O=
ԃ>j�E>�9�=�Н���=��K=A��=ƾQ>��r;y23���!���F=��=�7c> �#>"�>�'?�0?A�c?U��>�{��ݾ��̾��>'$>@��>�E�=��i>`+�>��8?�yE?ץI?I��>�I=>��>*D�>�%*���o�.tݾ�������?#+�?�:�>�w#<�6 �9����=������?�-?ϝ
?�V�>V����Y&���.������"8��
+=�ir��RU�<���Gm����|�=`p�>��>(�>lVy>��9>_�N>.�>x�>�&�<h�=�&����<p	�����=(���h�<��żV���i&���+�
���#��;)�;9Q]<Dn�;���=P��>1<>��>xX�=p}���3>ۤ���qM�"��=v꨾'�B�KQd���|�)�-���:��)>>��S>�v���u��.y?�T>E�+>a��?��w?N>���+�Ⱦ����W���W�%�=�g>tb1��8�>�^���J�d7־���>޷>��>�?�>
�H�)����h|>�P��f}�=m�>�:ؾ��ܼHj���~�a���߭���T�d����a?,�|�B�>v�f?���>,\�?-�?�������	��>�A����Q��ξ�B>N�w?BW[?�$�>�;��}��bT̾ˌ��ȷ>�TI�N�O������}0��j�f߷�=z�>����Ѿ�63��U��䏿I�B��hr�ͺ>��O?Ӯ?��a�[M����O����N���I?�g?3Ԡ>�?Q]?�O��s����w�=�n?t��?:-�?U
>�~�=����(��>��?R��?���?�s?H�>����>bt�;#>���.��==s>�[�=�c�=io?X�
?�i
?2F����	��\�<��@}]����<�=�ϒ>�Y�>(�q>;��=��`=�v�=�$]>Ţ�>-�>�Zd> �>S��>����%���?lx��oS;��?�>�ő>��[��C�=��~��0s��;�_��{�;=h9�:��<*B�=]@K�I��>�Ϳ�B�?�h�>P�-��?K���� ;��׼$5V>�-ѽ���>�5�>Hv�����>�p�>�P>��h>@U>>R&Ӿ�>��V�!��#D��mR�@z;wu>�e���/��A
���EO�I��d��j�m傿�1>��X�<�ڏ?Gi��|j� �&����R�?p��>l�3?Hm���z��V�>���>-��>�������p��G�߾
L�?F�?�gb>��>��W?@q?�t1��3�Z�d�u�T9A���d�G�`��㍿Z����
������[_?��x?I1A?��<��y>ٝ�?��%��𐾀��>�^.��.;�>�C=���>�����_���Ӿ:$ľ+���AG>̔o?��?�l?rW����=�]�=n�?��&?b}?�"D?�? ?L@?�nK?�R�=L�?#�,?J<?^�@?MD�>�Î>J��>��=�DU<zѫ��Ț��5�Ù���¼��=#�=R�>����؄D=E>ck�nO��=k
��ŭ��)>��=1&�=�N�>[y^?�`�>/��>H�7?q��@:��԰���0?��N=�!x��3}�la��=V��]	>��k?�ޫ?�`Z?O]>��A�~ZD�%�>�(�>*.>�g>�Ͷ>̾�ˬA�Lb=_e>��>��=rE�<��-��Lg����=��!>���>�|>�ۍ���'>~���)z��d>�Q��׺�-�S�y�G���1��~v�MJ�>��K?��?��=�\龕5��	Ff�=8)?�\<?MM?h�?i�=��۾��9��J�TH��>Q��<}	�����$��2�:�:�s>t1���|����b>C��h�޾��n�J��[�O=�9�y�Q=�a���վ��~�'�='�
> [���!�^#���媿Q&J?�1k=�����U��s��W�>��>6��>&7<���y��a@�u笾p�=%H�>�:>�蚼�ﾴ}G�J6�P`�>��I?��d?�j�?{zh�\�Q��P%���ƾ"��<�>tt�>���>>�?,?>��j>X��Le׾��M�d�;1�>�e?4C��7��gɽ�g�=�'��� >���>�X^<�Q�>gт?{�,?�:�?6�?y�!?�u�>O�׽�̾�C+?ԭ�?���=��L��"#��T7���F�;_�>�B?���V�>ܒ/?+s.?�F2?%mW?��!?�O>R7�QAH�z�>&��>�J�����te>�F?�d�>7N?��?-.>�z�Bՙ�I怽^<>�(>&�!?4L-?�)?Q}�>�/?�z�H}�=J�>��v?��?�wx?����"?�>�=y�(?��i>w�(>�$??
A'?I�t?�=~?��K?^��>� J=ɗC��L��21ȼ����=w�8>��>���=��=�O�=�m�����b��`�^�K��zv��-;�v�;PZ�>��p>z����./>�cƾV���?>l���
��6����:��ķ=�'�>:�?�,�>\�%�� �=���>+��>H�n[&?9?6�?�{�;�a��"۾�N�ט�>��A?�=�=?�k�o���t��i=5�m?�c^?�U�o���J�b?��]?h��=���þ��b�ɉ�[�O?8�
?��G���>��~?]�q?7��>
�e� :n�!���Cb���j�BѶ=Ur�>BX�7�d�k?�>b�7?�N�>N�b>�$�=Cu۾�w��q��m?��?�?���?�**>u�n�T4����ř���R?��>�\��f?��=c���^���YP@�������ϾIgC�9����؞�]j��|E������=G�?Ć?�Q}?�mX?e���ml^�<nd�C-��/i�,r����(K�͒N��W��3���.��"�����FX�=)~��]A�1i�?�(?�/��7�>Ǚ��u+��̾E>u?��'����=�!��|�B=.�\=��g���-��]����?1G�>�r�>�<?6~[�J�=�'�0��u7�����3>-�>�h�>��>�(�:2�+����Tɾ
ℾµսj�>�VM?U�??=]q?M�����)��ʊ�Y~��=��a�4b�=�4:=��>y�u�`�q�j�"�jK+�8M��d���VN�Iz��l=8oI?k߃=���>(Ҡ?W�"?�5�Xd�y�/��>Pp�>�l�?�M?x�9>��w��^(���>�/b?�c�>��>?����_A��?s�@�>y�>0�>G�g>W�w��b^����U����&��/�=�h?>�E���x��9>��a?�-��,��$��>P��=�����ھ0a����=6�?�'8>�f6>գ����f�q���,N)?��?����)��b�>#�"?~��>��>_A�?�ޛ>q������:mi?O�_?�{J?a�A?���>�'>=Rp���1ȽTx(�*9"=�4�>�^>�x=֦�=Y����Y�r"���@=V!�=U'��Ʒ����;�X��L�1<�$�<��5>3mۿ�BK�i�پ�
�#�m?
��爾%���d������a��F��Xx����'�\V�:7c������l����?�=�?〔�V0�����4����������>��q�E�����Q��q)���ྋ���nd!���O��&i�k�e�V�?>�A�c�̿�h����i�?N*?���?����+��I�Қl��Fv9ŷ��n��s��5�ǿ_@�xQ?��?}<��Z�=UW�>�r>^μ;	�=�έ�/h���>>?��G?^ �>mܽD��A?���z=>���?�/�?�@A?�))��f�9R=)�>��?\?>S/�^m�֤����>w�?`��?w�P=5�W��D�0�d?��;t�F����b��=z�=�� =b�
��XK>�q�>�!�B@���ڽ]�5>�ȅ>#�U���^�H��<o^>="ս�[��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�򉤻{���&V�}��=[��>c�>,������O��I��U��=L��wѿ���ld��%�=�-���<�ܞ��	ܽ_��=�"y�":L�2F�=$�E="�>Ny>�"�>�ED>E<�>$sM?7�Z?&��>.a�>{��3������@��n5���E)�i�h��������F/�����Q���#O��Y�Ȫ߾f�u�8�>P W�;����A�!"���'��2?1��>�S����x��-�<��������y�=�T5�����{G�Ε~�3R?��%?�S��Lx�/>�����޳���8?��ս-��	
��R�<�������P��>�q�=/5�Dc�n��s0?8?y���g����)>�� ��7=8�+?�w?vˇ<�Ъ>i�$?�A)�P[彲K[>��3>#G�>���>>ј���ٽu�?<DT?���딜��.�>�����|�#�f=S	>�t5��l���tZ>Bת<���"T�[���Ȯ�<v(W?ٚ�>��)�	��a�����X==��x?`�?�-�>/{k?��B?Ԥ<�g��{�S����`w=��W?�)i?p�>0����оw�����5?��e?z�N>hdh������.�U��$?��n?D_?,���v}�J��?��|n6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������n��=H�����?�P�?��|�Z~�����c�`8#�8�1;ax�=�A�}$�<����b@�k}վ��
���
?^=&�>��@6�a�U�>��m�G#ֿ�ٿ���F뾺^���Y?�ʜ>͑����Ӿ�)���R��b�`�h�7����X�>�>g��r�����{�k;��{��H�>�c��'�>��S��4���j���3<0Ӓ>���>o��>�஽߽�C��?>W��u.ο&��������X?�o�?�p�?dZ?_�@<?}v��{�,m�� G?ޟs?�%Z?i�%�s"]��8��j?�a��#W`�?�4��KE��U>� 3?�N�>�-���|=�>)��>�a>� /�ԌĿsٶ����U��?i��?}i�A��>T��?�w+?�b�7���c��Q�*���'�p<A?2>Ȁ��¶!�8)=��Ғ���
?�0?'l�0�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?%�>G�?�q�=�c�>dU�=`�N'-��q#>��=~�>�N�?�M?|H�>O�=��8�!/�QYF��ER��$�o�C�V�>��a?5�L?rPb>����2��!�A|ͽ�d1�7M�~S@�ߦ,��߽�,5>d�=>�>&�D��Ӿ��?�`��}ؿ�e��'�*��43?Q��>��?M3�*u�H (��^?"�>�������+=��
/�%�?	��?u�?W�پ�k��l�>��>���>Z۽�~��e���19>}�B?~�����n��M�>3��?��@���?2i��	?���P��Ra~�#���7�Q��=��7?�0��z>���>�=�nv�ӻ��U�s����>�B�?�{�?	��>�l?��o�8�B���1=^M�>k?�s?|mo�x�{�B>��?�������K��f?�
@zu@Y�^?(J����}�����ጾ��}=�4S=�`�>���;m,>�A6=����d1�<j>B��>V��>��>�'4>�q>�� >D���å�5����v���q�tUG�Ͱ�2aE�I��L����K������@��:���ȼ;l��$sӾ�t���vM�b��=��U?�R?R-p?�~ ?ֹ}�b�>H���k =$�!��E�=�>��2?�L?��*?��=���Y�d�<���%������=��>�mG>Q��>YL�>�>���:�]J>Ԡ=>� �>mL>�D0=T<;ߩ=�dO>�>�>zn�>V��>�8�b*y>�3Ŀ����������X�+��=�͕?�C��߄��᧿�S��zz����G�@�&?I~>f���J6ڿ�_��/�Z?;,i��+,������I >�~V?�1?�3>�����%����>����
�o�acp�a8��ԥо~���I>U�3?-h>6�a>7�}:���T��h��$�{>I�<?�c���)=�j3s�'�C��ھ=L>��>rF#����̕����w�p�\�\mu<
�<?�
?�z��鴾6*��6٥� �Q>~�e>�Iq=1�=y�H>{�w[ҽ��:�Y΅=�E>��E>�t?�n4>�M>��?���.eM��OV>6�>&��=��g?/v?eZV�Ĥr������B��\>�>M[�>񛶻d3�
�1>��?ڍM>����Y�@"�=������w<e���+����*{��T�����>P	%>��M��,y�yg���~?���(䈿��e���lD?S+?_ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��J��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ*��>N������A��X%x�M��<�8�>њL?�����^c��hC�c�?�?��ۣ����ȿ�4u��-�>�"�?Jٓ?�:r��H��p8��a�>mb�?��Q?~�\>�e׾28N����>��B?ŏO?��>����"�%?�7�?�j�?�3�=gM�?3"p?r�>ͬ�=N�ʿ�'���^>�X��ʮ>ڸ�=��G��v�F�����/QM��3�����>%��=?��>�T�D0��>"�=?ݢ=R�þ�z?���?P�l>��Ǹ>�� ?>��>po>ý>V��=.PK��$q���K?���?���.2n�/U�<��= �^��&?4I4?�a[��Ͼר>%�\?q?�[? e�>���>��H迿�}�����<��K>63�>�H�>�%��AEK>-�Ծ�3D��o�>qЗ>��>ھ:+���C��,B�>�e!?I��>�Ԯ=�� ?��#?'�j>>&�>r[E��8����E����>Ƣ�>�E?j�~??�?ٹ��[3�X	���桿*�[�">N>��x?�T?�Ǖ>H������.�E��HI� ��?�sg?�5��?�/�?{�??-�A?/<f>xv��ؾ-���f�>#�!?����A�2&�5�ee?.=?7��>zœ���ս"�ռ+��Sp��x�?�\?B&&?J��|a��	þ��<�;%���D�ko<��9���>-�>鏉�	}�=��>��=?m��?6��(i<{��=٤�>��=,17�ԭ��0=,?��G�xۃ���=��r�>xD���>�IL>����^?fl=��{�����x��	U�� �?���?Yk�?n��>�h��$=?�?R	?k"�>�J���}޾4���Pw�~x��w�^�>���>
�l���I���ؙ���F��k�ŽE�$�;��>`L�>Z�
?Uv�>]�P>�>�_��'�*��� �I�[����M}5��-��E�I�����������x���>����"��>U�?t�n>�-�>5��>��$��@�>3X>Ti�>��>�_e>�8>`|
>\f<�鸽�R?:x��#�'��辻����bA?�d?v��>�o��R����-e?�9�?�<�?s[t>Y�h���*�?���>>���]	?ё@=`A�����<[䶾�D�<��rH��̎>%sӽ39���L�&ad�$
?�r?�����˾:�ڽ6����B=���?+�$?p���U��&n�d�k��&{�ڋ��2���ž�f<����������������0�A�X>��?�ɕ?�������贾��Z��,\�*>k�?Z5[>{m�>>YW>'�;��7�gQ�X=�ʹ��~�>��[?�h�>3\?a}E?ӡ:?��G?UK�>dx>:D��`�?C�=!��>%�?V]>?j�S?��F?`�(?j�U?2�?����)߾TRؾ�0�>��>�-&?��0?=l?T�߾�sy=<bԽ|�=�ɬ��bp�x��=��}�o�нDw����>c�>��?�����8�I����>j>��6?l��>�?�>�~��━����<d�>ԃ	?��>�4 ���q�����	�>LL�?�����=�+> �=Ozb���a����=�����1�=�G���9A��y9<��=��=�c8b�T��׌;{��;���<�t�>.�?Ǔ�>�C�>z@��&� �~��ee�=�Y>TS>'>�Eپ�}���$��~�g�X]y>�w�?�z�?$�f=��=���=�|��0U�����S������<�?J#?XT?M��?R�=?cj#?��>�*�QM���^�������?X+?'��>�����;+L���4�^1?z?��a��?0)��1��߄ֽ�4>/G/��~�}@���RC��3�����n��2:�?H;�?V$��7��R쾩1���w��B�C?G��>,��>�G�>xF&�$�f����^�C>���>M�N?�>�JW?E�y?�[[?:Vl>�8����Dލ�iF�c�1>��8?ԋ?/��?��}?���>\s>�ַ�F	ξ����I޼��xy��p��&d>�5�>T'�>�$�>��>�̽Q����2��=͠>�o�>�ŕ>}��>#o�>�=�=��G?���>AN�����c夾A����*=���u?a��?��+?܍=1z�q�E��5���Q�>�m�?���?.7*?<�S���=u�ּ�ڶ�S�q���>i�>,=�>��=v�F=�b>�>��>�;��\��i8�]M�;�?)F?ϻ=T���9��]6��H�W��j<b&a�d ����򭛾x��<!b�����J����k��Cѡ��(��Ԑ��6����>m�=�@>�4�=@�(>��4=k?>">+�==g<�?���O ��T�0��l�s<�_�;{ =�
�=X�>>�ʾ�O}?U@I?�+?}YC?
y>?�>ת.�5�>�+}�-?_|T>�AR�ﻼ�ws:�n��+}Yؾؘ׾�c������>��H�E�>��2>���=[I�<a��=&�o=�ȍ=e6��L=��=Yb�=0��=��=��>�h>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>~�/>��=eXT���*�X�f��^e�B$V�k?(�;�.�ž0�>���=�ܾȵ���z<�v >a]K=����{X��a=�����%�=�Z�=�W�>Y�Z>��=��Е�=4�:=�4�=��;>�wӻ������=�Y�=��W>pH >2��>�%?f0?a�e?�Q�>�ym�_�оa���O��>��=��>F�x=��O>o�>�y6?3aC?�=I?.ߴ>��r=�S�>Lx�>�'��ki����j�����;=��?�ǃ?x�><�<+_F�:����;�7���?�;/??PR�>��	�M�ΐ�$�"�)��WU��˜��6{=��L���Y��P�<��	��%��م>�B�>x4�>��>�M�>';>#�u>��>��=k�=Ly�="�=�Ҝ;-?�;�m={�憡=p����9����n=T74�w�;3(=�9(=�};ad�;���=���>5A>i��>ay�=����>/>����o�L��߿=_C��K+B��1d�KF~�/�'Q6�p�B>Y4X>�����1��e�?V�Y>�p?>��?�=u?�>|.���վ�O���Fe�DES�ϸ=��>�<�Rr;�!U`��M��~Ҿ���>�>�0�>F�_>N�.��R@�'n=�gվ�m6��p�>���qX ��|�^�l�s^��º��Bnf�Hj�$JA?a\���l�=�}?��L?�?�)�>3������WN3>��z���E=���n���m��T?NR)?{H�>H��A�E��0˾gM��e@�>�0L��P�������/���M�V	���]�>�f��+оz�2�����"Ώ��C��Os���>W}O?���?��h�x��^M�Ը������?�?f?��>�u?��?�E���쾅�|��V�=Dn?���?��?2�>e�=�wؽ7�>�?/��?ڈ�?�sq?;j0�w��>�l�9�!>32��tp�=Y>6�=��=�?}}
?�?�����>�K���I��PQ��ӭ<�T�=���>��>��>��=B,�=ne�=L�M>ý�>Sؕ>(�r>}��>�~�>^ۭ���3����>�jV��#>XH�>��>�y>H���OU=E���g�G���潓/��ބ��!��OHC=ЈY=�=��>�Zÿ���?
�>ր�Vi�>��~�V�ds>;/�>:xP<xx�>6�>e
�>Ix�>_��>+��>ŧw>��=��Ӿ�=>
��D4#�5FD�ѻP���ξ�m~>�����z*�ك	��_��H�����g�şi�Em���>����<�$�?eE��i���(�$��	?��>�m6?&掾B|���>W��>���>�V��C|������V�ݾ�?=��?Cc>��>��W?Z�?��1�!3��rZ�f�u�'A�R�d�θ`�n���i�����
�c��_?��x?uA?�ّ<:z>â�?��%��͏�,�>x/�`";��<=&�>�+���`�3�Ӿ]�þ(��OF>ڗo?z#�?	T?dV�~@̼$($>%�6?��-?�v?d.@?<9?�g3�r�"?r
�=rq
?�?�D1?b7?�O?D*Y>��>�\�:3R�<>`u�x���'v�sŽDMs�z�.=7�f=I���;���"�=�1X<���-}?������Ƽ��]�!r;=���=Wԇ=���>�8^?'��>���>9?�7��!6�N괾�p1?��>= rm��u���|���m߾��>}�k?,<�?�b?��n>��@���K��>\o�>>4=>'Ji>$Ӵ>�I�:�7��p@=�q>�>S�=6O;��^��m�W2��p��<};+>���>�|>1���'>p����8z�K�d>�Q�HѺ�V�S���G���1�҃v��Y�>��K?u�?���=�]�y>��7Ff��')?�]<?�QM?>�?[$�=��۾��9���J��7�q�>$Z�<������h ���:����:ɺs>|5������?�a>���"߾��n�J�I�%�ƥ_=x��zK=���־������=_�>�!���y �K$���ت�'J?xVr=��� X�pW���F>_��>J�>��<����=m@��1����=���>��<>A����uﾩ�G�x����>xMS?�[k?�?U���"�l�1�ߓ�Bʠ�9��=Dc?P�G>��+?Rz�>�F>��j��8�i�G��b�lt�>�^�>������@�)���پ\�-�=by=?&��=��#?�n�?F��>f�K?E5?I��>ۜ�>�$4�(�`��q'?*��?���=��@�M�l9���F���>�)?�;�[D�>�~?X� ?�'(?*�S?�?��>����|�@�[��>?�>wxU�i㯿j�e>щI?�.�>i(V?�/�??@>��/� ���r2���y >zp>g5?:,?��?d�>3�(?�B��M�?�I�>�J�?D�?YM�?�=��/?'�D�z�?P�>�� >0�H?�<<?�r?�ӎ?��?`��>"��=j+�~�"��&���;�d=��>2�:>5a�<���<q"r�e&=��V=�B�v����`��z��6�>=�_�>��s>�	����0>A�ľ�P����@>����oP���؊��:��۷=���>�?r��>�X#����=���>I�>��C6(?��?�?4i";��b���ھ�K���>�B?���=��l�7�����u��h=��m?@�^?D�W�!'��O�b?��]?>h��=��þ|�b����e�O?=�
?-�G���>��~?e�q?R��>�e�*:n�)��Db���j�%Ѷ=[r�>KX�Q�d��?�>n�7?�N�>1�b>%�=hu۾�w��q��h?��?�?���?+*>��n�Y4��� 1����_?I6�>=ޓ�Y�?V��<ϴ��u����H�G���
&ľ�����ڰ�.���w]�x��>%߽#d>=?"��?;k?��~?�Ͼ�U����S��f�/JQ����_:�ܬD�>�6�J[g�f0i�Z��2$�����Ӽ�‾z�C��ִ?;q%?��.����>�w��J%��q;m�G>c����X��7�=�u��*@=�<U=�d�c*����?�i�>��><M>?�JZ�4F=��O1�w�4����O7>���>ik�>��>�7���)�_@ܽ�a;$_����ֽA�>7l?� =?�t?>*���5��{���M�Z��mȽ ��>I�3�J��>�8���^5�t�侗!���O�?>���B���s(�=��U?zB�=/>-�?�j&?�7&�=!S�	���F��kR>'a�>��W?q�?�QK>S,<l�0���>��m?�z�>���>Nň�'� �� ~�彈��>�E�>K"�>��n>P.�ܻ[�F��0E��e8�4��=��f?U�����_�M�>a�R?��!�:�A<Y�>~[B��N#�U����� >ި?�u�=<_D> Ŀ�5,��Vz�����)R)?�J?6ݒ�Ę*��G~>�$"?"��>�#�>�0�?l%�>hVþ��#�c�?>�^?�CJ?YA?p_�>c,=2����;Ƚ��&���,=%��>L�Z>19m=g��=Y���a\��|�s�D=O�=�kμ�7���4<q���=L< �<4>��ۿ�%L�C��*�������T�zR���?����q�Pg�e��񋕾�u��9��(��j\�V�U�Q[��"Wp�Ƀ�?c?�?? ���t��.ɕ��~�����>��[������YþD�!��I�����
2��|�ĪP��ds���e��??WK���ſ�勵�f��8.?�|(?�|?2����4�^��š�jA>�����龠���lп<\ʾe�C?i��>����E>$ �>�Z>�,��'=N���d���J\>�(!?��O?�3?X��>�޿��Ŀ�D;�G�?G�
@}A?�(����tV=F��>!�	?�?>�S1��I������T�>s<�?���?�|M=t�W���	�9�e?`�<��F���ݻ��=�;�=bE=u���J>zU�>���SA�?ܽA�4>Gڅ>�~"�X��܂^�Ã�<ȇ]>��ս;��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=^���!ĿM2�k:���g�L��<���~ʍ�k��<9�=�$�����>��#���>���>[-�>T�>��Q?��r?��>�F�=�p�{�-�\񺾜ʆ>KQ������ݾ���;�b�����!��s����Rp4������[����:�@Z��ҋ���=�ZN���G��d?�K�>[��A���#��m�ݾ������==������@�G���u����?ԦO?��V��=l��� ��� ��v<�k?�S���0������}Y={4���t��+�>C�w>e��� �_�-�a�pt0?�b?3W���䐾�)>�k���=T�+?_�?�h<QD�>�%?#+*��佮Q[>R�3>!��>��>��>���I۽D�?+�T?#g�W𜾆�>�=��'�z��`=��>��5��p輥"\>RZ�<!�����V�ܴ�����<�(W?s��>��)��za��}��3Y==��x?��?$.�>o{k?��B?դ<'h���S����aw=�W?4*i?��>����	о_���E�5?�e?��N>�bh���=�.�^U��$?�n?5_?]~��)w}����o���n6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>���������=	 �����?y.�?p���4�������d^��
�r���_TR=���m!ѽ�	��B7�aVɾ�e�}l��94�5��>��@*�5�%��>M��#���пy��VC���?�����>^��>�&���˾��u�������B�:�$��ӆ�AM�>x�>��������P�{��q;��"���>��?	�>�S��&������*�5<��>��>>��>�,��轾(ř?Ic���?οP���۝�}�X?:h�?�n�?�p?hz9<a�v���{�\��	.G?��s?�Z?Ss%�^>]�Z�7��Mb?	����3Y���4��:O��->��.??�>�ZD�N1�=N�>�?D}8>�7�Μȿ�V��A��@�?ͻ�?հ�u��>{'�?L�7?�X�BF���e��%�0����L?��V>�1���-'�<�6��~����>�6@?����B�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?K%�>��?�r�=�e�>�[�=��2-��i#>�$�=��>�p�?ϤM?�N�>K�=�8�/�ZF��FR�a$�@�C��>@�a?��L?GOb>*��k2�3!��{ͽ�d1��b鼲`@�|�,��߽�&5>l�=>>��D�Ӿ��?Mp�9�ؿ j��$p'��54?/��>�?����t�����;_?Qz�>�6� ,���%���B�`��?�G�?=�?��׾�R̼�><�>�I�>A�Խ����]�����7>1�B?Y��D��t�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?pQo���i�B>��?"������L��f?�
@u@a�^?*����������ھ�s��	��=��=��H>��
93<��I>��|=��=�>� ?"Au>��>f��>�ُ>�5=q�}��U����`+����f��#��=��u�Aj��|r���x'�_�;���ď� ���P)�%M/�q1ݽL@�u�>'�W?�X?�A~?Ϣ�>@S�uK>k�߾d/�wܽdE�=׶�<+5@?�E?} ?� >�z���hV��q�������aj����>��C>��>�O�>��>�VH�(f(>+&/>��M>?pD>�h�=!�=BL�=�>��>��>�č>q\=��H>����\G��bSz��λZ߸=Ѳ?��ǽ�+��6��A�̾PM�� �;ZX?S��>?.��(޿vF���L?�B!�\@3��O�U?p>�!P?�h?���0N�a=�?N>&E�����K(=��#�h�߀Q��T>;�?g�f>s1u>Z�3�L�8�u�P�����|>ZA6?ⶾ��9�m�u�:�H��bݾ�M>��>��@�X��������i��{=�r:?�?����t����gu�}\��j�Q>��\>q�=��=�]M>��c��HȽ�H��-=��=� _>�?`�>>`�=�?�>삝�D�j���>�O<>�v.>�F?�%?�9����=⊾",&�i��>�>F�r>���=�K��i�=���>��m>�;��ʁ��;߽��5�0
B>�a��i�c�h�ϽH�=�6����=���=�
 ��)� � <�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>|x��Z�������u�|�#=R��>�8H?�V����O�n>��v
?�?�^�ᩤ���ȿ8|v����>X�?���?f�m��A���@����>4��?�gY?doi>�g۾3`Z����>ֻ@?�R?�>�9���'���?�޶?ٯ�?	�`>94�?�q?5ݧ>�&G>P�4�3�Ŀ�$��k �>���=8>��>�&��s��@��<���D�bվ�`�>nǬ=F|�>}��n��
���>��������3��>$Қ>EHk>cOX>��4?:��>>�>4"�=tW=ŚҾ'_����K?���?���2n��M�<���=4�^��&?I4?�d[�U�Ͼeը>�\?^?�[?"d�>3��G>��@迿-~��Q��<��K>(4�>�H�>�$���FK>��Ծ�4D�Tp�>�ϗ>J����?ھ�,���Q��VB�>�e!?���>.Ү=� ?!�#?��j>e'�>4[E�[9����E����>d��>�G?b�~?�?2߹��]3�`	��S硿�[�=N>��x?�T?˕>��������[�E��
I�M����?fug?j6�o?g0�?S�??ңA?n%f>���ؾ����I�>Z�!?��ûA�JN&��	��~?Q?��>�8����ս-hּ����~��0�?�(\?eA&?����,a�a�¾(E�<f�"�$TU��O�;r]D���>*�>`�����=>�Ӱ=�Qm�]E6���f<a�={|�>���=�)7��q��0=,?��G�~ۃ���=��r�?xD���>�IL>����^?kl=��{�����x��	U� �? ��?Zk�?b��@�h��$=?�?S	?m"�>�J���}޾6�྿Pw�~x��w�Z�>���> �l���K���ڙ���F��_�Ž�WD�l��>��>d��>Y�?�=�5�>rt¾O�4�������ƾ��;��+�'h-���.��'�7���,���+�=�;���j���D�>J����>�?��>F�I>��>3��]K�>�/5>h��=���>c�|>��\>��>n^^=*��KR?����$�'��������g3B?�qd?S1�>ti�<��������?���?Ts�?=v>h��,+��n?�>�>H��Wq
?zT:=9�;�<V��y��3���1��>E׽� :��M�Enf�wj
?�/?�����̾�;׽푾���=9�?l�0?_��B�d��)n��V�J�N�Ӛ"��/��<.��:7F����ݐ�Dᆿv���G��6p�=?t�?������^��a�5eb��}s=Y)?�ԕ>UV�>X-}>�^1��.���d�:A��*�?��l?��>	�T?L�@?�O?�D?��x>�B�>0J��O�?�i�=>�>9� ?VA?��;?2�3?�@$?�A?Cn>�[	��X��L�ؾV�?F.?K�?�
?r\?����>�Y�/Kc��i��*��q^F�Q>��-:��ǽ$�"� ��=YK}>�W?��j�8�����dk>
�7?��>���>:���+����<��>�
?�E�>s �C~r��b�7W�>���?X��{=�)>i��=���к�\�=�����=
^��x;�>g<ww�=���=��s�+�y�@��:]��;�j�<�t�>:�?œ�>�C�>�@��3� �p���e�=�Y>8S>u>�Eپ�}���$��|�g��]y>�w�?�z�?-�f=��=��=}���U�����.���
��<�?EJ#?,XT?\��?t�=?ij#?ҵ>
+�cM���^�������?��&?�$|>eo�7`�����|)�8�?	?! r�����!��%��2���*S=��I�jE��(���6)6��V8>V6
�Hl��P/�?$S�?Tٿ�/�G��=׾uK���N�F?J�>d �>gX�>�,���h�}L$�s�><��><�e?C��>B&m?嫀?�O]?!gL>�[7�����jK���ر=sE>��O?l�?��?�z?�B?�)�>��=�ص�Գ	���3��j����2ް���>lK�>�
�>Z��>�fz>C��/��O��H=1�>�J�>���>��/?��>�>��G?
��>�]������뤾6Ń�=�ۜu?Λ�?��+?9Y=	����E��F���J�>ho�?���?04*?7�S�:��=��ּ+ⶾl�q��%�>۹>�1�>�ȓ=�zF=�c>Z�>��>�(�a��q8��OM�w�?�F?���=3�¿��u�ɸW��v��穵<������R�< ��=
e���=���F~
�_���1�W�K��cN��o����ّ���]�2��>�?T=�T>�:�="��;�4�'�@<'1�=9�z<��=�VC���������sļqa�р<�d%�ZW	=Y�C��˾�w}?�7I?��+?�C?2my>/L>{]4��w�>y��xB?PV>ԄP�����њ;�/�������ؾ}[׾��c�Ο�d>u�I���>�d3>v��=��<�l�=� r=Aˎ=�SY�p;=؟�=9y�=�=���=��>�*>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>ܭ7>	">��R���1�Ϝ\��b��zZ���!?PI;��H̾8�>��=),߾?�ƾ��.=�6>;ab=�g��U\���=��z���;=�l=}׉>o�C>�w�=�0��F�=�I=���=|�O>D��F�7��*,�c�3=���=W�b>G&>	��>�S?͑0?sd?���>��n�"pϾp���`�>�;�=�Ա>-�=z�D>Sڸ>�$8?ظD?��K?U[�>]��=Dܺ>�"�>�p,���m�	���R��`��<r`�?Mц?�{�>;�f<%�>��p���=���ý��?��1?'^?MB�>In���࿇ '�uB.��z����º�
=+�n���C�o΄�������T��= �>��>tA�>~t�>�A>{�E>�%�>�C>�#�<N[�=s�����<긫����=��z�͛�<(���XM;C�7u��_�t��u�;�M<�Li<q��=$��>lR>���>���=���<:/>Ի����L��'�=�.���1B�� d��A~�N/��D6���B>�2X>]���/��)�?�Z>	`?>���?w;u?y�>i$��վ�P��OMe�"�S�1��=2	>N�<�(m;�%O`��M���Ҿ* �>�1@>+U�>��2>���]�M���>�kо::w� �?Ń[�o+�=�⧽gbp�hF��uۥ��Q�/tT���c?)}�obC���?��A?��?�ӏ>��˼\�ݎ�>�l*�i>�n�nm���Y�=�K4?k�%?@?G~|�A(k��H̾���<߷>%AI��O���s�0����η�g��>������оo$3�qg������$�B��Lr����>3�O?�?W;b�^W��.UO����6"��qq?m|g?&�>J?�@?�%���z�<q��Wy�=��n?o��?�<�?W>�U�=��(B�>8?��?ߜ�?Tqs?S]T����>�;l�/>�g��R�=U>\�=<z�=�
?	�?�
?�塽F
���!G��6 {��=���=
|�>0%�>']W>�t�=oQg=��]=�c>}��>+�>��j>@��>-	�>󺿾��&�e�&?�?<hВ>�S!?,�>� ݼn�1E<5u�=W��t����і�����ނ�ᯇ<=s�=���=�>�&�����?׈\>���A^1?����P�=�~b>�8>>�Jۻ��>C4>>�^>���>���>��
>�k2>*�=FӾ�>V��5e!��,C���R���Ѿ�~z>���
&�J��a{��wAI��n��Ng�]j�n.��{<=��˽<H�?ռ��X�k���)�����ғ?[�>]6?:ی������>8��>zȍ>,K�������ȍ��g���?K��?�;c>��>W�W?+�?t�1��3��uZ�"�u�n(A�=e�M�`�y፿����
�q����_?��x?%yA?T�<!:z>a��?��%�Mӏ��)�>�/�S';��<<=�+�>*��J�`�8�Ӿ�þ18�:HF>>�o?5%�?�Y?TV��Zm��'>N�:?�1?sQt?��1?ő;?T����$?hR3>9I?~s?�J5?�.?	�
?�2>c.�=����(=�3��m�V�ѽ,�ʽ�񼠻3=.z{=W ��,<�s=v��<Av���ټy;@���G�<�<:=�Т=�$�=�Ԧ>��]?�`�>؆>b�7?l.��j8��ɮ�A*/?�R<=�]��-	��/^��^���/>�k?;��?JZ?;�c>�A�
C�1>Jc�>�&>�@\>0��>�k･pE�^U�=�>ذ>��=+�J�ȁ�ѩ	� Y��#�<�	>���>�0|>�
����'>�|���1z���d>%�Q��̺���S�'�G�@�1���v�Y�>��K?��?��=1_�M.��,If�?0)?�]<?�NM?��?��=a�۾j�9���J��?���>�M�<��������#����:���:��s>�2��z��Ic>�~�	-޾�n�J���66R=�W�	6U=����
־$����=��	>5i��U� �����Ѫ��I?_�k=u����W��A���
>���>6��>z�8��z�,;@��+���=�=��>7K;>g�����RG��'��Gz>�mK?�cZ?"A�?��<���u��9��'޾iq��t�i<�k?H�~>6��>��=��=❦�����(�j��M�6o�>/7�>��� �X��o���`��ڭ	����>�^�>x��=h�
?�uM?�?[?�)?]�?C�x>8��w�;�&?���?�i�=�KԽ,T��&9�L�E�{Q�>2K)?��B����>7G?�g?>�&?�[Q?��?;�>4� ��i@��a�>�B�>��W�gd����_>xJ?_s�>�hY?���?=>UB5�����Z�����=>��2?��"?A�?�c�>Ԩ�>������=���>�c?�0�?��o?��=�?t:2>���>@��=���>8��>�?XO?��s?Y�J?���>��<�7���8���Ds�C�O�bǂ;�nH<�y=���3t��G����<� �;�d���K�����D�������;��>̚=9�l��a0=�����u��?�>S�=�a��|��dr���h>h�>��>5��>��=<�|���>r�>ܽ�)*?���>�?���-m��������x�>O]?g�q>^�m�����׎�૽k�q?Bl?eOy����O�b?��]?<h��=��þq�b����g�O??�
?4�G���>��~?f�q?V��>��e�):n�*��Db���j�$Ѷ=Yr�>MX�S�d��?�>n�7?�N�>(�b>%�=lu۾�w��q��h?��?�?���?+*>��n�X4�alӾQb����@?��>�`��SO?��<��ྗ,�������雋�������v��\���U��o��9�;=J��Y�?Hl�?�׀?`�w?�>ھ�hj�f��)����L�����	���H�d�L�
�G�i�d�/��l�ƾQ2m��>�e~���@�?��(?�.�3�>�l�����Jξ�>?>N`����Ӟ�=�ߌ�Q�4=��U=�.f�n�,����V�?}X�>"6�>�Q<?[��>���0�8�7��[����3>�"�>�E�>9U�>���:�u+��W㽓�Ǿ�ヾcAֽ�e>��_?`~O?٨t?�K* �,���<�!�����J��ؚ>��y=��q>�t�P�R��1%��50��Rj�����O��~*�,	>��2?���>�"�>���?r�>`��x���9���$���<�K�>��b?h��>G�>�[��L&�^6�>��_?���> F�>�����1��\��ԙ���>~�\>��>�{Y=@3��KV��+�������[4���N>\%T?[�u�}������>#Q_?Bqѻ�{>t�>�03���-F���X-���>*?���=:�>_�˾&	ҾH��\����-?eY�>GV��N�'�@�=>�,?�?\�>�Y�?b�>�Uξ��'=��?o�b?�U?�rB?o��>@��<Dm��V̽7���?�"b>
<I>]�3=P�a=�:��w���D�j�b=��=;�����I�V<r��؝<�h|=��5>�Z��9�kK�W(�ߏþx�p���6�vм��-�VY��%����O�Bǘ�Rl�O��RJ��&��=�ƾ�=y����?�o�?��߾����V݋�]~�[�$��>�Z�����|@ �)/�b蔾�!�����}&��3I���m���\��t%?kz���3ȿ'���l�ܾd�?��?v�w?�9���"��F9�U`)>Em�<�)���������.ϿJ��W�`?�i�>\-�	o���z�>���>�zZ>w�n>\��j,B�<�-?q�.?���>��q�FhɿT-��M��<0��?a4@P�F?��L����]��=� ?4?�>s�J�/����ྯ��>��?�4�?DL>]�_�.3b�?WF?�T>d0+�!�;Z�>�\F>�5p:+�S�QE�>wnY>\>�;�a�x�H���>vĠ>s炽�,%�ۘ��Am�=j�j>�p�	�;Մ?e{\��f���/��U���V><�T?�*�>�H�=6�,?F5H��|Ͽ�\�*a?�0�?��?%�(?7ݿ��Ӛ>B�ܾ��M?�C6?^��>Ee&���t�Ѡ�=���7_�����H)V��
�=���>��>�y,�����O�[`��=�=�D�"漿 	���*��~=�zR>߳=1��TX��Π��yq�AHֽ�t�Gta<���=�o>Z`~>�(>Qy>1�h?e�{?3|Y>���=�����ݮ�B��� ��=��\��Jm�͏���r���������ɾ�W�F4��'��S�4P��u�=uzU�Ô�p
�3I��6�j�,? �W>q�ݾ;�S�?(�<�IѾDB��5EF�fʽT�ھ�D=�L�j����?��G?5��9�]�L8�B�������D?�)}�z��O$;��>�PP=��=1+u>IvI<{���N.��@�Y/?��?|1��4�����*>�d��=P�+??�9j<6�>�f%?�4*���߽Z>�1>�z�>~��>}�>����Wy۽V?ܭT?�c��&����>a���7ty���Y=�&>��4�
�R�V>K �<��$n?�����s�<}"W?���>i�)�M���T��UG� �==&�x?G�?��>�ak?��B?���<�X��+�S�Q'�"�v=I�W?� i?`�>R���оy���C�5?��e?[O>�$h�)����.��K�� ?��n?�\?�)��3m}������_t6?g�v?js^��t��m����V��F�>=S�>���>\�9�Pv�>"�>?�#�G�������X4��?X�@���?sO;<���Y�=�C?[�>�O�l>ƾRw�����4�q=�)�>����&lv����D/,���8? ��?���>7�����xx�=�咾�3�?Ӿ�?���9�W;;m��m��O��)�;�o�=�'-��"Z�E쾓�8��̾��	��<����¼�=�>"F@8�ǽI�>V
3���ῗ�Ͽ����%վ2>x���? Ӟ>�Ƚ	ۦ��$h���n���B��iD��){�$�>X�5<�
�>��A�����-�x��<u�N>>ļe�?"v�=D��������;\�>�%2?��?�1�p�P���?(u%�f����ͤ�![�a}:?��?�|�?Lc�?���>W%�(������~�"?�$�? �Z?�eV�&������j?�a���U`�>�4�XGE��U>b"3?�A�>��-�9�|=z>��>�n>"/�,�Ŀ�ٶ�������?]��?�n����>l��?�r+?_i�K7���[����*��E-�\<A?�2>Պ��'�!�G0=�HӒ���
?.~0?�{��.�nk?�op��ݾ02"��
��?��>:�>!�?��+>X�f�[)6�lQ-��?���?m��?Ԭ¾��+�/;?΃n>	g���
Ͼ6P�=�ű>~� ?��l>�[~=���>a-}�ġe�%��>���?��?��>�?���n�����>P��?���>'�?���=�"�> �>�m˾8�e��/+>2W'>Gk����?]�O?b�>�U�=S�/�~����;��vN��x���9�u%p>�i?�K?�4>���G��g)�$���?��F��;9@��8���T���>�X>6'.>#�?���¾��?D����b>��;�Y�j�@?4�d>��>�����ea�����v?�:�>�[�Zh���폿@�E�]��?x�?�P%?���Ӻ^�Z>r�>]?�>�K�N��fp���w>�sM?�\��Í��Xc�x�>���?B�	@�:�?i�z���?�4��ؙ��·�Ĝ�G�<Bv5=_x?�S��?�>-�>�K>pd��9���⃿�m�>�R�?s��?s�?0}?(����\[ >2 �>ϖX?�U�>ygu=���Yզ>�?H�:���kվ�j�?��@��@��(?��Ӊ��K������*���߀=+��=#r"=��F�o	=\��=�1>R�=���=��]>15(>��`>�P�>�>��>����$��]��A�@��/
��Z ��i����s����ᩨ�e2��(���"��W{��v��H��"$�
)�=ָU?~�Q?��o?r� ?k~���>�����y==K#���=\�>�1?L?�*?L��=PV����d�n��~��Җ�����>s�I>7�>�{�>JZ�>��q���H>@>>��>�� >� =��Z��Y=��O>�'�>�F�>�й>Y9<>�>%ϴ�92��A�h��w��̽� �?�}��üJ�2��X8��(����^�=�`.?�x>���?п����3H?����r+��+���>��0?�bW?Ϙ>,����T��3>$����j��`>0 ���l���)�C$Q>�l?Y�f>(^t>��3��Q8�0�P�BK���}>�C6?w���$9�w�u��nH�!7ݾ�gM>F��>m;Q��V��Ė�o��0i���z=қ:?"�?C᳽=����v�۞��\R>�p[>�=�J�=G�K>sjd�k$ǽ��G�a�.=~��=��]>�! ?�.5>[��=U��>��B�a�!��>�*4>�8>�69??�?��?�ʲ���B��Ó4���h>*%�>̬�>(>;�F�z֡=LG�>B�`>_-=�ߓ;������`��*U>5!y�;�Z�������=������=H�=L��g&?��=~�|?�¼�����DԾ��q���3?P\�>��=�L�=�A��%���>d�Z��?��@���?Y�8��i�V�F?��?�����f�^�:>�&?�><��ɾ���>7`!��쟾����<;j��?���?�$V�h0��9'����>�J?�̨�x*�>#ӌ�����1��|�j�	&�=���>.�?D8��?��ok��M#8?��
?�����;Ϳ���� r�>/��? (�?e�l�Ac�� ��jݼ>[��?�6?�?�=eM��쩽:��>�C?&G1?�F�>��#�d����?M�?�y�?��/>�$�?M�d?3��>o<��3�TV���ˏ��-s�H��;�>���g����M�����n�k{J�3
�Ԉ[>G٨<���>]<��Kӵ�;*=��L��L���x�=ǩ�>��;>��U>w��>���>�Ϻ>��7>��Z��vݽ4a��k�����K?���?)���2n�N�<G��=)�^��&?�I4?�k[���Ͼ�ը>�\?l?�[?d�>4��L>��F迿:~��D��<v�K>)4�>�H�>K%��oFK>��Ծ�4D�Up�>�ϗ>����?ھ-��!T��=B�>�e!?���>bҮ=�� ?��#?��j>�(�>�`E��9��J�E�f��>��>�H?��~?m�?�Թ�sZ3�����桿��[��;N>u�x?�U?ʕ>A���҃���lE�E>I���w��?Ctg?'R�(?#2�?�??6�A?1)f>��ؾf����>��!?vj��kA��^&�TG��?�?Z.�>M��-<ؽN ݼVM�����3�?��\?_Z&?��r�`�XR¾�<["���b���;h�S�xs>�>6� ڴ=i>T �=QJm�!]7��7<Dɺ=��>���=�v7�����~%4?�P�<#����V< �h���W��>��3>@��"��?� >,�r�� ��5g��������?pm�?���?� ���\� o?Ui?�q??�Ae?\a���""�"A�����Ͼ�c��/�=ǃ>���<�x�����!��^p���Baн�\?�-�>*�3?���>Ŗj=C <w��9�P�LE�B ��k�����=(��3������o=+�<���1VG��\�>$]½	��>�� ?>P�>��=n�>@�= �4>�>�A>�c�>��>�)>j�;=�9=#u��+�b?H�-�U�X������Q?t�Q?h�F>ͩ[>�.v��M)�U9N?'ȩ?���?�R�>�!��+.��	?�s�>&Ug��Q?.8q=�Ai������h�D�*��1�����~Ls>�8ͽ�C$��W��$��*m?j�?G�>�>ܾp=T�T���V�p=�؄?�<)?`)���Q�S�o��dX��S���(��9j�&���61%���o��ȏ�Jf��@���s|&��U*=h�)?�?�� ��=�c�����k��:@�ib>���>���>���>jC>'1	�e�1�?]�.�%�F+��
�>�|?�!�>��I?�;?�NP?�L?�h�>�}�>������>���;�>r��>`�8?�\-?\�/?�]?�*?:`>_=󽮣���&ؾd�?V�?t�?f?X�?�І�[`ƽ�B��W;����y�=Ƈ���o=�Һ<h�ҽыn�A�P=@�R>k�
?�U^���=�r���M4x>�-?bo?F��>�J�a����_�>X�?/�>���V�~�GS	���?�Qf?rb<�A	���'�>��=e��ND�=�]>���t�=�x�;�|�<S��=���q��=7�=vW�=rI�<[��<��ɽ���>!z?�؊>;��>����?��$�-<�=hL>��O>^�>�Qݾ���������g��4v>�\�?B��?��q=��=�W�=�-�����B��6F��@k�<�?�Z"?�R?*��?
�<?�8"?��>���.J���؄�������?�,?�h�>c��Q�ʾ]騿�z3��?�a?�9a����m8)��s¾��Խ��>�R/��.~�������C�u֌�_��|���?���?��A�s�6����Ř�_J��.�C?�"�>�K�>��>G�)���g�8�p7;>�|�>�Q?�>�O?�8{?i�[?�|T>�8�n/���Й�J�5���!>�@?���?��?y?�a�>u�>�)���F�������ނ��V=wZ>���>�*�>]�>X��=��ǽ2P��n�>�&h�=�{b>H��>���>Q��>|w>=��<."L?�<�>}������-�%%��{+�=��u?J��?ӢM?:;�=�s��>������>�ظ?�"�?0�?���l��=��+>^��f" ����>�E>�V>��v� ?w����>��$?$<�==���~���Y���H��xC?tDB?��ȼ�Kſ�Nq�^r����}'`<c�_�2���7|]���=�����G����t�Y�����Д�Fõ��.����}�!�>)�=q� >���=�'�< 庼r��<&�/=�<~�=j�j���k<�?O��� �V����|�d0b<�TH=�8�!�����?П�>.��>�0n?�L3����=Gk?��">h�,>t�]?��l��R�a���=8�=N�����*);�6ɾ��7��\@�v֔<�kV����=��w>�A�=���)h�=�_=?U�=y~a=ܙ�=�H�=��=�D�=��M=���=���=OAv?����Q��Jj�ZMd���T?j;&>,s$�����
n?�b:>ws������tfl?���?a^�?���>����L�>/U����>��C=>晽��>^�{=���2��>ܡ&>#�!��쮿����?��@�R?ۉ��_�ֿ q�="�2>�>}�O��O/�H�R��Bf�O�L�-.#?!�:��sɾ���>���=�ܾ��¾x�!=��)>ڭT=ce���[��*�=Xj��g=ڹv=��>��G>���=�ǽE~�= -=�<�=Z:N>h킼��9���.��7@=n��=׍`>��>E��>q<?r�6?�sf?7�> �r�	Ҿ]q˾L�~>S��=B�>�Q=|@>��>�1?�C?�P?�h�>g�,=��>�>>�*�6t�yb�Ṯ���<i_�? +�?���><�I=C3@�I��o:�����?'Q3?QG?35�>&��y�ݿ#m��Z1�Т���e=ƭ7=�J��U���@�Ō���Ě�V�=ݥ�>Ί�>H��>^��>��7>��q>�	�>�6)>w�-<܆^=׿�<ʨ�=�N=0��=�伕�M���b6�<�3ﻟK�?e�5m��v
����t���+;�>p��>�WH>�W ?Z�5>��2PU<�o����L�;2�=Nf��6�E�Zgj�n!}����
�Ƚ}ֈ>@��=�]������SN?Jnz>#5�>uY�?�Sd?�%_=n]���ľ����o[̾z�z��P=��>a�H��O��^b��c[����� �>�j�>�>k�u>��*�� <�m^F=+O���5�&�>����bS@�Z0��up�ZG������Dg���'C?������=��?4K?W\�?��>�.����ݾ��)>����.�<o��p�o�JF����?�F&?ޥ�>i��h�D�#�˾�u���ܸ>yrG���O�[����0�b�7��A���+�>tܪ�PѾC�2��J���폿z/B��$p��G�>~O?��?��c�_:��Z�O��&��a���e?�`g?�[�>�?��?.9����쾌1��3M�=�o?���?Z��?Kr	>6��=�[���T�>Q�?飖?
v�??os?i3>���>[6�;� >�^��f��=��>���=���=�?��
?��
?����*�	��p��W�a�^�<#=�{�=��>	�>�ds>lM�=uj=��=�\>$�>��>؄d>'�>�B�>����gm���?�-�=���>��/?3̋>�]�=��ν��<��u��31��3$�ǟ�!罍���e3��<�=�O(����>SĿ;�?{Ee>����?��@7���DT>1�D>Ȫǽ��>�S!>2�q>�G�>�C�>��>.G�>�>5����� >z5�*xD�59 �6f4��+��uH>pQ��>����7��E���j������8�y��`����;�]T�o��?�&�;R��� .��a��<��>���>J�?K[��V�I=�>�%?~��>�6־a���EL��g��G��?K��?Jm1>��>
h?|�I?dǙ��3��6�a�J���h��9q��rT�������g�h�� X����?��Z?�W?94�<�tu>�YX?�*��&���9>N@Q����7>�3|>��ڽ������پ�C
�"E�}�b>o�s?:~?*?����&�[$�>��?T�?؊k?u�?�U.?+�>�?[<=>��7?
�?�6?b(??�>�>��_<p�,�<h�=*�����l���E���f��;ƽ���9�<z�{�=nF
�K�<d��= ���=|�9�><a��<�|�=�'>b�>-�^?�1�>���>U�+?����k4���Ѿ���>��o����@پ�ž�'����<�=?�q�?'i?p#�>��K�'q�"�>��>�ҋ=�{>��>�.�I��R�=���=0h>][#�y��2n���ܾi"��ƞ�<}a�=�*?�^2>`ҭ�<�=*���wC���bj=�Ȕ�q���G����Q�#(���g��>��.?�Z�>�q>����ҁ��}f��3?�u?�<M?]#�?�����w�_H���M��^D����>L��i��N��P���A�D�G9h�g=�>�-���(����R>��������]��C�(H𾵹�=dz���u�<�>�Js��d�<�5�=�^>k2��Z!�㩑�������Q?(A�<�ݒ�J�J�w��>�ª>�´>T�(����I�>�T���53=77�>�4>#�l�����FM�EO�p<�> RE?CV_?}i�?1��Qs���B�����b���ȼ��?�v�>8c?AB>kح=������d�G�}�>��>���A�G�D1��a'����$�c��>�7?�>7�?�R?��
?a�`?�*?�D?�)�>����9����A&?/��?��=��Խx�T�y 9�F�`��>?�)?ʷB����>*�?ҽ?��&?�Q?޵?>�>�� ��C@����>iY�>��W��b���_>��J?ښ�>n=Y?�ԃ?��=>?�5��颾 թ�}V�=>|�2?�5#?B�?寸>���>���� ~�=��>�c?�%�?�o?R��=w�?s2> ��>�=���>�v�>k
?PSO?��s?��J?	|�>�w�<-W���	���:s���P��};�[G< Oz=����"t�́� ��<��;�����e'�E�u���}]�;���>(�v>�ڕ�s�3>�m¾�����C>��ռ�4���򊾤b@�gߧ=�J{>S� ?���>���Ɗ=�>�=�>S�e*?jh?��?�!;<0�a��Hھ-�J�L$�>�A?��=�m�?���B�v�<�e=J�l?t]?y�R�+��0�b?��]?�f�=���þӸb����]�O?��
?h�G���>:�~?��q?4��>��e�u:n����Cb�{�j��̶=�s�>X���d�J@�>��7?�N�>#�b>�#�=qu۾j�w�"r���?H�?��?���?�**>��n�54�=���:���TZ?��>�����?8���R�Ҿ߃�����U��{������b���ܥ�����s�������.�=�A?nw?Q)m?HWa?���6�c�2X��~�{V����~� 2I�B�W�E�V�n�f�������^��=��}�T�@�}��?�?(?Y0��J�>U#�������ξ��;>����o��Rs�=�A��<�4=
%W=�<k���/�R譾��?�շ>���>�k<?��Z��=�j�1���6�6\���1>��>{2�>N�>9�; �.�
潪�ƾK���ս�U>:�b?�RP?iBg?����e!�s�{���#�K4�],���w>��%=���=�N���`��y*�4�A�w�D��C���[��>�p??&H>P��>�/�?L�>h���H���᜾���[;��>��V?���>�^>�I轨��[H�>)�n?��>�%�>��������y��3�He�>���>d#�>�/>\u��U�.p��}Z��S�:�~�=�k?��w��_|��z�>�P?#�����K=�f�>㬍��~���Ҙ/�vG> �>)�=�,>�^��� ���x��<���%'?��?̛��4�)���~>id?)r�>��>zǁ?'��>��þ�;ۻ`�?�2^?�/K?�BA?f��>bz�<�Ϋ��~˽�U'���A=�R�> PT>7{Y=F��=����X�i���1=�=[	��Rʬ�2><U���ѽL<�g�<pZ1>M[�}TM��?ᾦ���������Th:���'�S�_��K�����܆����&�44��2C=f-+��I�����~Cb�`�?<��?�|�{mﾞ���z�[��1��ۗ�>aF�ȣ���)׾۽2Y�I�׾~X��u���J���f�[3X���+?�Zپ��ǿh<��
�I�9?ʣ>?\Il?|^̾��A���3��e^>�24>�'
>�M׾_���ȿS�ľ(�q?:��>`��҂�=s?���=5�>6d]>�r������:���?��%?(5?6��ҿ����3(�=6F�?�~@��A?G�(��k�VnW=�P�>��	?EG>>=D0�p��I���8��>�@�?Hϊ?�F=aX�֜�q f?�+2<��F�D컗K�=�ۥ=>�=�9���G>p��>�L��\C���޽�4>G��>0^�Ew�7b_�#y�<�[>��ֽHœ��P�?g�d��aZ��O �΁��%)>�XZ?ݪ�>E��=��%?�N��ӿ�yH�>�}?T� @��?��?�mؾ�>i�ؾUE?�/?��>.�5�*Px�7i>��<���<9���Xp���D>�?� M>ʔ:����f��
Z<�L>d�6�ƿ�%����,�=�`��]��	��.��IlW������,o�K@罗�i=��=�Q>��>a�V>�Z>�}W?ϸk?��>��>څ㽎c����;3,
�������������>ɣ��M� �߾�g	����?���ʾ��r��(=��|�)��ch�v03�9�A��4?ջZ>�y(�} 0�M��=wzƽ��j�&h�=���<xW�y�)��;�;�?YT9?�o���z�l�;<����[c���9?aNU�����E��%A>��E:x�(<P�>���=�<��3>����^0?	V?�v���F��C=*>� ��8=��+?	l?�\<a��>�?%?I�*�6��Xe[>t�3>��>���>��>����]۽q�?d~T?K��m񜾮Ր>�Q����z�U�`=K>��4��|�\�[>%ԑ<8댾�HV�-��-2�<��Z?��>}�&��������d/˼h4�<!�w?��?V�>�,j?pE?���<~����W�z�����=n�]?S�b?�W�=��P���ɾH��y80?�X?)@>�U�C����71��� ���?=n?_�?ef�����o�����
�6?�z�?.;u�0p��UD���\��,H?�֩>�v�>��߾G]�>�H[?r�
;���=���A?����?��@¸�?�޽ ���/�=��>w;�>0��bĚ�vK�U!���c �,?�s���a��:��0w��� ?xmr?s��>qͧ������=tԕ��X�?��?5����f<s���l��u��_�<N��=a1�G`"���L�7���ƾ_�
�����±�����>Z@*V��,�>�48��4⿘QϿ����^о�Sq�3�?8t�>e�ȽF����j��Mu�r�G���H�y����K�>s`�<0"�=�K��ݏ��|Q�޷_=?��>/�ݼ�>��*�y�B��+��kE>g ?0ɼ>�n�=�μ�[��?�o�Q�п�j��I�.��7?x��?�Q�?su?o�>�X�c����=Q'?�h?�y?�h>;�����;AKo??ȭ���W��,���F�ل">g�"?��>r�)��t=!�:>c��>�M>;@0��ĿW���;���!g�?��?���ŷ?m��?��?���IX���z��4%����29?�D2>/˾Y��a�4�Yą�W*�>�<?c�D���p�i?�x� �X��A�>84�U��>���IPj�f���﫺~BI�2B�����.$�?jy@i�?�0.�k4<���?ӻ�>f�1�� ���>u!>���=�>�>uJ>}��>��'��'v����=w��?��?K�? Y���U���;:>���?��>��?,��=�X�>w<	>�d��nӾ���(>#�=�����>u�L?��>E�=�	A��(0��:B��MN��]���C��Z�>:E]?��H?�x>|��kZ�}�UY��LB&�)6
�I�<��9�0�ڽ�/>��@>g>H�8��پx�(?�F�K�ͿR���h>��*�b?#а>��>Z޾�h۾`[�=8�i?^s�>B
��&��L%��7w余��?���?_Y�>u����=��<��>r��>��|�I�X�m|�'��>�/s?w5�[����Đ�ˏ�=��?�	@�ͷ?*���=H?ݧ�$˅��q�����r��I��=p1&?�)پ��?>Q<?qp>i�d�8,���W|�V��>��?���?���>�\?��e��p/��N�����>po?33�>�`��l�۾U��>i-?;������Y����f?�4@�@�R?������ؿ�y���&��4#���et=Q�d=Z�&>h
�n9[=%��=�ޗ<{��<�xa>�j�>K&t>'�X>:�$>Bw)>�>>v����!��饿�㛿d�B��>�.�
���i�B�3�^����0������ln���m���~W��S#�>Ȃ����=��U?N�P?~�n?&�?ô��̡>������<?���k=���>��0?J?I9(?*%�=����%�b��:���������S*�>��H>̏�>�l�>��>VO#���N>N�B>�5�>� >�kS=t2M��o=�P>Zj�>jl�>5b�>�,,>��<�����qĿ� D�5#�6��:o�?.!���J��k��v�Ž�@����>x;(?�;>����YϿO���B�f?ma���6��_>�b ��tH?
�v?L%�=L���-�$�c#�=Cl���h��h�>p�ֽ�DȾ�5$�oE=֨-?]>�cv>.H��Y#���(�Tɾ�>�*?y� ���nh�W ?��Q��6�> �>��=%W����>�R��LM��*���;N?���>�M&�YG���Z��� ���(>[�>����թ�=�l
>߲-�_��$W0��=�+�=
�>F�?��*>�5�=
�>t��`hO�s%�>C�?>u�&>Fd??��#?U���Q��Yׁ��-+��2y>8��>��~>d�>��I��^�=Y��>��b>�	��Ӆ�@��?$?���V>���P�_�wUr�k�u=�ᕽ;��=�M�=R� �.[<�Rf=��?,���Vjt�g�̾�����-?�Y@?�=��=Ƿ��c���[վ+��?�@hp�?�t˾��S�29�>�?�?k��J*>ܘ�>�^>o������E?�Ո�|�"�����½?�ɖ?Uό���-es�{��=�� ?n����r�>���Z��D����u���$=l��>�4H?�K���P���=�|
?c?<N򾺩���ȿCyv����>M
�?$�?��m�6��H@�r�>��?WY?�Ei>�l۾�MZ�4��>��@?W�Q?��>HF��'�*�?M�?���?�d�=:{�?A�T?\��>F<��4�T*��{L��9��:-b�8k`>��*� n�u~L�����c��
�W����R�>��<D��>ޔA�l����=�9W;�N��!f7�W��>� >�o�>m��>`��>���>�P>,*/���1� hʾ9v��|�K?���?-���2n�dO�<+��=�^��&?}I4?bj[���Ͼ�ը>�\?g?�[?d�>;��N>��C迿8~��m��<��K>%4�>�H�>�$���FK>��Ծ�4D�^p�>�ϗ>q����?ھ�,��hR��EB�>�e!?���>�Ү='� ?H�#?��j>�(�>PaE��9����E�{��>d��>�H?-�~?��?1Թ��Z3�����桿Q�[��=N>��x?gU?˕>�냝�nE��OI�N���.��?.tg?�S�?�1�?��??8�A?�)f>ԉ��ؾC���P�>>�?*���LJ����j~�8b�>��?�t�>;���������5��|ܾD?{�^?�!(?���`�}����<����pB	<7���2���f�=a>mr��%5�=�>�	�=��^��2��JE=$�=���>P�=�I.�k՘�8�U?%���J�,|>b�]��f�.>�:ew�>��|�Z�W?� �G��
���%����\ c?a��?�v�?âٽ�o\��??f�{?UO�>�)�>a�1� �߾�Z����*뽾f6�q�=��>�P2=��Ҿ����Ŀ�����V<�t���(?B��>��?��>~���Kם>�C,�8^�Ux��?%���P�3�H���3��i	��T��}�a������>i��ȝ�*�>��<���>D|�>9j0>Y��=<��>l;����=�F�>CT>qY�=�v>!�>��>�(C>�'��KR?�����'�8�� ���3B?rd?�0�>�i�&���6��H�?���?Ss�?�=v>�~h��,+�(n?r>�>����q
?*Q:=�8��G�<V�����4�����>�B׽� :��M��of��i
?j/?*����̾^<׽!m���͆=_<�?O3,?f9&�w8N�l��^���V�Eĉ�i�z�����&�(�Daq�s9������t\���|&��x<=AP)?\��?�����{꾏d����j���?��_q>3�>���>�W�>s�/>Lk��;.��Z�+�"��h��}�>H.x?��{>#�J?��:?FcM? !R?|��>xX�>�O���/�>��<��>yt�>��9?�+?��)?M�?tE*?z�s>�|�Ϋ���ܾ�`?,�?[#?���>��>�o��ȴ轕������l�\�g~5��o�=g�=D���ƽ�d=	J>�?t�4�8��m��(Uk>[�6?^0�>���>f����o�����<�>��
?�o�>�����q�.A��b�>���?Z��=,�*>�r�=�������=����4��=�e��j�=��"<�=�6�=�fk��"'�IH�:l��;+��<ھ�>ʵ?�m�>�\�>���s �U���r�=Y�X>%�S>�>��ؾU��< ����g���x>!z�?ꀴ?��i==��=m��=����7�����㾾�p�<��?��"?��S?�r�?��=?�8#?�e>�6�Sl���v��d=��u�?� ,?��>����ʾG�؉3��?<[?�<a�����;)��¾C�Խ�>�Z/�i.~�p��kD�rօ�?������8��?���?�A���6�qy辵����[����C?*!�>dY�>g�>��)�?�g��$��0;>T��>�R?��>��O?�:{?�[?E�T>I�8��0��7ϙ�@�2�5�!>�@?���?n�?�y?�k�>��>!�)�oྼe��N����Ⴞ��V=U
Z>���>9%�>��>��=�Ƚ�D��K�>�"M�=��b>���>"��>z�>��w>�7�<-~�?L��<0AE��z���V��9N����	n?�|�?��v?C�3=q`��!����R�>m�?�>�?Vbm?v�{���J>.�м��v4H�d�#?��2?�>�<���z'2> J=���>��=?Q����O��bR漁N?j0D?	�^R¿,@�H��ƽ=��h�<�~�*�ﾇI�;L����TE���T�Yp����d��Խ���!�%���۾d�h����r	"?�ę���X=��&�K�>t[b��c�=o�0=4�>�,A>�� �v�"=�]ڼR���M�$��A@;>�l=��w=�YP��r��ޣ}?�^&?�i
?�!�?0t�8�=��>�>O�O>�Z�>G�>�(?>I_��t_��#��]�K�M@|���4����*�b�p�.=H�(��6>�{M>�_>hؕ�W?0>��=|^>"@y=}U>��=���=P[�=���=q#>��+>�Oq?����˜���,P�09S�_��?������h��­��yS??�������/��$�?�?�`�?�{>�ø���>�bV��D<�ڸ>)=�x�Ǧ=�����+>p4�>ί:��h������u�?�@c{K?ZT��|jؿM�Q>�'>��>K*X��+�7$C�Sf�ͽ'���?5a@��~��۝p>���=�W;L���#z�=}�R>�W=A�8���Q�~�h=ǟ����.=`�3=�hz>"�+>gR�=��^��q�=�bf=^��=�XK>�I&=����]J���%=?�=B�[>��>)��>�?�^0? Wd?7�>^n��Ͼ�E��P8�>�	�=z7�>���=�cB>���>}�7?W�D?��K?���>n�=��>��>ݘ,���m��h��ɧ��^�<��?�͆?�Ҹ>|R<��A�&��#e>�� Žr?�P1?�l?�>U��࿚^&���.�Y����;C�]�*=jfr��DU�����qh� ��](�=�r�>���>�>�Dy>��9>3�N>T#�>v�>��<2b�=?ϋ����<����ݥ�=�T��b~�<Lż<��n�&�B�+��������;$N�;�^<��;�O>�>��J>菻>�k�=<�Ѿ~�=��{���D���=/�����9�m�d��,|��R3��U��`0>�-+>h}0�ޑ�Xi?l�%>�c>���?r�z?o[K>����Ӿ^����T����a��g*=Ck�=d
�K(�C�L���I��JϾf��>ǹw>�v�>��5>��"��;i�oa��3|������>���Z�N<^S���m������w��N�\��#=��
?��R��>��|?�?(��?IS�>_����E>�ak�.��]�'���#��;�?�?^�>6�/�Te� W���?ϽO?��}��iG�荿��2���7�����3.>i˺��	L��4������l�3�5�9�ȕ�>v+?���?�U;@�s�td�Y�@��������>X`�?��>�uP?:�?*�������z����=�(t?`�?���?�=a��=CT����>�A? V�?x@�?;�s?Bn@�p��>��;�>�������=�
>���=���=Q�
?)?�
?�䤽�4	�1�����l�]��o�<-!�=�~�>��>�v>V;�=�Nm=3ٷ=��^>��>'M�>��d>�}�>\@�>ݗ��=���mF?� �=�@e>��?i2g>�$=�2[�]ۂ=�iڽsI�W��뺺�]�P�� �=
��/4Z�j	�����>�S¿�d�?R�P>@��9%?H9�$.2�Z�I>�=�={���U�>��	��z>X@6>��>5�>���>\_(=U|־�k>�+��#�6�B���Q�8[Ӿ�{|>أ���X.�HQ�d����C��᳾��ʭh��1���<����<}�?c4����l�F +�����=�?�u�>5?X(��h���8�>�>�>���쳔��/��$�߾m�?i��?�6S>���>�\?g� ?����W8��kN��/����P�jm�$g��B��t\��>������Q?!~`?[3?��]=T	~>��q?����I����>�a0�D�<���=�{�>�����FD�_��?"�����J�:>��e?��?��"?R���N���{�>�!?e'?%?g?��>�N?�%>�v%?y�Y>�#5?�+:?�v?��'?0��><*k��m%=�I>��<(�ٽsaj�ي�F"��}��w��<�cC=^�׽��L�lּ/=�؃�m�H�}�	=;l=G6�=2����"�W�=r��>�a?���>���>�4?�(�@�/��i���n?/�3=����q������L��=�e??	�?�yX?�>��=�466��:>p�x>�{>��I>�R�>$-ѽ�	��r�=�<>� >T�=i`w�~#�aJ�M:�����<� >��>i">an����9>Q�;����$n�>U"��"������,|��j!���U��u?�X+?�
?w-ƽ���d���,a�඄?�T�>�A?3��?��D���о �#��i��0��W��>lV�����W_���l������<�>>fB��z��Ic>�~�	-޾�n�J���66R=�W�	6U=����
־$����=��	>5i��U� �����Ѫ��I?_�k=u����W��A���
>���>6��>z�8��z�,;@��+���=�=��>7K;>g�����RG��'��Gz>�mK?�cZ?"A�?��<���u��9��'޾iq��t�i<�k?H�~>6��>��=��=❦�����(�j��M�6o�>/7�>��� �X��o���`��ڭ	����>�^�>x��=h�
?�uM?�?[?�)?]�?C�x>8��w�;�&?���?�i�=�KԽ,T��&9�L�E�{Q�>2K)?��B����>7G?�g?>�&?�[Q?��?;�>4� ��i@��a�>�B�>��W�gd����_>xJ?_s�>�hY?���?=>UB5�����Z�����=>��2?��"?A�?�c�>Ԩ�>������=���>�c?�0�?��o?��=�?t:2>���>@��=���>8��>�?XO?��s?Y�J?���>��<�7���8���Ds�C�O�bǂ;�nH<�y=���3t��G����<� �;�d���K�����D�������;��>̚=9�l��a0=�����u��?�>S�=�a��|��dr���h>h�>��>5��>��=<�|���>r�>ܽ�)*?���>�?���-m��������x�>O]?g�q>^�m�����׎�૽k�q?Bl?eOy����O�b?��]?<h��=��þq�b����g�O??�
?4�G���>��~?f�q?V��>��e�):n�*��Db���j�$Ѷ=Yr�>MX�S�d��?�>n�7?�N�>(�b>%�=lu۾�w��q��h?��?�?���?+*>��n�X4�alӾQb����@?��>�`��SO?��<��ྗ,�������雋�������v��\���U��o��9�;=J��Y�?Hl�?�׀?`�w?�>ھ�hj�f��)����L�����	���H�d�L�
�G�i�d�/��l�ƾQ2m��>�e~���@�?��(?�.�3�>�l�����Jξ�>?>N`����Ӟ�=�ߌ�Q�4=��U=�.f�n�,����V�?}X�>"6�>�Q<?[��>���0�8�7��[����3>�"�>�E�>9U�>���:�u+��W㽓�Ǿ�ヾcAֽ�e>��_?`~O?٨t?�K* �,���<�!�����J��ؚ>��y=��q>�t�P�R��1%��50��Rj�����O��~*�,	>��2?���>�"�>���?r�>`��x���9���$���<�K�>��b?h��>G�>�[��L&�^6�>��_?���> F�>�����1��\��ԙ���>~�\>��>�{Y=@3��KV��+�������[4���N>\%T?[�u�}������>#Q_?Bqѻ�{>t�>�03���-F���X-���>*?���=:�>_�˾&	ҾH��\����-?eY�>GV��N�'�@�=>�,?�?\�>�Y�?b�>�Uξ��'=��?o�b?�U?�rB?o��>@��<Dm��V̽7���?�"b>
<I>]�3=P�a=�:��w���D�j�b=��=;�����I�V<r��؝<�h|=��5>�Z��9�kK�W(�ߏþx�p���6�vм��-�VY��%����O�Bǘ�Rl�O��RJ��&��=�ƾ�=y����?�o�?��߾����V݋�]~�[�$��>�Z�����|@ �)/�b蔾�!�����}&��3I���m���\��t%?kz���3ȿ'���l�ܾd�?��?v�w?�9���"��F9�U`)>Em�<�)���������.ϿJ��W�`?�i�>\-�	o���z�>���>�zZ>w�n>\��j,B�<�-?q�.?���>��q�FhɿT-��M��<0��?a4@P�F?��L����]��=� ?4?�>s�J�/����ྯ��>��?�4�?DL>]�_�.3b�?WF?�T>d0+�!�;Z�>�\F>�5p:+�S�QE�>wnY>\>�;�a�x�H���>vĠ>s炽�,%�ۘ��Am�=j�j>�p�	�;Մ?e{\��f���/��U���V><�T?�*�>�H�=6�,?F5H��|Ͽ�\�*a?�0�?��?%�(?7ݿ��Ӛ>B�ܾ��M?�C6?^��>Ee&���t�Ѡ�=���7_�����H)V��
�=���>��>�y,�����O�[`��=�=�D�"漿 	���*��~=�zR>߳=1��TX��Π��yq�AHֽ�t�Gta<���=�o>Z`~>�(>Qy>1�h?e�{?3|Y>���=�����ݮ�B��� ��=��\��Jm�͏���r���������ɾ�W�F4��'��S�4P��u�=uzU�Ô�p
�3I��6�j�,? �W>q�ݾ;�S�?(�<�IѾDB��5EF�fʽT�ھ�D=�L�j����?��G?5��9�]�L8�B�������D?�)}�z��O$;��>�PP=��=1+u>IvI<{���N.��@�Y/?��?|1��4�����*>�d��=P�+??�9j<6�>�f%?�4*���߽Z>�1>�z�>~��>}�>����Wy۽V?ܭT?�c��&����>a���7ty���Y=�&>��4�
�R�V>K �<��$n?�����s�<}"W?���>i�)�M���T��UG� �==&�x?G�?��>�ak?��B?���<�X��+�S�Q'�"�v=I�W?� i?`�>R���оy���C�5?��e?[O>�$h�)����.��K�� ?��n?�\?�)��3m}������_t6?g�v?js^��t��m����V��F�>=S�>���>\�9�Pv�>"�>?�#�G�������X4��?X�@���?sO;<���Y�=�C?[�>�O�l>ƾRw�����4�q=�)�>����&lv����D/,���8? ��?���>7�����xx�=�咾�3�?Ӿ�?���9�W;;m��m��O��)�;�o�=�'-��"Z�E쾓�8��̾��	��<����¼�=�>"F@8�ǽI�>V
3���ῗ�Ͽ����%վ2>x���? Ӟ>�Ƚ	ۦ��$h���n���B��iD��){�$�>X�5<�
�>��A�����-�x��<u�N>>ļe�?"v�=D��������;\�>�%2?��?�1�p�P���?(u%�f����ͤ�![�a}:?��?�|�?Lc�?���>W%�(������~�"?�$�? �Z?�eV�&������j?�a���U`�>�4�XGE��U>b"3?�A�>��-�9�|=z>��>�n>"/�,�Ŀ�ٶ�������?]��?�n����>l��?�r+?_i�K7���[����*��E-�\<A?�2>Պ��'�!�G0=�HӒ���
?.~0?�{��.�nk?�op��ݾ02"��
��?��>:�>!�?��+>X�f�[)6�lQ-��?���?m��?Ԭ¾��+�/;?΃n>	g���
Ͼ6P�=�ű>~� ?��l>�[~=���>a-}�ġe�%��>���?��?��>�?���n�����>P��?���>'�?���=�"�> �>�m˾8�e��/+>2W'>Gk����?]�O?b�>�U�=S�/�~����;��vN��x���9�u%p>�i?�K?�4>���G��g)�$���?��F��;9@��8���T���>�X>6'.>#�?���¾��?D����b>��;�Y�j�@?4�d>��>�����ea�����v?�:�>�[�Zh���폿@�E�]��?x�?�P%?���Ӻ^�Z>r�>]?�>�K�N��fp���w>�sM?�\��Í��Xc�x�>���?B�	@�:�?i�z���?�4��ؙ��·�Ĝ�G�<Bv5=_x?�S��?�>-�>�K>pd��9���⃿�m�>�R�?s��?s�?0}?(����\[ >2 �>ϖX?�U�>ygu=���Yզ>�?H�:���kվ�j�?��@��@��(?��Ӊ��K������*���߀=+��=#r"=��F�o	=\��=�1>R�=���=��]>15(>��`>�P�>�>��>����$��]��A�@��/
��Z ��i����s����ᩨ�e2��(���"��W{��v��H��"$�
)�=ָU?~�Q?��o?r� ?k~���>�����y==K#���=\�>�1?L?�*?L��=PV����d�n��~��Җ�����>s�I>7�>�{�>JZ�>��q���H>@>>��>�� >� =��Z��Y=��O>�'�>�F�>�й>Y9<>�>%ϴ�92��A�h��w��̽� �?�}��üJ�2��X8��(����^�=�`.?�x>���?п����3H?����r+��+���>��0?�bW?Ϙ>,����T��3>$����j��`>0 ���l���)�C$Q>�l?Y�f>(^t>��3��Q8�0�P�BK���}>�C6?w���$9�w�u��nH�!7ݾ�gM>F��>m;Q��V��Ė�o��0i���z=қ:?"�?C᳽=����v�۞��\R>�p[>�=�J�=G�K>sjd�k$ǽ��G�a�.=~��=��]>�! ?�.5>[��=U��>��B�a�!��>�*4>�8>�69??�?��?�ʲ���B��Ó4���h>*%�>̬�>(>;�F�z֡=LG�>B�`>_-=�ߓ;������`��*U>5!y�;�Z�������=������=H�=L��g&?��=~�|?�¼�����DԾ��q���3?P\�>��=�L�=�A��%���>d�Z��?��@���?Y�8��i�V�F?��?�����f�^�:>�&?�><��ɾ���>7`!��쟾����<;j��?���?�$V�h0��9'����>�J?�̨�x*�>#ӌ�����1��|�j�	&�=���>.�?D8��?��ok��M#8?��
?�����;Ϳ���� r�>/��? (�?e�l�Ac�� ��jݼ>[��?�6?�?�=eM��쩽:��>�C?&G1?�F�>��#�d����?M�?�y�?��/>�$�?M�d?3��>o<��3�TV���ˏ��-s�H��;�>���g����M�����n�k{J�3
�Ԉ[>G٨<���>]<��Kӵ�;*=��L��L���x�=ǩ�>��;>��U>w��>���>�Ϻ>��7>��Z��vݽ4a��k�����K?���?)���2n�N�<G��=)�^��&?�I4?�k[���Ͼ�ը>�\?l?�[?d�>4��L>��F迿:~��D��<v�K>)4�>�H�>K%��oFK>��Ծ�4D�Up�>�ϗ>����?ھ-��!T��=B�>�e!?���>bҮ=�� ?��#?��j>�(�>�`E��9��J�E�f��>��>�H?��~?m�?�Թ�sZ3�����桿��[��;N>u�x?�U?ʕ>A���҃���lE�E>I���w��?Ctg?'R�(?#2�?�??6�A?1)f>��ؾf����>��!?vj��kA��^&�TG��?�?Z.�>M��-<ؽN ݼVM�����3�?��\?_Z&?��r�`�XR¾�<["���b���;h�S�xs>�>6� ڴ=i>T �=QJm�!]7��7<Dɺ=��>���=�v7�����~%4?�P�<#����V< �h���W��>��3>@��"��?� >,�r�� ��5g��������?pm�?���?� ���\� o?Ui?�q??�Ae?\a���""�"A�����Ͼ�c��/�=ǃ>���<�x�����!��^p���Baн�\?�-�>*�3?���>Ŗj=C <w��9�P�LE�B ��k�����=(��3������o=+�<���1VG��\�>$]½	��>�� ?>P�>��=n�>@�= �4>�>�A>�c�>��>�)>j�;=�9=#u��+�b?H�-�U�X������Q?t�Q?h�F>ͩ[>�.v��M)�U9N?'ȩ?���?�R�>�!��+.��	?�s�>&Ug��Q?.8q=�Ai������h�D�*��1�����~Ls>�8ͽ�C$��W��$��*m?j�?G�>�>ܾp=T�T���V�p=�؄?�<)?`)���Q�S�o��dX��S���(��9j�&���61%���o��ȏ�Jf��@���s|&��U*=h�)?�?�� ��=�c�����k��:@�ib>���>���>���>jC>'1	�e�1�?]�.�%�F+��
�>�|?�!�>��I?�;?�NP?�L?�h�>�}�>������>���;�>r��>`�8?�\-?\�/?�]?�*?:`>_=󽮣���&ؾd�?V�?t�?f?X�?�І�[`ƽ�B��W;����y�=Ƈ���o=�Һ<h�ҽыn�A�P=@�R>k�
?�U^���=�r���M4x>�-?bo?F��>�J�a����_�>X�?/�>���V�~�GS	���?�Qf?rb<�A	���'�>��=e��ND�=�]>���t�=�x�;�|�<S��=���q��=7�=vW�=rI�<[��<��ɽ���>!z?�؊>;��>����?��$�-<�=hL>��O>^�>�Qݾ���������g��4v>�\�?B��?��q=��=�W�=�-�����B��6F��@k�<�?�Z"?�R?*��?
�<?�8"?��>���.J���؄�������?�,?�h�>c��Q�ʾ]騿�z3��?�a?�9a����m8)��s¾��Խ��>�R/��.~�������C�u֌�_��|���?���?��A�s�6����Ř�_J��.�C?�"�>�K�>��>G�)���g�8�p7;>�|�>�Q?�>�O?�8{?i�[?�|T>�8�n/���Й�J�5���!>�@?���?��?y?�a�>u�>�)���F�������ނ��V=wZ>���>�*�>]�>X��=��ǽ2P��n�>�&h�=�{b>H��>���>Q��>|w>=��<."L?�<�>}������-�%%��{+�=��u?J��?ӢM?:;�=�s��>������>�ظ?�"�?0�?���l��=��+>^��f" ����>�E>�V>��v� ?w����>��$?$<�==���~���Y���H��xC?tDB?��ȼ�Kſ�Nq�^r����}'`<c�_�2���7|]���=�����G����t�Y�����Д�Fõ��.����}�!�>)�=q� >���=�'�< 庼r��<&�/=�<~�=j�j���k<�?O��� �V����|�d0b<�TH=�8�!�����?П�>.��>�0n?�L3����=Gk?��">h�,>t�]?��l��R�a���=8�=N�����*);�6ɾ��7��\@�v֔<�kV����=��w>�A�=���)h�=�_=?U�=y~a=ܙ�=�H�=��=�D�=��M=���=���=OAv?����Q��Jj�ZMd���T?j;&>,s$�����
n?�b:>ws������tfl?���?a^�?���>����L�>/U����>��C=>晽��>^�{=���2��>ܡ&>#�!��쮿����?��@�R?ۉ��_�ֿ q�="�2>�>}�O��O/�H�R��Bf�O�L�-.#?!�:��sɾ���>���=�ܾ��¾x�!=��)>ڭT=ce���[��*�=Xj��g=ڹv=��>��G>���=�ǽE~�= -=�<�=Z:N>h킼��9���.��7@=n��=׍`>��>E��>q<?r�6?�sf?7�> �r�	Ҿ]q˾L�~>S��=B�>�Q=|@>��>�1?�C?�P?�h�>g�,=��>�>>�*�6t�yb�Ṯ���<i_�? +�?���><�I=C3@�I��o:�����?'Q3?QG?35�>&��y�ݿ#m��Z1�Т���e=ƭ7=�J��U���@�Ō���Ě�V�=ݥ�>Ί�>H��>^��>��7>��q>�	�>�6)>w�-<܆^=׿�<ʨ�=�N=0��=�伕�M���b6�<�3ﻟK�?e�5m��v
����t���+;�>p��>�WH>�W ?Z�5>��2PU<�o����L�;2�=Nf��6�E�Zgj�n!}����
�Ƚ}ֈ>@��=�]������SN?Jnz>#5�>uY�?�Sd?�%_=n]���ľ����o[̾z�z��P=��>a�H��O��^b��c[����� �>�j�>�>k�u>��*�� <�m^F=+O���5�&�>����bS@�Z0��up�ZG������Dg���'C?������=��?4K?W\�?��>�.����ݾ��)>����.�<o��p�o�JF����?�F&?ޥ�>i��h�D�#�˾�u���ܸ>yrG���O�[����0�b�7��A���+�>tܪ�PѾC�2��J���폿z/B��$p��G�>~O?��?��c�_:��Z�O��&��a���e?�`g?�[�>�?��?.9����쾌1��3M�=�o?���?Z��?Kr	>6��=�[���T�>Q�?飖?
v�??os?i3>���>[6�;� >�^��f��=��>���=���=�?��
?��
?����*�	��p��W�a�^�<#=�{�=��>	�>�ds>lM�=uj=��=�\>$�>��>؄d>'�>�B�>����gm���?�-�=���>��/?3̋>�]�=��ν��<��u��31��3$�ǟ�!罍���e3��<�=�O(����>SĿ;�?{Ee>����?��@7���DT>1�D>Ȫǽ��>�S!>2�q>�G�>�C�>��>.G�>�>5����� >z5�*xD�59 �6f4��+��uH>pQ��>����7��E���j������8�y��`����;�]T�o��?�&�;R��� .��a��<��>���>J�?K[��V�I=�>�%?~��>�6־a���EL��g��G��?K��?Jm1>��>
h?|�I?dǙ��3��6�a�J���h��9q��rT�������g�h�� X����?��Z?�W?94�<�tu>�YX?�*��&���9>N@Q����7>�3|>��ڽ������پ�C
�"E�}�b>o�s?:~?*?����&�[$�>��?T�?؊k?u�?�U.?+�>�?[<=>��7?
�?�6?b(??�>�>��_<p�,�<h�=*�����l���E���f��;ƽ���9�<z�{�=nF
�K�<d��= ���=|�9�><a��<�|�=�'>b�>-�^?�1�>���>U�+?����k4���Ѿ���>��o����@پ�ž�'����<�=?�q�?'i?p#�>��K�'q�"�>��>�ҋ=�{>��>�.�I��R�=���=0h>][#�y��2n���ܾi"��ƞ�<}a�=�*?�^2>`ҭ�<�=*���wC���bj=�Ȕ�q���G����Q�#(���g��>��.?�Z�>�q>����ҁ��}f��3?�u?�<M?]#�?�����w�_H���M��^D����>L��i��N��P���A�D�G9h�g=�>�-������нb>����D�=$n���I��?辁2r=�i���K=�u��tѾ��{����=��
>�ľ�!��d���|��`�K?��=gߩ�RJ�܋��#">���>�&�>���@W���@�����6�=Y��>��4>�������1G��t��~�>��D?!`?e�?�E��Gq�0�B�> ��h����ԼQ�?�C�>��?Ӈ:>�4�=͈�����d��F�_��>�C�>���ҼH�4���Ę���$���>��?G#>S�?�0P?JT?�4a?�D*?�A?���>ZS��<[���?&?L��?t�=�Խ,�T���8��F�f�>��)?d�B���>��?�?<�&?��Q?��?{�>� ��B@����>�W�>��W�Xa��o�_>�J?ԛ�>T?Y?ԃ?-�=>a�5��㢾�ĩ�]W�=�>��2?�3#?��?3��>{X�>�p�=��>��b?Z�?��o?w��=u�?o]2>���>O�=���>h��>��?&O?&�s?��J?Cs�>V�<e��s���t��]��l;!�S<Nn}=����u��R����<؆�;M���_|��S��C�g���.Q�;���>��k>�`���/>6�žE܊��<>R!���[���y���M=�a��=K7�>Ip?�֘>��Y�=,�>�ȿ>�/��s*?6�?��?��<��`���߾�J�>�>?���=M;n�"^����x�M�H=Ll?��Z?=�Y���J�b?��]?Fh��=���þw�b����a�O?1�
?K�G���>��~?b�q?Q��>��e�(:n�+��Db��j��ж=Zr�>LX�K�d��?�>k�7?�N�>M�b>F%�=_u۾�w��q��d?��?�?���?+*>|�n�Y4�KE;�Q���iT?��>(��-�?�$�oپ(F����̾������C�۾h܅�#v���+�������F=�pʼÐ?Ma�?*r?�W?�wݾs�R�|cN�����(PH�dl	�m'���\��=�s
F�y]|�3�����7J���;>��O���)�P�?kg>?�/!����>d���-��� ��ƽ=�����"�镩:^�
�D��D�=�J��;I�:���`8?i�p>H��>i?��`��;�O:��v/����>-��>�>>�n�>�=>����\<S=�a��u4��Ą���s>�qY?��M?Sd?�a��X�"�����/��q���þLe>�����7=�H���Nn�T�-���I���S�$��m/��~��8�;�nJO?0�>��>���?g��>��!���{���������j"<�K�>��?��>��>���/����>}�[?4e!?�0>/��CL��0����Q��ݔ>���=�v�>��i��>�Z��G��)��1�l��̶>��0?��b������WG>
(_?����$i>�>zPн��2��cھQ� ��2>\��>�l0=�jI>W^����Y+�����m7?�+�>BI`�R+)���O���?��?�@�>��?�o�>H��u�=J�?g�N?��]?s?��q>�~�<�i+>28�������g<�er>׫U>�9�=aQv;M?�_P��C�H�<�3�='c2��R���x�<�1�<nWm���=XUc>��ҿ� 3���	��^>����ݷ��勾T�=#+��e����g���н���"a�}9���߂��r�N�w�!�?� �?��վn�˾�ȏ�VKi���Ͼ� ?���.�e�]ݾ����c��	���9�W`)�;IC�d�W�f�]�H�&?N�����ǿ
���e�ܾ��?Z ?�y?� ��8"���8���">�Z�<7��d�������ο�/���^?�O�>�dﾁ������>P5�>}/Z>s&t>g��]���ѕ<n�?D�-?���>�r�Z�ɿ�K��KϬ<���?�@WlA?��(���%�S=H��>F�	?�?>��0��R��>��w>�>\>�?Uڊ?��N=�uW���	��@e?��<KG��ջ,��=_�=7�=�*�p�J>�`�>"��'A���ܽ}�3>���>��%�xV��>_��\�<}q]>BIԽ�u���؄?@�\�Y�e���/��`��a>��T?�#�>��=��,?�>H��fϿ��\��a?�&�?��?��(?����A��>!�ܾ�mM?�.6?��>6c&�߲t��I�=�߼ZD��!���V��Y�=��>�>��,���FO��������=�����ÿ��$����-�<����Un�R���3۠��4���7��s�V�����!�9=vr�=��6>fj�>uaS>��h>4\?t�m?�>d�2=��Ż=��@���E\=x���Fq��9���-��m��3 �+%;��	���>-�W�;jS@��n�=�$U�}m�����2Z�K�C��Q0?tv >!�Ⱦ�aG�tI=S��� ��#hq���轥~Ͼ�-��k����?��F?d��^JQ�y��挽W����W?���K�Yг���=�z�u=���>N
V=<���2��Q���*?�?a
������e�+>�n�ΥI=m�*?�)�>8�_<��>��&?d�&��+Ž>4_>^�->+ �>B�>z>`��`=���!?�T?I�h�����>'���3w�lv=�%>��2�����fe>��}�9�����<�`O��g�< +W?a��>R�)����Sn��l���==��x?%�?=N�>~k?
�B?�K�<�f����S�4��!x=��W?'i?ޢ>'*��о�|��]�5?E�e?��N>qoh�y���.�eP�?��n?~^?�]��e~}�%�����el6?�	u?��a����J`�~�X�K?�>��>���>�3�w�>�G?��R����s޾�-�9��B�?B�@���?1z��� <�@b�}^?��>�W�1儾���Î���7�=}�?� ��'���I'��n��PN?!��?���>���������=�ԕ��W�?��?�{��5�g<��?l��u��[О<��=��;�"�B����7���ƾ��
�����z��գ�>:Z@�.��E�>N38�c1�HOϿD��n\о�]q�<�?]^�>��Ƚ❣�l�j��Fu���G�-�H�ꃌ�SC�>�*;yUl>��+��s��[��eܽ1d->9>���R�>�"�N�Gȩ����=���>�j&?'��>=ʾ @־鶜?��6�_�ɿ�D����8���%?ǿ�?�^�?RQ�?zAs>U����W0��~�=��T?�̅?�g�?�,}��c\�k��=%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�d�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.��xp?6�~��d<���'�l)��6�>4c����`���D>R�w��o�+N����x��?�!�?c��?|�.���=�N�0?XE�>l�׾g�����M=Sk���H<.�>�>u��>>VC��*���N�>�[�?Y��?X�?Z���kh��K"�>���?Bж>u�?���=PB�>�9�=N���8@3���$>��=ڌ>���?��M?�3�>"�=w�8���.�(F��7R�_��Y�C����>�a?rL?{�b>����:�5�!��ͽ?Y1�}M�L'@�ކ-��T��4>V�=>��>$�D�x�ҾS?�4�/�ܿ7\��[�X�G^3?��>���>TD���l���o�Zlw?���>*3����ُ��1J��oѭ?y��?n�!?�J	���<~�=BB�>��><�Ȥ轤���h4>�mS?�✽
x���u�^�\>u�?�.@M�?A�h�{Q
?�g�oȑ��(���V�Wu>=��=ȿ)?����-M>��?[L�>$a��yĪ������f�>o<�?0�?'6?��~?֋����Ǫo��?�>���?�ݡ>� -�E��!�S>��&?������-���s?Z�@u@�IL?����1ݿ�E��"���e���
�=U��=� �=�8=G��=+�%>K�=2��=���>7k�>�	>E��=�f�>\4>%(�<�����nqԿ�w�H������zk������.�����������ݸ���:��VؽV��L-��`�ƽ(�=�xU?`�N?��l?�a ?��]�޺$>24����=���B�=ת�>��0?�K?��(?��=ኙ�_Ce���~�%>���]��GE�>��J><H�>+
�>z��>�!�<3yF>�=D>/�>�%>�*=إg<�;�<T�J>t��>)��>�
�>�9>Um>�ߴ�����h���z��̽��?�V��M;J��ڕ������ʶ�뼟=� .?���=` ����Ͽ�譿7�H?�����G���(�ˑ>�]/??�W?�P>����\L���>��O�i��%>h����l��)��Q>g)?��a>��>K�7��~=��s:�����]l>��,?�7Ѿ9Hj�2q���K�1�ɾ<}V>���>�����(��:���,���z���d=�+?g?��8§��kb�#o��.l>�`h> �=���=�z:>����BX�ZhP�<-m=�x�=">�?.�0>���=���>�C���TP�Σ�>'\B>�->҇>?�#?g���N���ł��+���x>si�>��}>,	>�OK�t�=`�>��]>���d���
��"9���U>,�x���Y�R�n�;Eu=�T��g��=�W�=�N���#;�M�=��}?C��d{��H	�����IA?:�8?_�>��!�0�D�	h��|�̾ˑ�?	�@~�?yB7�-�Z�2�8? �?�/�h�'>J?��>�p/��	���<F?w
���Rq�s`#�� ��Ӱ?W&�?��=�S����r��Т=|�J?�����>B��/ޤ�]����iv��4z:���>2�F?^���%O;�B�f��_&?�_	?��hO��=̿�s���>~;�?3P�?=t��r����9�B8�>��?O;F?U�>_ھ��b�9+�>�O?�q5?Qu}>lU4�����B5?u�?�L�?*K>�o�?[�x?>p�>�&;�A��ݯ��^��orQ=)ZO�x�>��<qE˾��E�*◿�Ņ�Xt�T���7>�	=哜>�����F���X=_g	�r�����Q �>��T>�?F>�W�>/�>+ռ> �p>��<P� ������J?n;�?����`n����<�=�3^���?]u1?$�] Ͼ>�)\?|��?�>[?ZG�>���1ך�d[������l<�|J>R7�>��>Cۊ�wH>�Ͼ#x>��>>�>`�n�پ,q}�BU�:�ќ>Ȋ!?��>^��=J� ?S�#?1�j>�(�>�^E�I9��a�E�˱�>ա�>�H?��~?��?.ع��[3�;��桿��[��6N>�x?�S?�ɕ>����ă��Q^E��\I�c�C��?�sg?]�?�1�?Y�??��A?�*f>���ؾg�����>	9=?�<��3<��T��1��љ?��"?9-�>:�>��Ͻ$cξ���Hؠ��Q?}�x?��?4+#��B�|�]=y*[=ؙ�=gρ=N�*>}Z�=�>�ӆ=�q��Q���	�>��>]�Q��链���<��W=LEW>��>H{s�@�5��B8?v�ڼ@m�6��=*�y�G�;��1�>�2'>,ak�mτ?�R���t�]�������졾4�?��?���?�S?�{Ae�q�S?�no?y�?��?���-v�?T��ｾ�BZ��W��w��=���>O5�<j;�R��?ب��Wm��f��c�����?�I?�A??��I>o5��yf�#�6���ھw�6�c:-���S�sgb����_y$��ᾍ!������¾����j�>ѫ��Mog>R��>�ׄ>%Ǹ>�ê>d���e>�F�>��W>C
>�K>�e>�);>��S�/;�@xS?]4����b+�����K?BGq?jW>�=��̇�E���	;?oͰ?3T�?w֬>[cS�du!����>��>���'>?�^�<���鬛>����QM� 6�������n>@Da==�y�R����-�>��D?h�}��T�����}��'{o=dO�? �(?�)���Q�r�o��W��S�f �E;h�
���j�$�˛p��폿V[��[%��9�(��0*=��*?��?��͊��$���k�5?��bf>c��>�>ݾ>�oI>B�	�ɵ1�R�]�_B'�����\7�>�N{?�p�>P�I?��:?��N?K?@�>�X�>�������>��=;�p�>r%�>��7?x_,?�g.?p?%'+?��^>������J־bC?Pb?x*?^$�>J:?�*��;S��{Ib���׻�v�������=�B�<~�ֽ/9]�y�_=�P>�J?lF�I�8�O����k>�x7?]t�>���>���-�����<�
�>ȫ
?z>�>�����hr��Q��5�>@��?��Q=��)>+��=�W����꺊%�=//�����=�O��M�:�ͳ <���=^{�=h�|�j����k;&�;���<2�>9(?�޻>�5	>-ɹ�f�6�w�޾p���<<>��7=�">���ݎ��[���5l�ke8>)t?���?t�ļ=��=.5$=�j�&ʾ����콾��ԽQN?m�%?�D?�{?.?�?\��=�i(�uҋ�������f��d�>�T+?^�>���B;����# 1��]?�?�<a���Ik'��ߺ�,7��>��*�~1|��X����?�&���W��IR��?�:�?��W�7�3��:侜ę��C��=@?���>9o�>y��>
+�> i��k��:>��>&�Q?
"�>��O?M:{??�[?mT>O�8��.��;ҙ��3���!>�@?0��?��?Ry?qq�>�>��)�n��K��A��.��݂��W=�Z>��>1-�>��>��=��ǽ�N����>��h�=P�b>t��>K��>�>w>�]�<��_?�K|>1��um�����to�8c>äQ?�>�?�X?9o+=,(�"�%��K�r�>qȶ?X�?in�>�̽GA�=j��=��]��q�� �>k�H>��p>cy'=>�w���?R!?�V>m	3��,3u����фA?=A>?������ۿ�承;\6��">6�齅8���i���[.�Bf0=�(�>�S>
>>jE�����^����X��[�����c��>oF�=���>��=��~=���<z!�=���ɰ�+Օ�&WŽ�;ۯ������ټ�Z%=
�{�<�t�<��h�y�?��>ں?d�z?�"�="�j�E��>u�>���=n�? R$>��)�چ��ýG*��bD���Ѱ��Zj�IT�DB�<2F�<m��=F>>��>�%��2+< ��=Yp�=܄��w<>��j>��3=f��;>�=���=���=�+v?�9���H��	�x���9��؛?Ӷ<�/=껬��8?��>��^� �������r?�5�?Pi�?�w�> �H`�>�跾�'�=�_f>#1|=��<үF;�g�}��>��l>H�0����� �j>���?Q6@��3?|[����翇�a>i�/>7>��V��?��h���:d���m�$"?�H�j����
�>�=0���H'o���P>�U�=P^���� �V_}��==�<��%>���=�>Z�=>��=�`�<X >��{=�R>>�t�>U���8�;h!=Y��=�>�I�>M�>R�>�?LT0?-=d?j�>sp��p;~����J�>ۿ=4�>��}=�>>2C�>"7?�D?��K?�ʴ>W#�=:J�>mK�>�Z+�'~m�x����9�<
�?sd�?�5�>I+�<�@�����=���Ľ��?d�0?��?���>���ŕͿ!�5�a��"������^����7/<�3P>#��=�F�=x��>��r>��>��/>��>"�,>��=��>���=�%�=�kF�m
J<����küo"x��]�����=i��N�����<�*$��U�vP)�1톽ѧ<u�>��>� ?ҟg>���>��=$����>b����u�H(�>faX��a�k�D�d4X��^=���P���X>�l=]�=1\��~,?8��=�>�g�?�$j?̬�#���i\���Q����g�QC������<�)�i�w�x^H�MJ��+��>4*�>;j�>l�k>�'+���>�Wub=I&��n5��c�>�ԋ�50�����q��S��Ȩ����i�����gC?I���w��=IY|?֪J?Gb�?��>�����ؾ�)>�j��� =&���s������?3�%?���>.;�6�D���ʾU:����>G�B�coO����V0��$��=-��P¯>h{��Y-Ѿ�3��4���֏�D�A��8p�
 �>sN?�C�?��f�/ڀ��P�?J�cx��'�?_�f?7ޟ>�?�O?[����꾒}y���=|�o?���?0��?$�>&�=�����D�>�?#�?��?9)q?��9����>!�*<�$>�i��|,�=r�>���=PY�=K�?�?�	?�䞽��C�쾩��!k�,�<��=�I�>�=�>G�q>7��=Ct=Xѧ=<k>�N�>�*�>��k>I��>��>�܈���?���<��>�|?"�9>���=!�>����&�z~r��9�̻SH=t�<%�k��ƞ=rA0�w�>��ÿf��?�ij>�a�j?�Ծԫ�9�X>�x7>���B�>��=�Z@>j��>��>x->�=�>9c9>�۾��;>�(2�f~.��.G�z�d�����o(�>����C@�;b�-���1����b ��y��W�A��V��)��?�9~�K�r��	�q<���>�q�>3�?��I���ʼ��=­?$#�>�����6���ɾN2�?~!�?��z>W׸>��M?�=?����.���L�Ҁ��&yN�n~��c�sX��9Q�����9���,A?y(a?Y{^?E��=�`>���?>�B�����g>��4�����zL=D�>M ��"{O����C�s�����I >��`?�?ٚ?<�*<������?�8?�?#�+?��>gfL?�t�>c�?��>�?���>�V?WH?H��>Y>���>6�p����=�Oo��;?����\&�JH���U=q��<��K��n=�J�;؂=c�<D=��m�9μ��`=�ቻ�=Wc�=��>��l?q�?'s�>�E1?Il;�mҾ�����>򦪾ЅY�>˾p=Ͼ��۾��=��<?�&�?�C�?�C�>�,O�'\�	C>�\����>q'�BX�>ۄ�dTҼ1X%>�dq>�R =��b� n��8�����JG��$,�=����>�0L>�⽧o�������m��=�Λ�.S�ξ�J�F����ۺ�Gx�>�F?��?�������֮p��
n���C?�n�>��M?3��?��=;Ež�O��^C�s���ir>K��y�3�`����/����/�����)5N>�鮾Q����!`>+�����l�wdJ� ���b~�=+��(�{= [�a�̾-�n�k��=��>�Pľ�_��N������hJ?舆=�R���A����?�=w�>��>�X�K^�)�B�􆫾�q�=�w�>��->����\�fL�b���f9�>�LE?�T_?�k�?x���r���B�\����p���,ɼ/�?dp�>�R?��A>���=������x�d��G��	�>�t�>���`�G�8��� ���$����>3?j >��? �R?{�
?q�`?�*?NM?�.�>~�����?&?}��?���=X�Խ͹T���8�<F���>2�)?�B�Y��>=�?x�?K�&?�Q?Ĵ?S�>0� ��C@�h��>�Z�>u�W��a����_>ԪJ?M��>,@Y?�Ӄ?K�=>ń5��뢾�ȩ�]g�=�>s�2?�4#?g�?��>��>����y�=}��>�
c?�+�?�o?���=Y�?�]2>��>��=y��>�}�>3?�PO?z�s?��J?��>��<~&���N����s�F�P��:�;^H<y=׭��Nt���� n�</�;Ł��:��V^���D�x���4�;�;�>�g_>�W��cE;>�Lɾ =���@H>b�䷾iD���	����=/f|>�3?���>:�6��c�=�/�>���>���J/6?�?�]?ւ�<�_���Ѿ���٬�>�8?��=�8g�H���b�}��~�<@�l?�[?�d�8�׾K�b?��]?Dh��=���þ��b����d�O?5�
?;�G���>��~?e�q?W��>�e�,:n�*���Cb�
�j�Ѷ=Tr�>JX�Q�d��?�>m�7?�N�>/�b>"%�=cu۾�w��q��g?��?�?���?+*>��n�Y4�	Ӿ����(�G?���>��p�d?t=<�P;�S����߾�y����˨�j���L����n�����]�G=�
=tc?���?��`?5|?�!���p���B�4=��0�W�ض��(��zM���9�<�=�
�c�����þlA�dB�>u�b�]�5���?k�3?H��y?x���;�	4�,��=I�����t�=>���Re���9=�i2�Z�1��˸*?�d�>	��>��*?�"_�N9�8'���0����3��>���>N��>�>����;0�C�ȼ״���,���N���r>�Jb?�L?��p?���0�r����!���`��x���?>���=���>M�g���(��&���?�|ko�����=��C��N/�=oZ2?(��>¤>~��?Q�?���<��B�x�+'/�P�<�η>��g?���>�T�><ݽ � ���>��T?�x#?��>�&�m�k��"��+X���s�>��H>��?��Ͻߏ�Zml��1��#铿ª?��>޿2?ǆ�4	����>��?`ƕ��̔>���>��<6�L����X$���0=��>��u=�ʒ>x��+�޾��~�����r+?J?ϻ���(��b>��"?�^�>p�>4�? p�>7�̾+g���?��]?i�M?"5D?���>'��<�7t�ֹ�����y�<c݆>�tk>W[�="�=cF�,Id�/���p=:�=p������N�i<K����D�<Z �<X7>�a����B�����,L�,.澩4k�hE�Τ����ž��1����۷:��Ј9�B������co��\x��D���?dX�?���V�NN~�
�k�����lZ�>B7���������1��K5��߾]x�����8���Y�0z8�N�'?�����ǿ񰡿�:ܾ5! ?�A ?5�y?��9�"���8�� >]C�<�,����뾬����ο9�����^?���>��/��v��>ܥ�>
�X>�Hq>����螾�0�<��?1�-?	��>Ďr�/�ɿa����¤<���?0�@KA?��(����0dS=���>�	?�"?>�H1��@�Y����>;�?؊?3�R=>qW�I�|Ce?k�<IG�P�̻��=��=�+=[��mK>!f�>:����@�PB߽T�3>��>+/&�W��T�^�\�<�H]>ϕҽ���b�?E]���b���-��$���X>��R?5�>���=��.?� F���ͿI�\�չ^??�?�?�%(?m�ƾ���>��ܾ��J?�-4?P�>�G'�_1t��n�=}ܼ(�;�ݾІS����=L��>��>�-������I��������=�������pa-�S'1�~�E<�=��>	�����!����u?-��-����=�=��4>` u>jta>˂M>��W?*�l? ��>�I)>pV�r���Y��<�M��%��t���8�$q��0pᾄ�۾���ر�[���ξ&bM�yi=��X�]���S���W�YE���-?�>���f�D��]=iĮ�쁮��fּ��ὕ>̾X�/��Wg�f�?�@?�
����N��	��=��&#��V?W��t?���������=s�L�H?�<8��>��y=���r�3�
F��o0?�X?<���@\��V5*>2� ��=�+?W�?):Z<�"�>^E%?��*���(`[>��3>�ң>��>�	>����S۽�?��T?$������]Ԑ>\����z���`=�6>(,5� ���[>�2�<�=V�J'��Ne�<�)W?���>B�)�j��i��0���c==H�x?!�?"3�>�yk?$�B?wä<:i����S���sw=�W?�'i?��>�r���
о�|��9�5?��e?��N>h^h� ��:�.��T�"?��n?�^?MН�x}���T���m6?��v?s^�xs�����I�V�i=�>�[�>���>��9��k�>�>?�#��G������}Y4�#Þ?��@���?��;<����=�;?l\�>�O��>ƾ {������Z�q=�"�>����ev�����Q,�k�8?ߠ�?���>���é�3��=BՕ�Q�?K�?(k�� f<����l�{�����<Mh�=��;�"�����7���ƾa�
��u��@M��⠆>�Y@�5��S�>�_8�N6�|IϿ���7rоi�q�;�?`a�>ʚȽX����j��?u�{�G���H�6Q����??f�:�j�>�{ؽ{*{�sT澱(>�M>mj=��>}?<�P仾9���n�v߰>�@0?�?IdI�����?��:�]ҿ���[Xi��`�>%��?��?���?��>p�y��|�J�K?���?݀?�����˖�Y|>��j?yb���U`�E�4��HE��U>n#3?ND�>%�-��|=q>��>�q>m!/��Ŀ�ٶ�������?���?=o���>���?zr+?�i��7��$Y����*���,��<A?�2>���^�!� 0=�uђ�ȼ
?�}0?�|��.��p?���f]6�J���6�.Po>��@>�=T8?��=����y�
��qz�?�k�?ul�?7����6���R?$�d>@̾d
�z�ȼ�U8>L7�>���=��<��K>^Pf�/B����=	��?F��?�!�>v.��u��Lu�=��{?�G�>�?l]�=2��>n>]������`>ge�=�A���>ڮK?�l�>��=�O7��Y,�J�H�NS� a
���E�Ժ�>y�^?��E?�s>S��$�3�;}�Vӽr� �a-W�
;��K��Tν+�4>�d<>h{#>�
7� �Ծ��?B���ؿ����(��4?�)�>o<?G��Փs�u��ɕ_?�g�>���D��y(����|�?q{�?��	?�ؾ�YӼ&>��>���>�ս���������7>��B?�A�'h����o��A�>�	�?��@C,�?�h�`Y?�1	�l���EQ�������\�C�)���0?4�ܾې�>��?[�Y>�x�^#��3��贩>s��?Rk�?�r?˭�?�Q���H���>y��>��u?�f�>�$��ݵ�r�>Gr?�?L�������?�@�	@�9[?s����hֿ����fN��o���"��=���=v�2>��ٽ^�=��7=��8��9��X��=@�>��d>�q>�'O>a;>ٓ)>���%�!�%r��n���:�C������Z�>��0Xv�:z��3������%@��3ýjy��	Q�42&�>`��J�=�W?�?I?\�k?�	?�8��B�=�ؾ��=��񽼢�=��y>�U ?;??�&?#��=�����f��{������?���E�>l6Z>���>���>�X�>���<��>�B/>���>!@m>t�=v���Wh==�]>ab�>��>�-�>�<>�>�ϴ��1��՘h�#)w�Rv̽T �?���B�J��0��A-������tF�=�Z.?�c>k���=пp�8H?����.�l�+���>�0?�aW?��>��p�T��>a��Κj�Ad>> �:�l��)��Q>@t?�'e>�ls>��3�r�7��N�X���ν}>Av5?�+��+�;�Awu��oG�ڤھj)P>rB�>N������"���F��k���h=��9?P?���|����z��D��B�Q>ܔ\>�)*=���=��L>��X�ѿ��D�-Q7=~��=Y�X>tO?�+>3�=H�>�'��t*Q�0�>+-A>\�+>��??�'%?5��?������Ds.�)�v>��>)i�>]>��J��P�=\@�>��a>�A��M��] ?�!W>�}��_�2w�-�y=����D�=��=~y���;���&=��v?ÿK���c�7տ�"�U?B-?�/�>�@=��d�����a㼾�Z�?q�@�?�)R��c��U?4�?�G*�%��=�>d�>�P��F��lH8?;��=2�����U㽒5�?KB�?N$5�{n��V3���U���D?25���D�>oK�e秿o���Z<o���<��>T\?�?���=c:`���.?��?g$۾ꔩ��mĿ,�m�ol�>���?���?��w�歙�n�<�c�>���?�pK?���=x춾�<�|�>��7?�.?ʊ�>��2�1D���C?���?B��?L�=>�E�?�n?$D�>�yǼaL��K��d���pp�=��幜��>�8
=_z̾*�L�J���艿�^j�> 辑B>F��<æ>`���������=��8�VfϾ��}�T$�>�
Y>�u4>hB�>U� ?Qf�>�Ї>�ռ�y�]n��*y��o�K?���?2���2n��Q�<w��= �^��&?^I4?qn[���Ͼ�ը>�\?g?�[?�c�>G��B>��D迿C~��X��<��K>�3�>�H�>�$��(FK>��Ծ�4D�gp�>З>����?ھ�,���K��ZB�>�e!?���>�Ѯ=ҙ ?��#?��j>�(�>/aE��9��Z�E����>ڢ�>�H?�~?��?�Թ��Z3�����桿��[��;N>��x?V?gʕ>R���惝�5lE�BI�����T��?�tg?cS�$?92�?�??V�A?N)f>��<ؾ}�����>B�D?|$���w-�Y��7@��b�?7��>�J�>�8�>��u��>����M��5�?�k�?�GS?�����s����إJ=�̥=�h�0�=> >Q[�=ݟ��@-�g>>��,�>T>�7����¾Se���=y��>hÐ>z���@3��=?ߡ�tXW�{C+=�y� 0���>>w�>,Q��kq?aU��Kn� W���+���Bc�8�?���?I
�?���2�j��P?��t?�'#?��?����/���q���t�ƾ����+]�h=�=�D�>WXH;Ί���������k�
�B����:?�?�G?�?j�g>G>� ��3g7��~��$���E��P�~�;��h)��
��z��dS�����-�ȾQk�$[o>)�ս4��>��!?s�a>�h�=W�]>4Y���>��>f�>��Y>)�K>��>�x�>�ͽ �� (S?��"���)�kI���0��=?i�?vY�>}q��+���Sj��'+?�L�?}�?�՜>�����`-���)?��>�;i��TO?/�>����<T=_X*���WHо)��)�>�-���X���5�̾M`?:�.?@�=���u\������1o=�L�?��(?F�)�d�Q�&�o�r�W�#S�����)h�mu��4�$�H�p��.^���#��F�(�[*=F�*?,�?(��5�����#k�{?�vVf>�	�>�#�>#پ>xI>��	�[�1� ^�dN'����M�>�W{?ī�>��I?;?R�O?�L?��>���>�,��D�>��D<�ޣ>��>��8?9-?�6/?*?�*?i]>i��9H��,�ؾ(C?�?�_?�� ?��>h��[羽�q�`��nq�n�w��Ut=���<�Iؽ� t� ,K=3�S>�V?I����8�������j>g~7?�~�>I��>���}7��#��<��>��
?�T�>����r�{c�]�>W��?���0m=S�)>���=
���f9к�[�=�¼m�=:Y���h;���<�f�=��=�s��j��*�:���;@�<
��>2�#?e=�>"#�=A�ͽ��P�-��s�4��\F=��<�Ҁ>ָ��+��׌��x�d�>��?�޺?��Z2��6 >01=��Tھ�➾�?���;�7��>��D?LiX?@|~?r�>�?z�`�xW2�w�������A�!�>P!,?⊑>�����ʾ����3�ǝ?;[?�<a�q���;)�֐¾>�Խ�>�[/�a/~�����D�E����������?���?�A�$�6�Iy辷����[��Y�C?"�>`Y�>[�>�)�<�g�I%��1;>���>
R?�"�>��O?G;{?*�[?WfT>Н8�^0���ә��3���!>�@?���?��?<y?�r�>��>�)�c�hP�����n��݂���V=Z>
��>�)�>t�>��=��ǽJT��i�>��U�=��b>o��>��>x�>�w>�2�<�ub?��>�f��B��n��.t_���O�M�5?h{�?�E?��>>Ws��U\�qD�ٍ�>��?v�?bv�>����<=��>�rB���|��=�>૙>�s�>?��:I
��ˁ>;��>W�>7��%\3���^�}�R���&?��i?����s�˿
0g��3��0����\)�v�1�
�	�}����=�4=�t�=,�L�?Fm��t���
��P<���hh���i�ƞ?��>�b�=���=}(';7�޽��?�M��=N�<Mh�<p���x���>���GF;�|���M\;է =�2�=����;�ؾ�I|?�?o�"?��g?h>�,���D�>vO�>� �>�O?{6>wg2��w���w����=t*����K�о�K��sL�\�2<���#�b�3=rB>�/�=���=5Y=?�=>��<�Y�=�:>u�d=��Q=���=���=.e%> Vw?����Q��-`������4M?���=�١=�d��[7?aq.>�k�� %��o��2�u?��?��?�y?~�t��?�>���`�=��>@#�*�=8�1>�����>�
�<,}5��㮿g�=�'�?c#@�X%?�v����ӿbvO>mA'>'ى=ԣK��,����]�a���U�.�?��=�ܾۚ��f>'��=cZ���-�����=�P�=�@�<��� �m�뜛=���/5>̖�=Ou>9s>a�t=��̽��=q�G�AB�=V�4>P�>��&ɼ�D��J=�n�=)ۇ>�p.>��>�?'10?��c?��>Y�r�;�nƾ�y�>�#�=��>G�z=�>>*Ѷ>�}6?�
D?XM?��>�=a�>�ץ>��+�s�n����料���<]��?�C�?@��>cC�<��B�<?���>��'Ž�?>k0?��?��>�U�j�࿘Y&�]�.����DW��+=�lr��[U�5����k�P���=�o�>_��>4�>Sy>��9>w�N>L�>�>
:�<�p�= 댻��<���J��=ۗ��q�<Lzż�
��ʳ&�}�+�'���d�;0��;��]<3��;��v>��>�/�=J�>N�*=�ۙ��&�=D���;��B�=&�ƾ�4F�H�Q��TW���#� `c���R<d�=�qȽ������*?X6�=Ơ�>��?�YO?3���b����̾�њ��!�����8�<�4�=T�5��E1�=Q~�J>M���þۣ�>�Ŏ>?��>Gm>̋+�� ?��y=���W�5��	�>����`B"�����p�?���柿+i�ҕ��D?�N���{�=n�}?�I?��?˝�>2<����׾�6/>hD��'"=��_Xp�� ����?v�&?��>�?��D���˾BҾ�n��>q�G���O��m��j0�E�?��L���.�>	媾[kо*�2�ij��J���6AB���p����>�QO?�	�?�pc�$=��4�O��#�6t��ME?3ug?���>�?5�?U���`M�������=�#o?���?��?��
>@?�=�g��!�>�1	?���?���?��r?�>��z�>)p�;�� >М�� �=C�>,�=�Q�=b(?S�	?�U
?������	�b��O�$^��t�<���=�>Ț�>�Kq>��=��a=ef�=��\>�ݞ>=�>lUc>tĢ>���>]�������D?�|�=֥�>"�?��W>��y����eXν�M����mb�����7����'�u�<���=⇾��>�O��6�?���=%8�S0)?�������۰�>�n>mp$=�k�>���=��{>h��>��>B�p>-l�>��=�)���>�p-���<��i8�=vX��*����>��������q���(<�Ԍ�W������j�S[��IxH��b=���?K�Ž� ��_)�y#��?���>�m8?����p�B���=7
?�s>��ʾ]P��i<�������?��?!h>��>	�9?�?V[��:��<�1�?h��q�]�gl����v�Y���%\f�$̾��޽U2?Oރ?�"U?z>��+>�}o?�x���s��W}'>�%����D���f>'UO����Xľ��Ͼ)P����=��c?�er?��>�9:�ʙ��t��>-?`�?%j?
��>�?q�=��?Ů>P�J?��6?�^?�~�>�X�>|^g>�|*>�C�&�%=�T���r��=�%�V���v��=Il��s1.�ęS����=�9�=�#� 𺓿�=�|�+-�w��=�*�=&AR=�W�>�oX?2[�>u�>�z'?G�p��&�?.�m}	?��$碾*I��2���4�\��=�p]?0��?�^?�(�>��B��y,���>��>^\->�kG>\s�>�S˽Y�"����=;�H>)�=If5<��V�����o3���P�<bM�=��?�">!yٽF�=�p��EH��㞎>�Zp��oľ/�v�A�>���#�a�U��`�>�kG?7�
?�P�=]#Ǿe6����o��z??ў?*iJ?��?Ov�=~��a��WR���ٽ�,�>���16��㦿�H���S.��� �I>>w�� ����t]>JP�����tz���?���ž �=�R��M�=b��e���̀���=�L#>a���6��qJ��'|��(G?�s=���B 4�̶���>K��>�7�>���Đ�nGF�'���,=� �>�E;>p��C*��J�2���>nW@?��e?� �?�v���#�V��V��>G�����8<?��C>[�%?82==܎�=u����;��l�R_��?D��>"�7��)D����M_�����ޡ>k�7?s��>���>QNm?f>?��p?|�H?�O?+q�>�?�:���t1?`ƅ?bU=����ib���_I��K���?��]?{�<V8>��?��G?�"?��[?0�?^�n>ӥ�:>H�]��>��>,-c��(ǿ-$3>���?���>�`?�͝?u��>�8�4X��T4���}T>�I<��>?�J?]8?�o�>��>�!�����=.�>+Z?N��?�b?P��=�< ?��>��>z�I="r�>Ĝ�>t�?��J?�q?E?]��>ìE<�᤽!e�K��c�;7�+<�
9�%o=���.���bKM��=.#�<{lj�Sּk����⡽b�̼�:��7R�>�s>!����0>b�ľ�I���@>��[��+Ί��a:��=L��>��?���>�R#�
��=ݯ�>�1�>���Z1(?�?!?h�;�b���ھ��K�w�>�B?���=A�l�|���-�u�\h=�m?��^?��W�W.��=�b?�]?h��=���þ<�b����/�O?6�
?)�G���>��~?G�q?��>��e�6:n�-��Db��j��ж=r�>3X�	�d��?�>>�7?@N�> �b>6%�=�u۾�w��q��t?a�?�?���?g+*>��n�P4�3�ᾬ!���|j?�;�>b���~�&?�[��*þ_���m��fḾ�׷�����m��R�������;U��~���n=zw?��{?��d?�q[?��ȾW�\���O�l���jQ�/~�0W��i0���B��I���r�< �x!�!����|�<��{�Q�C�ʌ�?�'?�V/�)�>���^��t�ʾ�[;>�Ӛ����F�=�璽W�G=swd=W�`��"+�l���0�?�w�>2��>,}<?Q�X��Q<�@�0�v�6�����U*>��>���>�*�>6����i/�k���`̾�X����ؽ�^>��Z?oP?�G�?F5O>��-�˨���HF���&�ST3��]X=��y>��ھ,9}�o�/���?�#E��PS�#l������s>�L?���=/��=��?OA?����κ����&
O�ퟢ=1�|>f�r?$�>m>�ɳ<}ha���>�$y?�"�>@DX>�Pg����g�����~���>tj�>�=�>��>Q*��P��'��"��WU�g��C��?V�n�4r����>��i?�R=���A=҃�>vp��47�:^���BF>d?�M��a�u>��X�����������ކ)?<4?�f���T��B�>�???�>ɕ?���?�>\Yp�$A>��;?��h?&�)?<�H?�P?�X>��ؽ��"�$/��k>'�j>	�Q>=�<�>��{࠾�U>���>�[.>��۽j:��p;=�5�Dν�	�=y�_>r�ܿB�K�SɾԒ�tJ�a,	��1��Q�����8���Y�"4��S(�`{Z��=6�'��|z��0���f��B.�?�n�?�1��%4���P���ww��7��:?�II��������h~̽+���\ƾ/����<���I��m\���a�Ӫ2?�"���"ӿp�����׾��8?v"U?��p?ý�m;/��XS�\��>���=��=��־�t��d�ǿ����.�i?�/?���z�Y��>䘱>�>�>�=����;QIA=k�?4�)?:�>n�iҿ]��
��=���?p@�uA?��(����~V=���>n�	?��?>Xm1��C�~����W�>�6�?��?��M=C�W���	�D{e?�<��F�#4⻄��=�`�=�E=Ǳ�l�J>�;�>�b�{2A�c7ܽr'5>j��>�Q"�Έ���^����<H]>b%ֽ�_��5Մ?�z\��f�o�/��T���T>��T?�(�>%+�=C�,?�5H�<~ϿǱ\�'a?E0�?w��?@�(?�ֿ��ؚ>��ܾ��M?eE6?K��>
e&�T�t�π�=�U�TH����(V����=ҩ�>A�>�|,�C��}�O�-p��Y��=XQ��+Ŀ����m�	�=׃�;��c�vw��������"����Ke�ջ���t�=N>4hT>��z>�o[>޶J>�lY?��q?��>���=0(�k����\��SL�=�^�eb!��ƍ�4p��ة��v侊bӾ a	�1�����Q+�-M��W=>
G��o����,��^��$���8?�^�=no�v�F�]A�<>���-�N�'Cc=�߂�e�̾Y�#�n�g���?�G?�q��P�T�5�f�<2ɞ���`?P�E� ;s�%��>���q?v��a>�=�Ǿ���iXE��*??�0?�x����F�=���{��<�)@?�*?�$>s ?*K9?��tTu=�o�>�b�>��>�-�>@��=_����5��2?�i?�Qs���˾���>"�ľ�n��-
<�G>�#޽�.�a5�=` >���hϖ����<v=�'W?��>%�)���cb�����|e==��x?��?.0�>yxk?�B?n�<rd��^�S����sw=��W?Y'i?��>�����	о>�����5?��e?�N>�_h�5��P�.��S�$?��n?�^?��u}�	������o6?�?n\�Gʣ�D˾k�+��`?��>-�>܋N��`�>��6?����}���ɿk:�MT�?7�@��?L�=�ϛ�G�'>�,?(۰>쑮�U�e��>.���Ƒ�8�?��P�������G�s|����t?���?;�? ����c	�pu�=���̥�?�L�?�_Z�u�=Z^�W�j�T^�������=6z���ڽ���ݜ<�-C۾o���������l^>�@����-�>Ăi��ٿ����4��ؾ� ��M�>��>
Fy�o����t�|�6�W��@�ڂ"��Ԣ>��>[���DǑ�,"|��:��(�����>q���>o�T�dg���I���O8<{�>'!�>,�>q���0���ƙ?�q��-Fο�'��#����X?"n�?�F�?�?�<;iw�]�z�����4G?�r?�^Y?��-��]\��'(�6�j?����+n`��y4��3E���U>^ 3?&&�>L�-���|=��>5��>�9>}/��Ŀ�̶�����n�?M��?�a�`��>���?�Z+?�Y��(��ڢ���*��Ty�86A?#42>���a�!��_=�������
?h�0?�'��<�-�_?��a�N�p�1�-���ƽfܡ>�0�h`\�������.Xe�d ���>y���?~\�?��?b���#�2%?��>����BǾyi�<���>�,�>g:N>S0_���u>B
���:��i	>���?�|�?�g?8�������V>��}?$�>b�?�y�=a�>�c�=�򰾣-��o#>[-�=��>���?D�M?J�>NX�=��8��/��XF�xFR��"�I�C�J�><�a?P�L?�Mb>�)���2��!��ͽ�i1�x,�8W@���,�\�߽�-5>'�=>�>��D�Ӿ��8?U�7�:u忠�h�2x����u?l��>��>;��y�Z��熽4�p?j>ˣž�ض�R놿�Pܽ���?��?���>�ſ�=>�=�wi=f��>�!�>�e �O�J��G¾)5�>��D?��c�*���Q��`��= �?�
@X�??d��	?(��V��)P~�Lx�`d6����= �7?�:�Q�z>M��>�T�=�jv������s�̺�>B�?<��?���>��l?ko�H�B�Ê1=pB�>��k?�X?�o�����B>��?��� ���k�bf?��
@�v@�^?/��޿�A��M���������={O��B,>]����=����(}��@�$��#\>X�>g��>u&q>�U->۞�=5��=W߀��q�Sģ�#���9�B�y��	7��Y���C�o�;�ھ_���f�ֶ��?��y0�t���B�<��=��U?� R?ep?�� ?]9y�J�>e����H=*{#���=?�>�;2?�L?̓*?��=m����d��W���H���Շ�&��>�lI>�y�>�9�>��>�p�9��I>�/?>ƀ>�� >��'=�&ߺ�^=��N>�H�>��>�Z�>� $>��>�®���}�r���Z��U%���?��� C�kO����v�貾uN�=��0?�c�=�^��_�ʿ����Q&L?]����!�@E�0�F>�?4?�]?��%>[.���ӽ����=b��Ծ����>�� �����=/�#�O>\�)?Q�7>�r>=�)��v8�t�?w��Y[�>�+?Ñ��J[��=Bt��/'��H򾯀>G��>�ߒ�/4��������N�D���z=��$?��	?��%����ӽ�����>\��=f8M�^�>=[b>�:=zN��,_N��ͻ���=%Ʃ>Ik�>P�=U�=���>��p��Y�R��>e�>=�>��.?��7?���;53�tf]�-�$��M�>_L�>7�M>vڣ=#�V�q= �?��I>0ke�΍��yQ���u{G>I\'�b�ս9������=����Zo�=M��="��LT6�n�=$�~?���K䈿R�9e��mD?�+?�=_�F<��"�E ���G��)�?g�@�l�?��	��V�2�?�@�?�	��õ�=�|�>�֫>Oξ+�L�l�?� ƽ�Ǣ���	�@(#�US�?��?=�/�xʋ�(l�"7>^_%?_�Ӿ���>���&���櫆��u�5�.=���> H?�����V�R�@���
?�?8���[��M�ȿʌv��K�>��?��?�9n�"T��d�?�_�>(z�?�X?��g>��۾ЕY����>ǟ@?�Q?�p�>/��7�(���?��?Lԅ?a�@>���?��]?`>�~�>�M��n�������1	��#_�>V0>$�̆�N�
�/L�� ����j�����c�$?�I�=X��>TR�������=ڈ�=C_���뺽Ra�>��k>yӳ=so>�?ٍ�>��*>5*|���l��Gk�Yv���K?��?���5n��9�<��=b�^��*?R4?ךY���Ͼ�ը>C�\?���?[?k�>����9���忿H���ܖ<u�K>b$�>"Q�>����kWK>!�Ծ2D��i�>җ>�飼�:ھ�(���ॻ�>�>^b!?��>��=x� ?�#?(�j>�'�>�_E�z9��g�E�2��>��>WI?��~?W�?�չ�*Z3�����桿.�[�k9N>.�x?�U?�ʕ> �������EiE��>I�������? tg?�Q彍?�1�?��??��A?�(f>���pؾ몭���>|� ?�-��NA��Y&�����?[�?ʇ�>�Ϙ���нq�鼨q�5����?Z�[?�%?�m�`�GHƾf?�<�����( <�.C�F�>�>>�6��m	�=9A>�Ъ=�l��7���<��=�>}8�=*�:������5?^�ٽG����=�u��y0�ܱz>��=9��>_?r�i����� �������MIP�v��?�!�?���?Eo�1c���?�?�?���>/꾁�ξ�J�}��`|��{~2�H�t>���>�7Q>ɾ��.s���n��l*������>���>U?�w ?!�E>���>�韾��$�������V��N��e1�F+����0�+� �O�(��Ⱦ��~�Mʖ>kL����>�/?D*U>װ}>?q�>��o�G��>�2�>��>M��>r�B>��>p'�=,�Ӽu��KR?����I�'�V�辳���z3B?�qd?F1�>�i�5��������?���?Us�?�<v>h��,+��n?�>�>,��6q
?dT:=9��<�<�U��F���3��g�J��>-D׽� :��M�cnf�Dj
?�/?���<�̾�;׽W���G�=8Ά?�3,?z��/�L��o��=a��|L��I5�F�u�����6�,��^s����V-��S〿o{&��m=� ?��?�a��Η�Yl���8�,�>���>z��>s��>:L> �������_�$~'��t����>(��?t2�>��C?SjR?�
O?�Y2?>�k��>^���?w�Q=i*?B?��0?��3?�EM?�?��7?to>}��K������g#?Q??R+C?L�>��?������ ����;IΪ���d�.�=�s�=͗�� ��;f�ؼ�=�U?ۢ�D�8�����mk>Q{7?y�>#��>����(����<��>Q�
?�H�>�  ��xr��]�UK�>���?�0�K_='�)>��={H��_�Һ�&�=W��"��=�,��ϫ:��!<���=���=׵t���s�M��:�\�;y�<�t�>��?�>ED�>m?��թ �����^�=6Y>�S>�>fEپ�}��$����g�^y>�w�?Kz�?h�f=	�=Z��=f|���T�����1���!��<��?�J#?�VT?Ζ�?��=?�j#?��>=+�yM��q^�������?t!,?��>�����ʾ��Ӊ3�ܝ?i[?�<a����;)�ڐ¾�Խɱ>�[/�f/~����<D�R������R��4��?쿝?NA�T�6��x�ڿ���[��y�C?�!�>Y�>��>S�)�{�g�q%��1;>��>jR?S#�>��O?<{?��[?ziT>�8��0��Cә�rK3���!>�@?���?��?Yy?�s�>t�>�)���XT��/��;�ނ�GW=�Z>���>�&�>3�>���=<�ǽnP����>��b�=��b>��>n��><�>��w>�B�<��I?M��>쾾�c�����d�� x�^|?��?�8?�;g��Q�It$�,fپ�	�>O��?[�?��)?a�c���=pk:�h���.���P�>��>n�>�ɩ=$Q=��=B��>���>�F�����76A��@O�V�?l�S?U��=�Vÿ)l��!x�*��P�˼�E���`L�V����r�A�o=�ڈ��
�j�����G��<��׏��.��+ɒ��k��z�?��=��=[�=��;�Q����<�M=�^���×=C�ּ�~�<�='�ց/�;c���)�PO<	L�=Ʋ�rž~�s?E?��*?�B?�l>�{>K$\��3�>�l����?��^>B��������i:�h��s���Hzؾ�ؾ�-h�ض��<>ɊK��|
>��0>�Z�=��<��=uY�=Q��==Z�x(=��=#D�=�и=I)�=�h>�A>�uw?������N��D����9?x�>`H�=��˾BA?��D>=i��Vo��*���~?ң�?�P�?�
?�d����>㠾h�Z��=\<��P>e�=�8�ퟸ>�<I>���������Ž���?�I@�=?���'�ο��(>�f,<���=[�E��[S����j���,=�/?��V�\�G��6�>$�.>����N׾Xc>v\>̈́�����|��ok>�D:��`=$">跪=JI>>P->�����=�U>f�B�U�O>�f0��W`��-��q=ި�=u�k=H�C�)��>b�?%a0?zXd?�5�> n�>ϾQ>��I�>��=OH�>�=qB>[��>��7?�D?;�K?p��>���=��>��>b�,��m��n往ʧ�>��<f��?�Ά?�Ӹ>��Q<@�A�?��f>�`(ŽFw?�S1?ck?{�>S���ۿ-m��'��(���	�c�<n��3+ ��p#�p����^��>���>�@�>�ҩ>)T�>��(>jy>�v�>�4>���<S����Q<�y�=�<�Q_������<
:=�j�<�#�	x����=�މ;h�=z�=7�T��@><v�>�>?F�>v��=�4���)6>�8��Z&H���=�f��z�A���j�m��\"����>Gl>�m>���mv��m��>	�H>Î?>�l�?��f?�
>����#��E%�����m�B<Uy1>A�>/��9�N� \�z�Y�/Ծ0��>�1�>� �>�{l>T�+���>�w�r=�1�V35����>�ٌ�9���	�3q��I��'���R&i��fC�s�D?T1��� �=�~?�I?�ӏ?��>�;���׾�0>E���=����Zp�T씽�?Q'?���>�X��D��H̾G���޷>vAI�F�O���-�0�ܡ�_ͷ�ꏱ>������оE$3��g������ݍB��Lr�\��>��O?��?�9b��W��5UO����:'���q?�|g?��>K?�@?�%���y��r��,v�=��n?���?K=�?<>)7�=;E��s��>)	?܌�?%Q�?��r?�[@����>�k;ͥ">�Ǖ�3�=ES>h]�=x��=�w?�
?};
?��� �	��{�\�6�\��]�<��=�>]�>�r>}�=��n=V�=a�[>jp�>���>]�d>鴢>���>������%���,?I�">��s>�"?֦%>$�;0�ѽ���<�i>��Z���y��W���"��^=�=m	>��==P.�ܞ�> 2��Ë�?-�7>-��0�)?���-D�<UZx>� �=A�F�@�>��>E�>X9�>;�>q�=4��><�9>����>9<�U}��M���"�mw�9��>]�j��]�w��C��B���O�������AX�X9��O>�ى�;m��?!bo�3U���#�Z�2=�8?���> �3?>j���_��o=b��>ѧ�>	���Ȑ��	��̸���m�?���?�;c>��>K�W?�?̒1�$3�vZ�(�u�j(A�*e�K�`��፿�����
����(�_?�x?,yA?�R�<":z>P��?��%�Vӏ��)�>�/�%';��?<=q+�>*��6�`�|�Ӿ��þ�7��HF>��o?5%�?rY?5TV�V�Q��_>�8B?;?�[x?44!?c8?�d�P�)?�/>�?}?�3?<�2?ՙ?οI>P�!>�ʻ�l�<e����;��W���e����%�<��=�	�<���ڏ�<c�&=?��<�<q��	���6<k�< =T3=�yx=f�=��>��]?���>oE�>��7?\*�fB8��f��q�/?�xA=����bl��]���
���>��j?e��?YfZ?�c>�_B�A�B��>ĳ�>��'>4\>���>��F���=ښ>��>�<�=ZaK�m򁾫�	�V���J^�<>�>���>R�{>)��#�'>�F���z�K�d>�HR��ͺ�U�S��G��1�*�v�)I�>��K?��?l7�=9��f��QGf�v)?�C<?�5M?X�?�*�=��۾I�9���J�~n�P��>rI�<=�������~�:�2d�:��r>a>��C��ü`>߻�L�}���p�<�  =�{�#>�h$��N^=���~¾�����=�,>�ߏ�j��e������/�S?�>��Ͼ��h�����R��=�c�>�Ϲ>#�[;��=�DJ�ϩT�@q=��>.T>\D��-����F�����:�>\�9?��_?Q��?���<5;��E%X��W��T`"�%T���F ?�;�>���>3�=� =�/ξ�p�b_u�"�T�� �>�`�>�:2��pQ����L��/q!��,g<�?cX�>f� ?V�?3>�>�0h?a>1?G?ˤ>^4���ʍ��!4?��?�=>%��e���(��ca�jL�>�$V?��>ˊ>f�F?\�8?Pa3?3�7?h?":!>@��ؔF�|�>}ފ>�5��ÿ;.>&�j?6F�>�R?4�?a?p���ǟ��9�=<�6>dg���BN?��E?�3?��>���>�ڡ��\�=���>��b?�7�?	�o?e��=��?N&2>���>��=>y�>~?<KO?��s?��J?��>�O�<A��n��gs���P���w;8J<�x=8����s�ߟ����<�_�;����>�� 1�vE�T?���t�;�_�>��s>�
��.�0>@�ľ�O����@>���-P��eڊ���:�޷=��>��?��>�X#� ��=,��>^I�>S���6(?��?�?�!;�b�8�ھ�K���>5	B?���=��l�������u���g=��m?��^?e�W��&��H�b?��]?�g�=��þ��b�_���O?f�
?��G���>��~?V�q?O��>,�e��9n���Db���j�pҶ=zr�>TX���d��>�>��7?�N�>1�b>�&�=t۾��w�q���?��?��?���?�+*>�n�$4�7ѾG𕿍zV?���>����؅<?L�'�=��R���/����z�Lˮ�n@��hx����o��p3�s�L�G��=��?ǂ?�x?��G?��ؾ ��R�E��ϊ��lV�;微�1�#-���B��jH��h��v������q[%=�Hz���D��;�?oc&?W�1���>ŗ�^�뾴;Ð=>:ؓ��[����=����EU=��V=��_��F&�ͣ��M0?�>���>�?;?g�Y���>�8�.���9������3>��>�I�> e�>H���[+�V���?R̾���R�н(H>c:P?�W?�z�?�a�=�X6��&������y=� ��n�.�L�g��>�Iؾ�����_=���K���w�"���>��Y���&>ڶP?8C�>�5ͼ��s?�VZ?��Ǿ�k����|>���_=d�>q�\?�a�>���>sޱ�BtB�c��>r�l?���>!��>� ��,���{�s`��� �>=��>j��>�Nm>5�*�jW]�� ��
R���;����=mPh?�W���f����>��T?�Q�:�<@�>n�<��y�{���y:��>ܡ?���=j�?>�������6ty������2?)� ?lq3���Q���:>"%?=ف>NI�>d4�?�0?�������=j.?��Z?��?d�M?��?��=-��m�ܽ�v2�F�I=��>&7=>���=�(>���$~���}�e"=Tub=�?= ���j=���_jf<i��=�;O>�'ٿRzS��޾���n������;� ������Դ���Q'��𕫾����v�~�=6�(�����3��򐌾t]�?���?Eξls��!���V��:Ƚ��?����l�������L4��V��lu�%)��,����S���x�Y���)?����#ӿ����. ��?�H?}�?Yw�x�?���8��ˡ>0b�����=qJ�����9���$y��yjk?�&?o� �gu+�f�>*��>�j�>�.#>�Y��O������k?J�$?3�?Tv�?�ſx˫��VH=7��?w�@�|A?1�(��쾢V=��>��	?��?>�P1�H�x���V�>�;�?���?~M=�W���	��e?7�<�F���ݻd�=�G�=gS=��
�J>�V�>K��CZA��AܽV�4>�م>Wz"���!^��_�<��]>��սp7�����?�
T��^���)�������->`�L?���>��W=-+?�F>�U�ӿ! o��T?u%�?_��?��7?1^��PC�>6d�f�L?;uB?�b�>C����|��~�=^�;�Ҿ�<�'ؾ7?c�=�=���>g�M>V�:�/���|��(������=�;Zȿ�����j�#=PWϼpi������½v�P�U,���b�c潽�D>_>p�C>5�}>Y�U>��e>[�Z?��l?з�>�m�=����t������;Ê����!�53l�g@��ͷ������Ծ��f�"����i�Ծc�>�Sq=.�P�P���ğ(���\��6���/?%�=ʒȾ5�F��!����ʾ	ݤ�ո���m���־#M3�%�r�tנ?N,H?Uv���'\����#v�w��G�Z?}g��������v! >�`�K�;�O�>&��=��ؾ�:�(�Y���1?�P#?Pҟ��?��z�>�3�����;z%?��?WK�=6��>�V,?W�;�-����`>=gD>���>�X�>Л >�������� ?�e?��ým��<��>΋;魶�!�˼�K>����0�f9G>׋�=�
��Y����{��}=�(W?���>��)�6	��a������#==z�x?��?�7�>2wk?��B?m��<q`��\�S�*�+�w=��W?�%i?��>/���}оw���5?��e?s�N>Ejh� ��_�.�R�$?��n?�[?F"w}��������n6?v|?��T�����G�Q0%�w}�>��>{7�>ROA�FF�>}@?v��T��Ɔſ��'�۪�?@U� @�Q�=�#�_��=2^?|��>�Q��,�̾iH+�ԁ���S�<I��> f� ���R�Z�+�3�V?���? ?����4�_��=&��1��?g�~?b�� ;5=��=n�%'��B'�/��=�����Խ
���3�a��U�����]!�<Vi>��@vC��V��>��۽� �(
ɿ&����ƾ�6o�v�>è�>?-e������:��{�u��SW���V���E�E�>��>�Ҕ�2��K�{��o;������>�h���>e�S�	$�������5<	�>2��>���>�[��8���ř?!U���>ο|���֝���X?�g�?�m�?�o?�7:<�v��~{���_+G?��s?mZ?�;%��H]�W�7�h�j?P`���V`�6�4�JGE�U>�"3?OB�>i�-�߰|=h>���>g>�$/��Ŀ�ض�������?Ɖ�?�n���>K��?s+?�h�l7���^����*�qM.��<A?e2>���ں!��1=��ϒ���
?_�0?Fu��/�U�_?�a�T�p���-���ƽ�ۡ>��0��e\�yM������Xe����@y����?K^�?a�?յ�� #�T6%? �>_����8Ǿ��<���>�(�>�)N>SH_�Բu>����:�i	>���?�~�?Kj?��������V>�}?�$�>��?�r�=�a�>�d�=�𰾁�,��j#>�$�==�>�g�?��M?M�>MY�=��8� /��ZF�GR��#�(�C�G�>��a?v�L?]Lb>����2��!��wͽVd1��C鼡X@���,��߽�(5>^�=>G>�D�{ӾGM.?C>&�M5ܿ�5�����o�S?L��>�8�>�y��y���c�'io?&�>!��1������:彽+�? ��?W� ?������b=`">�>��>m��6�*�u���>��F?H�;�yʄ��搿�K>d�?��	@���?�i�K�?8��𠊿��w�9��25�ro�=��4?Iw���Ju>�h�>��=�q�4^��{r�)"�>-ذ?���?�B�>�:g?��f��7��N=.�>5�d?���>�P�;3D��A�L>��?:y����������h?��@d�@�c]?�'����ſt���}����&�V��=iD�=��>�6�� �W=ŉŻW�ڽ���s��=���>�k�>��v>�>J#$>C�E>��z�_a��ʖ�mk����Q��r��e�9�B�J��Y�{�i.�ʾS��E�H=V���d^����ebZ��_����=��U?R?Wp?j� ?F�x���>h���E=f�#�i΄=m.�>�h2?#�L?��*?@Փ=;�����d�^`��4A���ȇ����>�sI>��>zG�>�%�>�nV9z�I>�/?>��>�>.Q'=8J�Ad=��N>SM�>���>�{�>B�>��_>2Y�����&`��$ ��~�>���?�����?���!�-/ɾ��K>[$A?|��=�qx��Aȿ�����A?��b�dg:���$��/T>~?�� ?:F$>:h��V/��P�=!���=�,���>�v��⦾����q�>@�6?�)]>>(�>�:���<��Z��@���&�>ng<?1��+a
��{�f<�,����p>���>��K���Kt���*��-�E��c�=L�"?U?AR�r����9}��������>!C>�'�<6��=׾K>�[������[���=�� >� �>L?�*>�?�=[ã>�f��}�N��X�>�B>Q�+>��??�O%?x��u���u����-�5�v>Ka�>�'�>m;>�J�_�=���>R�a>Q��]儽oj�{�@�D�V>�}��&`�g*u���x=ָ��4��=�	�=C ���<���%=�~?���*䈿��e���lD?W+?w �=��F<��"�D ���H��E�?q�@m�?��	��V�@�?�@�?��/��=}�>׫>�ξ�L��?�Ž:Ǣ�Ô	�$)#�hS�?��?��/�Zʋ�9l��6>_%?�ӾI��>,��`7��a���u�^&F=N1�>�H?�����
p���@�C�?��?��ǣ�$ɿ�&v�9#�>�a�?@��?n�5	��^_>�R�>�p�?,�V?�^>g�ݾY�P�.��>��??C�R?eԱ>��Җ$��K?@�?��?�B(>�G�?�Z?���=�ą>��a���2���������F>�Ry������E�����]��0�o� �\�?Z!>=�O�>�~ѽ��L����=7m<�i��'(^�Ok�>��>����o>eC?懋>j�q>d���bT��g���Y�P�K?���?����8n���<O��=��^�6'?eQ4?��W���Ͼwި>��\?���?��Z?<p�>����:���忿�y��/��<�K>|(�>EE�>_����<K>��ԾFD�rr�>9ȗ>����:ھ�,���]���A�>�h!?&��>�ڮ=֙ ?��#?��j>�(�>1aE��9��]�E����>͢�>�H?�~?��?�Թ��Z3�����桿��[�6;N>��x?V?ʕ>`���񃝿�lE��AI�v���P��?�tg?�R�)?:2�?�??b�A?e)f>���(ؾd�����>��!?���K�A��Q&��A��t?~`?6��>T:��#�ս1*ؼM�������?-\?:&?����1a��þ!��<"�F�d��� <�B��>so>�x���)�=��>�ΰ=�3m��56�]g<��=l�>���=�7������-,?��;�Z����b=�v�eu4��>�>�S>�Xž�fS?����5M���ѱ�d���v���埓?��?HƗ?��I��p��wD?5ns?`
?�8%?�sʾ}���ƾH���{4��ۅ�$��=���>��ٽN��|���C%���I}�����%0�.g�>�5�>��>��? B>(/�>�~I��r/�1��Iު�Dm��j �L���0�����*��d��Ӓ���־�(ꦾ�L�>�����>�h?<j>���>��>�¼����>L��>�`�>o?�>�y>�>8>�]���R��KR?����+�'����Ų��i3B?�qd?Y1�>�i�;��������?���?Ss�?=v>h��,+��n?�>�>=��Oq
?�T:=�8��;�<V�����S3��c�7��>�D׽� :��M�Xnf�mj
?�/?M����̾�;׽�j��߼�=��?�"?'����P���l���b�2P����S�h��皾o�-��Ju��䒿sͅ������p)�̆e=e� ?�c�?ϓ ���������j�QB�`�>@��>0�>��>��:>�0��"$�Yk��%��������>Tg�?��>�0F?��E?͓>?<�4?T�> Ο>��e*?���=(��><L?�6Y?�,?A3?}�	?#�)?�7�>͖���B��߾O,?�iD?�r?��>��?ج�{CL��ɽW��=h�������n%>pk�=��ڽ�$���ȼ�m+>�X?���d�8������k>s�7?s�>y��>F���,����<��>ʵ
?�F�>y �,~r�"c�`V�>���?q����={�)>��=����+�ҺPZ�=����P�=$5��9~;�1k<ׂ�=x��=�0t������:���;m�<�t�>5�?���>�C�>K@��!� �G��pf�=4Y>�S>�>4Fپ�}���$��w�g��]y>�w�?�z�?P�f=,�=n��=}��}U����� �����<��?9J#?�WT?j��?}�=?[j#?��>+�dM���^������?w!,?��>�����ʾ��։3�۝?i[?�<a����;)�ސ¾��Խӱ>�[/�i/~����>D��텻���X��6��?�?HA�V�6��x�ۿ���[��{�C?"�>Y�>��>U�)�~�g�s%��1;>���>lR?�"�>E�O?�={?��[?%mT>��8��0��Hә�"�2���!>@?۱�?<�?�y?u�>$�>�)��ྲR������߂��W=$	Z>$��>�(�>��>U��=g Ƚ�_����>�.^�=�b>���>���>6�>p�w>XV�<f�I?=2�>7����� ޢ�s�p��C��&�s?=��?��<?n-=�u	� �4����u��>���?���?�&?�`�v�=�+��ǯ��u��W�>���>3�>W��=�d�=eH>4��>��>�k	��D���:��=�?qtG?��=!�ſҼq�X�p�����V+c<�����e�*���;[��[�=�x��ϫ�輩��[�w���c���ص�߉����{����>)Æ=eX�=0�=���<�P˼!��<q�I=/M�< �=Gq�m<��8��Ի蝈��%��|X<��I=����˾{�}?8I?�+?=�C? �y>0?>�p3� ��>���VC?
V>��P�Ŏ����;�<���L����ؾ$x׾_�c��Ο�
I>aI���>`>3>�6�=Ly�<Q.�=@s=��=��O�$=�,�=z[�=�b�=H��=��>�O>M�|?�t��5��j;�E�O��zI?*��>K�	>�i߾7?��>�S���$�������?H��?�,�?�(+?n�*���>�����;>���<�U��S��<-A�=4�=���>5<\>�!� 8����p�PJ�?h�@XB?<ل��(ϿG�/>��6>��>s�R��y1�h�[��Mb��&W�]�!?�o;��̾,|�>8P�=J�߾sǾX;,=�>6>�wb=qj��n\��ҙ=���R7=Fm=(Ή>xD>s�=�m�����=��H=�I�=Q>I����1��.%�o�/=+��=�l`>�|%>���>�?�_0?�:d?�)�>%�m��)Ͼ�.��eo�>P��=�@�>-C�=��B>3��>u�7?�D?��K?���>���=
�>��>�,�Q�m��_�����y�<L��?kφ?�۸>�P<|�A�ޙ��a>�F�Ž'v?[1?|q?F�>�|�~�R�����%��ν!(7�w���Z����<��D��qX>[�?�t�>NT�>�#�>nqY>z�s>�ƫ>M�>(�A�ޥ�=:�=jlj��!ܽ#��-b7���=��>��<Cw+=�Z=��t�漃����(���<�h�=��>Xނ=A*�>�2>������c>JNR���R��/<�����e��l��郿u�-���ٽ4X>]s�>A�T��$��D[�>���= �(>���?�`_?|3>NIw�@Z�&	���t�;����6>���������O���a���_�g�q��>�&�>�>�>��l>S�+��?���s='��15����>���D@�����Rq�hC������!i�}�-� �D?T*��� �=�~?�I?�?�.�>�����׾��1>Q����=8���n�.W���?W'?��>�뾥E��H̾D���޷>�@I�,�O���W�0�%��-ͷ�(��>������оj$3��g��������B��Lr�T��>!�O?��?Z:b��W��IUO�����(���q?�|g?+�>�J?�@?�%��z�r���v�=�n?ʳ�?Q=�?w>���=�	���0�>�(	?��?&��?��s?c?�,o�>�;-� >[옽J#�=΢>�r�=�)�=�q?{�
?d�
?�g�� �	������^��+�<פ�=:��>�x�>��r>�%�=m�g=N��=e>\>���>�>��d>��>�K�>䛾k�o��>���=u��>�<K?<�N>�V>#����G߽�4�>;?��t�u�}�@�4F��s�H=_��=@�<.���ˈ�>��ο���?yY>�$%���=?�L���}��>��>]���|�?�a�>T�>���>��}>�>KJ�>�`@>5�ξG�>�<�`k!���D��P���ľl��>�����h,��Q
���ڽ��L�jn��~���i�󒁿ys=�a��<Q��?���m���%���C1
?��>K
4?UΎ��m��h�>��>���>����0��o-�������?<��?�;c>��>J�W?!�?Ȓ1�F3�vZ�(�u�l(A�/e�U�`��፿�����
����'�_?�x?,yA?�R�<+:z>R��?��%�Zӏ��)�>�/�%';��?<=q+�>*���`�|�Ӿ��þ�7��HF>��o?9%�?rY?8TV�F����>t�e?G�Z?t?_�?�+?ol~�-A9?1A�>��?q�!?g�Z?��+?�F?T.�>��F>�lA=A�a=2�D��W��Չ�+ ���"< ݩ=T�>>E��=Jf�<������z=d����-�� �����;�i�<n�Q=.;>3ٵ>��`?E��>s#>��*?��ҽ��=��ڑ��@F?��>���6^`��a���Ѿ�W�=�l?3�?-X?|>>C���H�#>C��>m�>�W>��>ܾ
�#|r���u;_,>չ>1��=R����zH��1����G^=3�1>���>��|>o����&>����[�z��e>rTP�D���TR�VH�3�зz��:�>l�K?Lg?���=��	t����f�!u)?:U;?��L?&��?꼐=vrھ�%9�<�J�U �y�>w�<���gޢ�͡����;��*P��p>퟾B���Td>��	'澾4p��6F��<�4�=[��(M=G��;�ؾ���I��=�>b��"E"�?���𐫿�GK?�~�=����Dd�\t����>oG�>�/�>ـ6�3�'�=cA�������=���>4�D>撠�b4I�#���l�>��7?3�f?��?��M�#�v�\lL��S���P<=��?*�>�?B�=��>�B������MO��U�_�>��>K��`�I�����c¾Q��k�V>�j?<��>�A�>�3>?��3?ޯC?9�? �
?��>�Y��^���%
$?��?��->�2�����_5��FZ��M�>$�X?�,�=J�>�1?��>?�g�>/�5??�s:>�/Ͼ4FT��u�>)
�>�"c��ĿW�=��H?s�>�~?�_?�	�>D�4���о��\%N>I�U=�?�h+?^%?���>���>�Ǭ��=���>�f?E�?��l?;(�=Ś?~	X>���>%��=�D�>�>�>��?�L?1wp?�E?5��>^;�<�2���Bʽ��U�����rH3<֊�<���=ˡ�<dv�y�-�[=�K<HVJ��"N��*ϼ��!���ü���;�e�>t>������0>��ľ�(����@> v��
!���Ċ��e;��^�=��>�%?���>t#���=�z�>�/�>����(?:�?@?�GI;Șb�~�ھ�L��~�>�
B?��=��l��x��&�u�r�i=��m?�d^?=�V�D���1�b?�]?Xg�:=�0�þٴb�%��a�O?��
?�G�n�>��~?��q?��>��e��9n����yCb���j��϶=aq�>�W�t�d��?�>�7?N�>��b>� �=�v۾��w��q��?L�?��?y��?�)*>��n��3� sݾ=G���~V?}O�>NL��+"?J䊽k���Jwc�P.��L߷��*��ڤ�ّ��V}��D���<O�����;�=,�?,i{?�q?i�[?G5㾚w��[`���o�.HL�Po�/n��&E��-���=�Fˀ���%5��S���;��s�DF��ϲ?%�"?�T?�=��>'.���:�X�þP_(>g�������6�=�±��Xy=��w=
N��� �D����?׹>k�>�T<?4Y�]2B�=�2�W�2�×�]7>�Š>?�>m��>�����F����h۾�:��;�սT_�>T�k?��S?Cma?��rCB����*��I<�Ŏ���#>&�=���>�r���z���&�(I�>4���`*��F��eN(�8�>��K?uh[>>ۖ>�D�?5�$?
�ń��F�x��9��i��>�p?y�?��s>�{-=|P����>>�l?��>7�>|����d!�_�{�6�ʽn�>�٭>;��>�o>ٯ,�?'\�$n��~���l!9�1��=��h?:��C�`��߅>�R?d(�:_nG<��>
�v��!���򾖱'��>�r?;��=�;>�yž�"��{��.��\�*?� ? �P�D�.xm>e|?(\�><g�>��R?	�>W��rB>��C?��j?�0 ?	?���>OI= �<����rZ\�"�=	�>kl�>�iZ=�.�=(M��ɦ�������0Ӂ=i�6�{��=1�=�3��.�u�x?���E>\[տe�N�Ѿ�\
�*+�n���P�B��
=����<?����?꾾Օ��]q�cu��Tk&�̝����m����R�?���?bfȾ���������S����
[?���z��<����1��Y�Ⱦ��4��ķ��c�I>������Ӏ?�!s��л�������&�DT?waU?�x?)�#�|
⾏1U��J&>I�:�Y.��©�ݖ�&�ȿ�X���HL?��?�f��þF�?R�>87�=��y>v�徎Ί�	�7���>��Q?��>`IM��ѿ̝��>=K��?m�@�|A?h�(�����U=���>Ȑ	?"�?>WD1��E�����}J�>�;�?���?��M=��W�&�	��}e?��<��F�f޻U�=_A�=oV=����J>wV�>}}�&jA�8nܽ8�4>�څ>u"�����|^�,u�<�w]>$�ս*��PՄ?�z\�Tf���/�SU���Q>H�T?�+�>2�=ױ,?�5H��}Ͽر\��(a?�0�?l��?��(?^׿��ؚ>��ܾj�M?�E6?���>d&���t���=�/��m�����?(V����=��>g�>!�,�y����O�U���m��=�t��OSſ��ѓ��><�f	� �"�EO����Z/�YW���j��=	�g� >�+)>5�r>��>��>�Ѓ>�2[?ֿc?\P�>�M#>��y�Ζ�����w��=3�������D/��P���������ʰ��p	�9����Un�ɭ;�߭x=�MO�����T-�$�M�ޫ-�$�D?��=�վ)gK�}MV��������J�<�{���T�:7�1�{�k��?�lX?󜄿��n��+�:��<�(<��d?�@��Wľh̾
|�=��ֽe��;X!�>�=�9羳�M��l\��/?�� ?�6��=���,3>�fս���<�/?�H�>�̽<�{�>r+(?%û���L�ݏV>t1>�,�>��>�/
>Jծ�(����=?[aT?zб��Ø�9��>:����Pw�3,g<�{�=}�6�݋���_>��%=����yļ� ����<C@V?�բ>e����&�(���`ռ�T�<Uny?�?�j�>��W?�=?J�=@߾�WL�����a�=��U?�>Z?v�>`�s����Wα��9?��c?�݇>��l��o��1�v/�	�?%vd?��)?���x-v�-���W��v<?�~?!$N�������־���ε>��>}��>� F���>��L?�3������DĿ��#��y�?�@��?F�I={��mU	=�"?��>���"��5��l��֕�<e?Fľ����I�e�׽4�g?�i�?-�?��¾���
>����- ?�
u?����踚�pW-���H���߾�����>�}�P����h�-O�G�޾�
�阨�Q�ýh'Z>9�@��9�2{�>x%Ƽ����0���܄�}�0$�� �>��l>��hڻ��~�����bq�F]��Z���:�>��>hߔ�&����{�0b;�����;�>����>Q�S��3��*�����6<6�>ܤ�>���>�z���	���ƙ?+%��(;ο����_��Q�X?3j�?�p�?�d?;4><Ow�>~{��H�a"G?�s?&Z?��%���]�>�8�&�j?�_���U`��4�xHE�U>�"3?�B�>P�-�ʱ|=�>���>g>�#/�{�Ŀ�ٶ�7���]��?��?�o���>m��?ps+?�i�8���[����*�i�+��<A?�2>)���P�!�P0=�IҒ�Լ
?c~0?�z�o.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}? 4�>{��?�K�=���>� �=KѰ�ء8�$0$>��=`�@��Q?�M?̣�>H��=�Q8�k�.��'F��R�H���C�9?�>��a?��L?�b>虹�r�1�y� �1�˽��1���1�?���0�#r߽�6>�>>"�>��C���Ҿ/�-?K��|���p�M����r?���>�3�>Ko꾿4�����=�"p?Ǥ�>��"�ÿ������Z&�?��@�?y�����~�U>{D{> u�>����d��Ld=x�{?�qԾ4���ܖ��~>I �?.�@��?���1�?6�������]�j�HP�)�A��#�=�^/?�����=�9?�=�dv������5|���>0�?��?/?hd?�zi��G4�Pd=Q/�>�@?5��>yz[=J^��)->��?N�3�m����$�w?p�@}K@�2Q?�����ݿ�z�� ���>P����>��=�#�=cս,��=o�=��0�A頽C�">�V�>-��>��>��8>G�C>X1>i���d�J���A>�����O��>^ �����*�2��tL�_���־56۾�#�	��;#������&�3Q����=��R?��T?pp?���>u��v�>cZ�[=0�/�풩=#��>pz.?�E?�&?ʄ=�.��P�c����.�������>I�b>	��>�9�>�.�>C�� $a>�9B>.\�>=!>��u<e ���c=|[O>��>�R�>w3�>j	>^�Z>���������l���&ֽ�a�=���? �վ��$�]	��1���Oh����=(�J?��=�ʓ�
ҿ�U��nI?Z�=��-��NjF�� 
� �?
7j?չ�=�&���I0>��s=Ti8�(l����$�P��[s�%�J->��?�4X>�l�>Ph0�cF���\�𞛾�H�>�#B?�NǾ���WFy��F�fL۾[�7>3�>�B��%�;��M���GeK��:=��2?v�?�轎����@I�^l��4�L>�${>=%��=v�Q> �	���%�_�Bj&=X6">�ҍ>a?qs(>:��=�#�>�b����M�F�>D�D>�G,>7m>?��$?�W����	��I�+�̦w>�6�>�H�>e*>�7I���=%��>��b>@o	�S���r����>�C[X>�{�4^�R:x�Oj�=7w�����=8M�=J���>��Q#=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ<��>0������n��@�����<��*?h1?Ȥ����(A龰�/?�N�>J�þRY����ֿvcz����>��?C��?�K��߫�	���?��?PF/?�)�=z������à�>)�N?l+J?f�?�RF�7�h�>j?��?C��?��g>�;�?�_?�HZ<S�<`Q�~����ם�+J-�����a�>෼0��j�Z��՛� ���ð���ar��Y=�k�='��>�* �؇z�"/���4!����w�T�_�>%-�>�����S�>�4�>���>�f�>���=�N�;�҄��tK?��?�Y��Sm���<m��=C_�X?��2?{7t��pԾ<e�>Y�]?u�?hZ?�:�>$���H���2��Y����l<��P>���>�@�>�:��b�G>^�Ӿ��7��>��>p��$�ھ�Ӏ�o��9�>a ?�B�>�A�=֙ ?��#?��j>�(�>6aE��9��X�E����>���>�H?�~?��?�Թ��Z3�����桿��[�6;N>��x?V?�ʕ>\�����iE��AI�����N��?|tg?�S�(?62�?щ??a�A?�)f>��*ؾ������>��!?+��~�A�#S&�M��#?�J?���>"]����ս7#ؼL��`U��f?x"\?%<&?����&a�F�¾��<	n$��\K��o<�C�ر>Ay>�=��]��=��>7��=�hm��F6�W g<"��=�|�>���=b97��n��T7?Dk����ʾ��=��M�c	3>�(�>���RA?si�󯗿�C��tF���V��菞?�t�?�Ӓ?�z��!r��E?Ms�?���>��&?��Ѿ����|�� �l�z턾�{3�S>�W�>I4�=^
�v���m���g���ܽ�Y��M�>���>u��>Պ?̴	>Ź><�y���(�}�����Ab�;�'��8;��]0�f��m������]*�	=̾]Y�����>
Wʽ���>Pe?�:B>#�T>+�>v����>��k>��{>�@�>��u>��.>:M>F��;�Y׽�IR?������'����6����0B?�dd?D�>�Vi������?���?s�?p9v>�ph�w#+�d?6�>O���b
?�;=WN��ʉ<�Q������Ն�������>Op׽'":�x
M�8Wf�:j
?I+?E����̾�8׽Ɔ�����=8#�?l{!?� �OZ�v�?rR��U�mpN��4\�s����� ���w�2b��mr��*���@�,�U�>;�� ?X��?��������}���1i�K,���!>�Ӭ>d
�>�
�> �9>�����,���T��-�6휾`u�>�Os?�Г>�x;?%�D?�>?�iU?R']>�r>��� �?��=� C>�>�/F?2�B?�h6?��?�?Ѓj>�)��������þ�8!?^�:?A�'?YY�>���>�=��H��=Ε&=�hF>?#�Q:�����j�=�ݼOڼ�v>Y
V>�m?�%��7�;5��Dkk>/E7?\��>=��>����S�����<[l�>Ӷ?�>@����hq����5V�>-5�?���.S�<�W,>)G�=Ag����g��=�|��{؊=�岼k�F�f�;�%�=�,�=�� RK:2:��9ޯ<%p�>m�?D��><�>�6��+� ����E��=J�X>^�R>�>XMپT���#����g�c_y>�v�?Ux�?D�f=r��=P��=mv��Y��=��]�����<b�?�L#?&ST?��?��=?�g#?-�><&�BK���[��`����?��+?���>��	f˾���D>3�L�?��?hMa��	^)��¾	Xս�5>��.���}�����9D��@��]������"k�?�ʝ?�eC���6�	�羢͘��/��ҚC?:��>^��>��>�*�O�g�f4�F;>z��>FR?��>�O?�{?=#]?D�S>�k9�zح�懙��TN��?#>�??�ǁ?�5�?�u?���>�>�;-���߾)������������QxG=�U>8-�>���>-v�>�Z�=g߮��^����8���=$Aa>C�>��>���>B�y>�<��G?i��>����(�H6��_���>B��u?ɲ�?B-,?�#=���D�|����>/�?]ʫ?�6*?�)T����=��ռ�Է���s����>sr�>��>6��=x�5=��>!��>�A�>�z����%8���P��?+�E?e!�=	ƿ��q�b�p��Ǘ�e�d<��Ke�yʔ�`[�V`�=8���>��=˩���[�t����~��A絾󝜾��{�_��>�o�=>��={�=6�<>�ɼ�^�<K=q�<�=m�o�z�l<g�8�QBл�Ɉ�I#���Z<<UI=�R���ܴ���r?�*T?�I:?;5?�Q�=�ۇ=�dZ���>�V�"?k�f>)���Aľ�$��$�������K���d�KW��͕><�B<;�%>�>��=����G9>�o�=�ud=�)�=��I;�\�=β>:H�=�>�f>[� >�y?!}�������H���-�~�/?�>��=#�Ͼ�Q8?��O>-ߊ������P���?(��?�Q�?�u?}�]�8��>NZ���d�;]��=������=���=��%�#�>��y>�Y%�#9���S��+X�?� @��9?�g��O�п��>�">��%>�`V�C�1����ۡ�N�(� �%?&�6���"��>�Ϯ;PK��nؾAC�:c)H>�C�=��ݽ�O����<�\Խ<Ƞ=���<�b>��O>8sQ<��$�D>���=N�->��u>��=��%�6�>=8z=�y'>��Z>m�>Q��>�:?��0?ad?��>B\u��Ծ8Bþ���>@�=��>rě=��P>�~�>;�6?��C?�I?�
�>AKO=0(�>�7�>z-��q�h꾫�����<Gω?��?1`�>���;�?M��Q�h#<�[˽5?e�2?��?�>!��(iۿ��侗�GM>��==�1=����e7�T�
�4�����z��t�=m�?��?�i�>���>pLS>N�>^�>�O�=J~<�=��d�R	����&��=�'u��a�y��<�IỜ�8=���!ҽ/��;.;߼ā><���<��>]A�>a|�<G�>$��=��߾g�_>����Y��6�샼��TW�Zju�Q�v�� 7��ҽiI�>A%>��{�aӕ��?�Z>߿�=."�?;U?|o>��@���_��Lc�-�T���=�j�=����N��Fa��wD��t˾���>�>��>θl>�
,�:%?�o�w=��8c5��>C{��@��S+�G;q�+A��j���ii�M׺z�D?�E�����=� ~?ެI?��?p��>�����ؾ�)0>%G��)�=e�e6q�,j����?8'?:��>���D��H̾4���޷>�@I�+�O���Q�0���/ͷ�&��>������оr$3��g�������B��Lr�]��>!�O?��?n:b��W��HUO����7(���q?�|g?<�>�J?�@?�%��z�r��w�=�n?˳�?P=�?r>�)�=�����O�>�[	?�ʖ?��?'is?T�?����>`��;'�!>nݖ��$�=��>\��=܃�=�k?�~
?M�
?�͜���	������1�]��4�<j��=f��>�C�>��r>�d�=lUh=�-�=��\>�۞>̏>��d>a�>�N�>U��e
�U��>�Ra�h:d>t�$?�(>h!�=�����P����=->r����q�Vd;{�>+j�>R|&>�gT����>�̿a��?ua>9��EK?���������>:�">�����>���>)Y.>�п>�"l>G�=qcb>N,>{�о�]>�c�|�!�p�F���P���ž*D�>����K���
���ｍcH�md��Q���,j�@n���<��\�<
7�?����p��w$����#�?*i�>�n0?�������&>.l�>�ǌ>?��������掿>T޾�s�?Q,�?;c>��>�W?�?p�1��3��uZ��u�S(A�3e��`��፿����
�t��!�_?�x?&yA?�Q�<�9z>)��?��%�Hӏ�n)�>�/�9';��=<=�+�>�)����`�0�Ӿ�þ�7�oIF>t�o?9%�?fY?0TV��n�=*׊�w!,?=��?��?9�:?��?Q�پycg?��'?�=?� ;?�R?vNA?���>W�>q՘>�O}=��=]�<��e�H��TV��lF˼*��=�>�K�=��2��+=���=�,�;u�E=�g;>�.~��ۼ��2<m=��=Ѧ>�]?�
�>��>�7?���Y8��1��G)/?z4<=ު���튾d����E�>��j?a�?VRZ?$d>��A��$C�L�>��> �&>al\>�x�>f��F�P�=&�>b�>8�=dwI�������	�<]��j~�<F�>n��>|2|>�����'>�v���4z�s�d>��Q��̺�e�S���G�P�1���v��X�>��K?��?��=RX龛(��yIf�A.)??]<?�LM?w�?���=��۾�9���J�JA���>i��<�������"��g�:��(�:h�s>�0��5��ׅ�>�Q����j���G��W�j(>�Q�ޅ3>�7�􍍾N;#9,<-�'>͖ѾsU���Ho����Q?N�=�kӾ��������=���>��>��=eW��V�<ӓ�l�>�P�>+ >%%����񾷯8��XԾ���>]�<?�%_?U�?�4�����=NN�:ג��ݽf�Ń$?)&J>��>�.N>�l�=����O���v��rq���>6��>����F��̾sp�(�B��zW>�a"?�%�>NC?Vcf?�@?�ki?}C?e5?�k�>月<5���H�+?^s~?Տ�=�K��N��T�a�X�b�]�?�$O?	e= $�>�j?(�>?l�)?��8??�?�q>c ��cY�Y �>S�>�h���ɿ�ʡ=�|b?G(�>�o??e?}��><��d��+{�=5��=�#�=Qo6?��-?g�I?N�>J�>�<��h�=
��>�]c?(b�?�l?�D�=<�?�}8>���>�Ƶ=\7�>���>�?!DO?_�q?��D?��>�3�<M8��R���၆��d�,v޻?��<>ؓ=�<��MS���4���<Qt�<�qܻ�K�����ag�Ps���ϖ<�f�>�t>����>�0>�ľ1?����A>����������-�:�M��=0�>$?`�>"�"�S��=<�>O�>�����'?��?O?3�D;�b���ھ��K��$�>|B?<g�=��l��{���u�йj=��m?]�^?J�W������b?��]?mI�4=���þŴb��l���O?T�
? H��ϳ>>�~?7�q?*��>��e��-n��
���Bb���j����=ZZ�>�J��d��'�>��7?u>�>R�b>>�=\|۾w�w��y��/?5�? �?@��?}%*>��n�N.�w��S ���a?�@�>�S�� \&?vJ���ȾQ���X؂��S޾xݦ��g�� ����2��X#�E�������4�=�)?Eq?>�p?��`? ����jb�]��ƀ�p�Z���F��3�F���D�??���l���ě�����v =B�Z�SR��0�?��#?�:2��?����ҾJ�;�T�>ٗ��8��/'W>�'�f��=�mt=��i�� ������?K׫>���>X�D?�TW�ge5�XY/���<���
����=���>vi>�y�>P~�<��!��ce�5�����b������>_h?�\M?Uk?`s�;W�T�UK��K �wۚ=-���z=0Un=��&>�6����H��h9��T�M���&a6��犾��	Et=��f?��>��"�
7�?�kU?���ӹѾ�zd��QC�f�U���>#��?�?���>C��|'O�p��>e�??Q�>��a>,�I�#�	��P~����`�>G8�>G�?�h>r�n��bS�
ё�&�JN��M<Яn?(�s��3w��a>�J?v��2���TZ>�W;�	��������|�?>8m?��@�&>n&��s:澗[��9�о,.+?-d?(�/��M1��C�=�$�>�?�?�Fk?�>>sb��8+Z>N/A?��b?�=?y�1?i��>/�h={�ʽ����<�t��=��>Ȗ">r��=@8>�CM�H}W���s��ԍ��(8="��9���Xc<>1����Ļ��߽�.>/`ο�F�⾟���d������%q/��׶��Ӿܼs�sK���\��7Ǿ
�����<x�x� ~i���u�C����?ܧ�?�P���ɾ>����g�@�ʾ�u�>S�>��F!�CӾ�:�Iת��x�������/��.���Z��|���:?kl���׿}���W�w=?�V?��?Z	�EXF���[��>�nd=���=����C�� #ѿ�yn��e?�M�>c%	�����K�>�o�>J�>Q׽�:Ҿ�nԾ�� T??;G2?�O�>�:��ԃڿ��������\�?k�
@�{A?��(��쾙�U=���>��	?G@>��0��@��ﰾ�B�>�=�?k�?7$N=(�W���	��xe?��<
�F�K�޻Q��=qd�=m�=���=�J>�_�>{���zA���ܽ�w4>M�>h`"�"��
1^����<�N]>^)ֽ���5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=����ƞſ��&�����s1=]��A�
�����62�o��`����}H�����=��>iQ>��e>�O>��A>-�]?�'n?7�>��=��7�Fȋ����S�=��c���}��k��j��O@���ھbE�D��(�$���7�Y.�=��L���d1�N?Z�Ѧ0�jw*?�1�=[���K��� =���s���A�;e��"ľ}-��y��:�?p�L?a�����[��&�gP"��q��Sd[?���.���v�����=Ρ�;�].���>�p�=�Kվ��2���X���1?�$?�r��������=|o2�.>�aG?6�>
�5=@N�>
5?���=�f7=��X>�<>�ɴ>���>nd�=��'�]�?6&L?�o��2[\��X�>��޾����M�2*λ<�`�N�)��Y>��#>����sp�|z.�u�=��V?r�><&����8�����E�P�d=o�{?�?�8�>�1h?p�A?|5@=��辝9Q������={jX?��c?p�>�ق��\ʾ�f��G�3?�c?�d>h�v�M��#2�M���o?$�l?� ?�x̻&�|�*����i���8?s�{?�B�sS���x龳������>���>�#�>t�W��`�>��'?��y��y���0ɿ��X�u��?Z!@+@��o<�jѽ���=�_!?ܩ�>ar��c�5�%�ā��'�
��� ?|����.��^�(��-��&t1?I�?��+?��ξ\�[>TUþ슮?�؅?�ҙ���=���"\���!����V��=H�ʽ��=�=��_ ���YD�r��b����Q>k@[��$�>ii���E�Ŀ���������Ӿ��	?�H>��þ�f��Qr���b��B8a��b?��X���>W> 	��Y����|�<��%D�3��>����j�>' ^�3������%o<�e�>�K�>�ф>�ҵ�'���ؙ?����|�ο�������FX?ɦ�?1_�?R~?��<ҝz�C�{�����/�G?�r?�kX?��7�ޘ_�Õ3�>�k?m���'�c�A�2��0E��gf>�81?2]�>.���a=/>��>�+>ܵ.��ſ���{���	�?0f�?�~�N-�>	�?��)?;���������v*��l�4�@?�J6>�}ľN"��L@�����/?��4?���0��]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?2-�>��?/��=�B�><.�=�鰾ݻ(�˗#>�&�=�@���?�M?l�>���=�8�D/�|LF��@R�����C���>��a?�zL?�)b>�渽�'2�!��2ͽ�r1����x@�n�,�a}߽<g5>~�=>;>7!E��Ӿ�7?4�J��ր��I���Of?��`>U�>=������Հ��&�|?�"�>��%�¿nd������6�?���?���>��;@�=Q�=�=b>�3�>�f�K�8��Ə���>Tp;?H[�G����瓿dW�=_O�?��@���?��k�KL?ކ �~%��+!t��6	���r��]�=�80?�!���&e>���>�y >�p�>���n��d9�>%��?f��?[�>�_?_��)�)�8=�-�>�x]?Q��>N4�<)��,�;>	�?'4&�^2����� �_?��@�@>}[?k��ؿƨ��\н��$��k�>L�:�jh�=�q�~Qd=�1�<'�ܽ��5�{����)�>aƙ>&T�>��[>��C>��)>R
������������q.��	�:q�u�����^P���!�F�h
�������#;hx�02	�ߤ½"�=|h�=PT?��Q?*o?O�>H}��(>@+��C=�T(�J�=�A�>��2?\�M?�-?��=������d��G��_����F����>�#[>�]�>��>Q�>��	�1%K>2�D>i�>+��=��<��1�7�=�JN>�k�>���>��>U�p>TjR>��������X���W��W�E>r��?Cd�2)��B��
�?��
���:$>z3?���<�
���Nȿ�n��oa\?����`J��A�*;�>�DW?`�\?*��>Y���O�:�>z���6Ž��>D&�(ˊ��:�% R>ra,?<tD>��>��.���I��煿�žO�>�;?�7�nJ,��煿O�1��2��p��=bg�>��ż#4��Y%��p#����<^](?��?����ľA���d���0�>��Z>u�����:>A,>�^2>�c$�fd �OZ;���=)e�>�}?ʢ->�z�=�C�>em���'Q��/�>�5F>��,>��??o�$?�����CЁ��$-�X#w>_��>c��>��>xJ�j��=�0�>�b>�x���	X
�
�A�q:T>*����a�_mg��y=*喽�W�=��=c��{>�p�-=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ��>X��b���j݆���u�j,=���>�H?����G�U�]�>�z�
?�$?���=Ȥ��ɿ��v�\w�>7 �?Nǔ?�m������?���>rx�?\$X?V`f>�H۾��X����>;�@?0�Q?h��>#���%&��?��?ϛ�?1�s>�B�?�r?%�u=�>��������Q����b>��>�d�>�ر;���a0�2�����ҳ������\?*�D=��>�� �ʐ��5�=V=�[����,?��z>�/�=�r�>���>S-�>_��>t,�W����߾�����I?��?�+��fj�G`��R�=�0��?	?/�2?
�A��־G�>ra?���?��_?���>�������������>�R�]V>�l?��>"��T�4>�;ư&���>D�>�h��L�߾id�lD=r\�>�,#?5��>��=� ?[�#?��j>�>j:E��-��D�E�]Z�>��>�??��~?��?�๾<g3�����롿��[�CN>y?�F?L�>F���K����lB��%G��y���~�?_�g?�d��?O%�?�u??�A?��e>�����׾zڭ��>U�!?����MA�DR&�8��5R?�?[,�>�M��6�ٽ��޼������"?�6\?4&?�X�1a���¾��<�1,�W�/�k<�M���>`�>�{��xB�=��>`�=g�n�1�6��o<Qʿ=G��>n`�=�8��Џ�j82?���< ث����=m
��aj2���E=��=>3W��$c?!	y�����<�������¾�s�?���?.v�?��v�o�o�'*?))�?K�?��	?���k��&�UU8�
��؎��>�=Qe�>$�k��������a��ȗ�I\d���X8�>��>���>�	?M�=>��>k:���a>�fR���ξ��U��$��oC��@�k���xu��o���;=�վv��>��d�>I/ ?�=�>!�>D��>�D̽1!�>O�>�Ӗ>�.�>D�>�]l>�.>xg�=�]h�^*R?7ɾ���&�������PiA?9�d?\�>q�f�髅����/� ?���?P�?�Gx>�Rg�"N*�G�?͙�>V)��!�	?E�?=��	�vx<]ȵ�wO����'��g�>��ڽm:���L�;>e�??O?����cξ�Qٽۣ���	>�p�?"�?&T�4O�)�{��PW�q�a�Oe.���4��c��H�'��G����������،��V���>��?E��?#;
������l�)�c��4�_��=�?���>"b�>�W:>��!�/M��h$�#���&+�>���?��>a1?Ǹ@?*�g?��3?�DE>���>�x>�S�?1	L�G��>M �>�2?y�J?��X?ز?�z:?��=?��E�ʭپKf?e	F?�B??kh�>P۸>���9�����=���>ӞU��K�/���H���}^	� �<oG�=[�6>�w?����V7�"�����h>�76?���>��>pc��CC�����<�?�>�V?��>�(�� q��9�b��>7,�?\��c��<d�*>�i�=����8�:���=ZHؼ{�=V���_�J��)<�h�==��=�RH;S~;N+�C^�iɩ<�t�>5�?���>�C�>�@��-� �b���e�=�Y>S>�>�Eپ�}���$��x�g��]y>�w�?�z�?�f=��=��=�|���U�����A���U��<�?AJ#?"XT?_��?~�=?_j#?�>+�eM���^�������?v",?���>����ʾ�+�3���?E[?<a�����;)��¾��Խ��>M^/�V1~�����D�į�����'��� ��?���?�A�C�6�|��x���@Z��ĔC?)#�>NY�>�>��)�W�g�;"�&9;>���>R?�#�>��O?c<{?�[?�hT>'�8��0��Gә�=3���!> @?���?i�?�y?s�>b�>�)�&ྷS��@����d����W=�Z>���>Q'�>��>���=ZȽ�_����>��b�==�b>H��>���>V�>O�w>s�<��H?�"�>�ѵ�E�������$U|����?���?�;?�>�=Y��<�*��ܾ���>��?���?��-?�\��mQ�=�d޼���|���>�>�>M��>>6�=1��:>M�>y+�>/����	��9�s2��U�?�9O?w>ƿ�q��Kq�&����$h<)㒾{�d������[�闤=&u���G��ީ��:[��L���T��aﵾg���A�{���>]3�=*��=�<�=^��<�O˼�z�<�|L=�C�<A�=��p��At<�;�i�㻐���QL7�
�W<�H=���8�˾�}?�:I?*�+?��C?��y>?<>��3�C��>�����A?s#V>o�P������{;��������ؾ�w׾�c��ǟ��H>�wI���>j43>9�=�N�<�=<s=CĎ=m�R��
=��=�X�= m�=���=t�>�^>�6w?W�������4Q��Z罥�:?�8�>g{�=��ƾq@?}�>>�2������{b��-?���?�T�??�??ti��d�>L��~㎽�q�=I����=2>s��=z�2�T��>��J>���K��D����4�?��@��??�ዿТϿ6a/>kp7>$�>��R�T�1�~A_���b�UY�U�!?�;��˾�P�>s��=�W߾9�ƾ|�/=�6>@$a=S��]�\����=7�z�?�;=%�o=D��>�*C>gû=%ޯ�=h�=�jJ="��=;P>�l��5�1��3-���5=��=�Kb>9�&>ޒ�>r�?�a0??Yd?|5�>~n�N Ͼ�:��`M�>��=I�>��=�uB>=��>r�7?��D?��K?Y��>Ҧ�=+
�>	�> �,�j�m��o��ǧ���<G��?5Ά?�ָ>��Q<�A�?���d>��.Ž�w?T1?�l?��>�K	��j׿����w~���c=���u����־T48�!�˽�B\�����;�W�>\E?��>a�>��>�"�>�	�>Sg>�R���=ܣ��3t=�c�=,�=�tF�q�=k�=s#>�|�8@��<�L1� ~������������>�S�>�F6=�>���=KB��?�=|���e��$�=�Q��b�Y�~f�B[����H�4:%��"�>�v^>�ѐ����Me�>9L>�~�=�c�?�Ob? �>kU��1��:|���J����<AB>���>t
�uX��m�$9�{������>��>�>��l>,�7 ?�Ȩw=Z⾐^5���>Sx������0�E9q�W@������^i��Pغ^�D?IE��	��=�~?P�I?���?o��>Z%���ؾe>0>(Q���=��3q�hs��B�?'?.��>=���D��H̾ ���޷>�@I�
�O���K�0���Lͷ��>������оe$3��g������ߍB��Lr�l��> �O?��?�:b��W��IUO����9(���q?�|g?S�>�J?�@?�%���y�r���w�="�n?ĳ�?E=�?l>���=�۴��$�>�(	?bÖ?���?{qs?C�?��b�>�E�;�!>�����<�=α>�b�=O��=d|?p�
?��
?Lo����	�~����IB^�'��<ԡ=���>���>��r>���=�h=���==5\>�>��>�d>`��>�K�>�}�H��mI?�;���>��?�4>Z}�=a7��z<�>�ͽ�<�������P�7>�M>�H>+�=�?�>&�ӿT�?q>_�6�,t,?�S��)>��>���>�Vb�o��>K�>��;>b�?�X�>s��~�o>���=��Ҿ��>1��0r!�yVC�uR�r�оRH{>�U����%�X
	�����MI��	���G�W�i��0���J=���<TM�?�����k�&�)�������?`��>�'6?�+��Ɋ���>���>��>����|��X���J����?���?�;c>��>&�W?�?!�1�X3��uZ��u�q(A�De� �`�|፿��� �
����_?�x?/yA?T�<:z>8��?��%�aӏ��)�>�/�';��A<=�+�>�)����`�G�Ӿ\�þ�7�uIF>��o?;%�?lY?"TV�l��=rzN;��??1�X?�[u?�,??�:?�P{�R�9?�6_>�9?�>?x�?�1?��#?,��>A�>��&���$�������6��&߽��;�nA�����;J�6�a�;:��A�=����%���K�O<��ڼ6δ�c�r<\ӏ����=���=�1�>'�]??��>L%�>-G7?����8����{s/?�E=dс�f(���K�����DE>u�j?@�?�{Z?gxb>�A�t�B��q>�H�>v&>�\>�Ѳ>���G����=�>n>��=�eJ��⁾��	�����׸�<�� >���>0|>@Ɍ�ɂ(>gZ��}9z�#e>Q��_��&T���G���1�S�u����>�L?��?�=�n��Z��N/f���(?*g<?,�M?c�?��=��۾�:��J����Р>�<�	�}���|���:����:��s>��������1e>�ګ�[����8�M�ʾ�EL>*�	���;,�
�?�9���dx�=�d?>4���A&��l�����W�F?�`>}Ϙ�Z��;<��=2�>�`�>�,=����RO�	���BE=��>��@>�+��}־M�����AO�>:�I?�c?��?,r@='��g���ξVh���ٽБ<?��>Z�>�m>8>}|���B��tn�l>f��O�>1�>�6�:4��q��o��u&�:a9>��>�}�>�0�>��M?#l2?K2??]�?��?�i�>�'k�H=��س,?�=�?���=$5�8�"P��d`�M�>�l?���=GU>�#?��>?�s?��@?�6??2>m$���R�R��>��>�zY�Rп��O�^�?t3?�m^?؟�?�@�>F?�������=�X)>��<�!9?�>?z�?u�>���>��u��=B��>�7`?I>�?��n?�{�=�?��=>*��>���=���>��>�|?�iO?�Kq?�H?4\�>ayQ<����餽�1)���P�{7A��<��=9��=Z�ku����<
|�<R����=�Ƚ���4�ѥ���=�;�g�>��s>����1>�ľ/��y�@>�����9��kɊ��:��8�=[��>�?���>:#���=/��>�D�>>���&(?x�?�)?ؒ;��b��ھ��K���>+B?�,�=1�l����6�u��i=��m?��^?ϧW����M�b?��]?7h��=���þ��b����a�O?=�
?:�G���>��~?d�q?M��>�e�,:n�*��Db���j�$Ѷ=Vr�>HX�M�d��?�>k�7?�N�>=�b>[%�=eu۾�w��q��k?��?�?���?+*>��n�Y4�s羏��k8b?v�>����v$?
��:!���O��쥏��Tľ�g���ᴾ�(��mM���J���^��>����=�,?�Qu?�@r?>[?X����_��SP�k���V�қ޾fq��>���<�-zI�µs�+����3���j�= �p��wD����?�L(?p�F�Ԣ�>\��pݾ
	Ǿ��%>�ڐ�o�1��q=Y�ý�J=��= �J�*���O��}H?��>� �>RH;?��W���8���&��:��7����\>��>�|�>�!�>4��9��. ��UҾޖ��l%��sng>.�c?n�a?�km?���=�zA�l����e^8>0!ʾc��=�q�=�5�>W;C�eo�2�4�/�D��1����[���~���>�??��T>��=C�w?Z?q������#�
=����Y�^��>1#x?�} ?�*�>�5��*����>{�l?#��>�Π>���M!���{�+�̽���>�Y�>�>�>�o>҅,��#\��p��4���QU9��o�=ݒh?-m��va�@�>+R?;��:&&@<y�>S�q��)!�\��AG(��>3�?�t�=��;>ž���ۇ{�����"22?�0(?_�?���Q�7��>Fo?���>w,0>ؖ?r�?�x޾ cV>h�[?�h_?Q�>SY?$��>S��<�������.�����=C��>Jq>xI'>�y>���ރ�=tžٗ�<��=aj+=ǰ�=���=�H!�s�彘G>]Vd>@�˿��R�#�ؾ�����������sj���5<X��� �����h&ʾ�\��:�S3�=:jX�9�k�b�>E���W�?a��?Uq��s��� ��:rr��0ھȅ ?�G�Lz��Ֆ�$s�����Dt��gh�� ����X��:b�H�}���'?��^�υɿ���3��_Y?�=N?Di�?.I��4*�n�Z���>���<kp<Z�羄?���
ǿ���5�k?�6 ?�A�"���9�>�͎>���>T�M>�֏�����.�۽Y'$?8�7?:��>#!��ʿ����r`p<
��?��	@�|A?��(�U�쾨wU=<��>s�	?��?>�l1��2�ް��1�>m9�?��?�N=��W�(�	��ue?��<M�F�b�޻��=il�=e�=O���eJ>�R�>y���A�G�ܽ�4>�څ>ˈ"�&h��.^��y�<�`]>�eս	��5Մ?*{\��f���/��T���T>��T? +�>4:�=��,?V7H�c}Ͽ�\��*a?�0�?���?*�(?,ۿ��ؚ>��ܾ��M?eD6?���>�d&��t���=�6����p���&V�u��=Z��>u�>Â,�����O��J��W��=gI��uǿ m�w��:>R<�
�=@H(����fV�<����,2�|�=�3>��C>Hq>��b>��D>��`?��l?@�>"�>s� ���[������1t=�/���F�3�_��Os�dɎ�jE�"B׾8��t(�*��Qq�sA3�^�L=V�L����x:/��H���8�>�H?���=��Ӿ-)>�����ež�د��"=�����k�)�*~����?��Z?���u[�g����Ž�>��l?��-�����ƾ��=S����=�k�>���=Eؾg=��Y�ކ0?�6?�"��⪐���,>S�轏%#=F�)?m�?gp�<P"�>R &?���ͽ\>%�2>�I�>�o�>1!>;뭾Bv��s?B�V?!&���]�>����jS|�wNX=�x>(3�ʀ��Mdb>�<tu��t`�w�����<P(W?X	�>�)�fR�:$��!��;�==�x?�?�1�>�-k?W�B?^Ȱ<i����S���
��?z=c{W??�h?�f>B
����Ͼ䦾
�5?��e?�O>Ħi���꾙/��K���?�n?�K?c���Fv}�/�����a6?��?L2G������LξI�]����>䭸>5��>��<�Y�C>��W?[������dɿ��.�Fp�?P@j� @E��<��`�Do�<�?.K�>��bW��])�<���
ș��?�!��������[��>�Wn?6܊??�ӻ�R�
�p�>��z����?�n�?I[_�����C���_�m������>�;�2Խ�+��#L��i���?ɣ�����2>Ij@�з����>Q��=Irտ�FÿX���n���6p�ҧ�>˝�>������}�z����~�G�U�WZ��K�>s�>㽔� ����{��m;� ���7�>�!���>�S�O+��Ú��P;5<��>��>G��>Q3��(��ę?jT���=ο������ŶX?�h�?;o�?s?3?9<�v���{�����,G?�s?�Z?g%��I]���7�%�j?�_��yU`���4�uHE��U>�"3?�B�>T�-�[�|=�>���>g>�#/�y�Ŀ�ٶ�>���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���J�!�D0=�TҒ�ü
?W~0?{�g.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?g�>��?�G�=e}�>��=9���3��U#>>��=P�?��?4�M?�7�>-E�=��8�v!/��ZF��VR�s)�ĶC�q��>��a?M�L?2;b>���"2�p� ��uͽ�R1�9�|L@�W9.��f߽U�5>�>>k8>��D�ӾU�/?v�����k��f����O?���>�]�>��-��K�=�?0�>������}��%|�ٳ?��?��?C�N
��{�=���>{#�>`����)���DV">��m?���G���ؙ�#�>�o�?��@D�?kv��	?�G������p����j�����=�p2?Db�-�#>"�?�=EDt�����te��Z��>���?�l�?b��>]a?�e��59���=Ⱥ�>��K?���>�p�<����Y�/>��?�8��6��m"���m?}@�>@�L[?u���N-ٿ2@���|�Jl��N�=x�-�=%�K��*Z:م=���=�߀=	�!>��>�h}>�#�>#�>
x\>[�{>y���^�#����r��B�E�V�����百e��Mc��/��ě��N���3}����ԟ0�������<u��=��U?�R?bp?�#?慽�>���5�=�%�Z��=�O�>Ɉ1?�K?�*?��=�\��nge��L������Uo���i�>|�J>���>F��>�,�>ܫ;>G>�Z>>��>N� >�=��@�=B�P>�V�>��>닸>N�;>�s>�E��B��K�i�%�u����q�?K᜾��I�Kn�����&���PJ�=�.?��>�ߑ���Ͽ-��o�G?������)�Ok>�$/?�;X?p�>�����2P�_�>�{�ci�$�>/��8:n�p�(�P�M>��?-�I>HԊ>>'�&�B��턿5v��'��>ݥ_?����Ľ��5�&RѾq�5>���>����� ��ꈿ?D+����=��?-� ?�l���[ǾS)K=������_>�Ⱥ>��o�Z&�>]��>DƦ<]G��g��,��=�ǅ=���>�E?42	>���=h��>Q[���W7��;�>xFZ>a�*>X�4?i�&?�#��v���Ų��w(%�|>;u�>���>�S�=��<���=��>�h>�C��m��Lܽ�V��bQ>�2n��!\��v���W=/��.�=��l=�f�
Z���@=�~?���(䈿��e���lD?S+?] �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��J��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾS��>���KV��R�}�~qw�~�(=�?H�L?Y��߂����{�`?���>,!о[䢿�ɿ�t�1S�>���?�Ò?��i�̝��1�Ӄ�>`��?� 4?��>�ؾ�Ob���>��<?I�I?He�>ý-�}�𽄀?���?K�?aO>�	�?�r?}�;>M��>�-�����5��̄�����I�l>�wK=�Ծ�P@�mM��;j��l'��@���?ζ<�*�>~3��K���~=Vc���!��Ek���� ?6��=E%�;���>\��>�0�>^��>��s=O��g������L?���?�:�h%p��Ӳ<�>�= �_�X�?�7?���:?hϾ�>^F]?�w�?.�Y?ǥ�>������K@��=���`A�<�J>���>4��>��Z���S>��Ծ	7D��A�>���>�����پ��}�>� �A��>>� ?M��>�{�= ?Ŝ#?{�j>�(�>�`E��9��Z�E�
��>1��>�H?��~?��?�Թ��Z3�����桿̒[��:N>��x?�U?�ʕ>S���򃝿bE��BI�c���$��?atg?`T�?;2�?��??��A?�(f>����ؾȩ����>��!?p��A�_Q&��:�r{?�U?���>N1����սbu׼9���}����?[)\?Q<&?O��:+a��þˁ�<��!�.�V����;#�D���>7�>����Ǭ�=�>(��=�%m��>6���g<XS�=�u�>@�=77��C���,3?v#U��۳���>�����J��4o>E~>�b�O?�[t�7����{��yΗ���]}�?Y��?M��?�F�܀t�T.C?�u�?!��>�Z?�l������7)�Iw�$���3�ϕo>:h?k �=�j�ur������9f���䭽�U�k)�>Nq�>��>��?\�U>ē�>(��^1+��������a�L�#�q@�!�4�<���Aq�Mֽ��t�H$˾���K-�>�Wֽ&�>�g?�J�=��>8��>
�ཎy�>Kaf>;}>�B�>FR�>�8/>�/>��=����IR?����۟'�ؐ�_��&HB?�jd?���>� h�s��g��=�?:��?,x�?v^v>q`h��+��t?� �>���6G
?fz;=C���ӧ�<|��Խ�_2���K�ʚ�>�!ֽ	:��M�ٷe���
?�;?����l̾�ֽ<螾��~=���?�J)?�#'�։Q�Ywo�tX�VS�*P!��ce��F���{$��fq�,U��`���Zc���(���3=�)?q��?�L�H�ﾉ�'�j��~?���]>��>��>	O�>�eO>lv	�$�-�E^���(�l+��܋�>�P|?jI�><u=?02?�jN?�@?�ݾ>y��>�ԥ�Z;�>/t=K��>�?�S?��K?U$6?Q�?y5?|��>8������,p�??��???�?���>CB�>����;���A$<�P�=��u�#�ݽ��>��3>-�<��м�4n<S�f>�a?O���j8������wk>d�7?C��>�!�>ł��E���c��<�_�>�?鼏>{����Er�*�_\�>^y�?�I�cp�<�*>_��=����p$�E��=����E�=�쇼eU9��(<߾=�d�=_�^'i��:��;�԰<<f�>ę?�ڊ>Jm�>����Co ���F�=9�X>�/R>ޙ>��پbu���$����g�@�y>�t�?Ys�?�e=�j�=�(�=�џ�f��Q��!ƽ�B��<0X?�*#?��T?
z�?n�=?AA#?c~>z+��?��_���o��C�?�,?C��>~��}�ʾw����3��?zd?�3a�_���H)�ݍ¾jս�>�L/�<(~�����D�>���)��3�����?$��?*�@�I�6�W�N�}T��-�C?���>o�>��>A�)�T�g��&�7;>���>hR?��>N�O?[{?h�[?`�U>T�8�������E��� >�@?{w�?೎?�x?yK�>��>9x*�ǽ�`���l����ʂ�][=��Y>�}�>+��>�%�>���=��ǽ/��)}>�/�=Vb>�V�>��>���>]�w>�v�<h�H?�d�>����2]�ұ��mt�j��v?\��? ;?���<����5���h�>��?�o�?�"?k`���=s	żE�������Q�>��>F�>�on=n�0=	>+>���>P7�>������O�9�M�e���?�IC?|�=�ƿ�Gr�,ao�	ǘ��W<:��K�e�H㘽��]���=򉘾R����� Y��՝�q���$~��b���	�z�k��>t��=;�=bF�=F5�<������<p�L=��<�&=om��rY<k�8���лHȃ�A�:�h�><�VL=��
�O�ʾMt}?��I?f,?E	D?�[t>[�>.�/�X��>)~����?�U>�V��e����9��ܨ�瞕���پ�jؾ��b��K����>ۃD�?K>?�/>h��=���<��= {r=O��=+�ѺU�=N��=$�=2�=��=�>�>{0y?HU~�f���H���l2?��>S��=�.оP8?ZCY>���h꽿j���{?�}�?�7�?@I?%�_��n�>tᠾ��z:N]�=K��_��=*��=�3����>JXv>.�"�|Y���Q�O��?�]@j�:?ډ�

пM0>3K7>Ż>��R�	[1�*�Y��a��kY�G�!?�R;���;�:�>�)�=��߾LǾFj)=�%7>z�g=V���%\�$��=]v����B=aj=5?�>�.D>o��=����=Q&D=�;�=c�O>�(��/�2���#��z4=Y��=�7d>��$>��>L�?a0?DYd?8�>�n��Ͼ�<���M�>C"�=�F�>���=�B>���>!�7?ݳD?V�K?���>n��=)�>_�>3�,�`�m�(n�j̧�Ŗ�<֖�?�͆?Vָ>�R<ʍA�:��Bc>�.Ž�x?�R1?�h?*�> J�Tѿ_f���q3������p����B��7���A��='|0��'��:��<�e�>�(?��>�e>�="�>h�>��=��I�'��W��	�>C��<.>U�X�9�>�i��G����膽c��$�=e�n�2��Vw��05����=52�>�>�= �>]->۸�<Y>|Un��V�(��<�˾�_N��h��X��!�>����# m>�IK>+;��36��ݼ?2�b>�9�=���?m~?�o->��^��ɬ�hfս#���=B>�
�=�5a��f?��]�m�:�Q�ؾ9��>\��>��>�l>�,�1#?���w=T��a5�#�>G}�����h(��9q�!@������i��Ժ��D?\F��]��=8"~?,�I?)�?Ҍ�>�����ؾ?0>�H��"�=��'q��d����?''?���>����D��H̾N���޷>�@I�2�O���V�0���0ͷ�4��>������оm$3��g��������B��Lr�\��>&�O?��?`:b��W��KUO����^(���q?�|g?/�>�J?�@?
&��z�r���v�=�n?̳�?T=�?w>��=���E��>{M?�a�?Y�?�s?}�@��_�>�`�;3�>�x��)��=�u>Ǽ�=��=�	?��
?�
?����$
�$F����<�^��z�<��=[v�>�>�rp>�T�=��j=Q+�=I�`>)ݡ>⢐>_Qc>=u�>E.�>BG��Y��
?�>�B�>M?���=,;l>�x ��E�����=Ȇ���N���Cg���۽"�=/97>�:�>9����>�˿���?�ۚ>j�>�߰?N��|�=8�>�߀>�(R:���>O��>Ѳ>b�>�9x>��>�>���=�B��?(>�t������W��D�����>)���f���RJ�i�\���+���(]澈?j��%|��u>�nd�<Cy�?�,�����������8����>���>
C)?����"�o�)>�?�#�>;�����0��Ԑ۾��?U��?~9c>��>|�W?D�?�1�h3��sZ�˫u��(A�Q
e�'�`�_፿)�����
�H����_?��x?tyA?�/�<57z>�?��%��я��$�>#/�8);��Q<=:,�>*����`���ӾܶþY1�_PF>Ŕo?�$�?8Z?jUV��7>�7,>��5?4�?�W?�
?iS=?����%?!�>�I+?1\8?�M]?�[j?},?_1�>py<>v=�[�=@LؽlOf�[���S��H�=��[��J�<�5��2,�=
�<}��= ڢ<ޝ�nHN�#k�6A�<�L/=���%,�=.2�>(�]?O��>q��>��7?����8�[%����/?��H=�����B�� �� ���>I�j?�۫?o�Y?F3c>Z�A��`C�kM>I��>�8'>5b^>��>N�󽄍H��׃=ݲ>��>�9�=�I�������	�����=K�<Ͳ>���>)|>2Ս�n�'>����*z���d>>�Q�?ƺ���S��G���1���v�$C�>�K?��?_��=S龅H��Bf�0)?L^<?SMM?��?���=��۾6�9���J�i��>���<`������#��Q�:��>�:�s>1$������_>�3�&M��p���H�����Jj=d�I�9=�d���Ҿ-��%�=��>x#��0� �}▿u���r�J?k��=�f���Z�F����>���>�%�>�b/��ꀽE�@������=;,�>�Z@>������^iG�հ���{>iV?�i?Yl�?�P��'\���T��$1���þ��=�8?��>2�&?��>ld5>�Ǡ�D������<u��C�>� ?�	��=Z�8��D���;��Ĕ>�?�>�� ?��8?Ъ?<Kc?/!?��?��H>V9������J:*?���?��>҆��(��
_d��f����>��[?I��<�;>�?�>�;?��L?�
]?j�	?��=�X$��l�4��>�0Z> �`����"5*>7�)?OW�>uE�?倫?��>LO�M[��ܲA��˿=G�+>��?�fD?��O?�H�>��
?�ԾӧN>��>/�>��?Yr�?��>��>��.=��?P�p=�k�>��%?;�+?8O.?�DF?n+?ފ�>INo����zq������&�<����T�=]� <;�;�= yڽy�N=?�#��V���:=1�����n���];��|;5_�>X�s>t
����0>��ľ�N����@>�~���P��Eۊ��:�۷=���>Y�?���>�W#����=���>I�>��#6(?.�?�?�!;g�b���ھ۰K���>D	B?���=A�l�Z�����u���g=/�m?.�^?a�W�X%��I�b?�]?+h��=��þ��b�щ�Z�O?>�
?�G���>��~?h�q?Q��>�e�*:n�(��	Db��j�4Ѷ=Tr�>OX�Q�d��?�>d�7?�N�>X�b>�%�=_u۾$�w��q��s?��?�?���? +*>x�n�V4�_���ld��O�\?�f�>hإ�6s"?0����n̾�P������Ӿ����糾�)��WΪ����y�8)Ľ��=�?�Kp?�Fx?`6[?������c��-c��ρ��S�*����F���=���?�>G��Er�&y�{���p$���UJ=U�w�Q�D��߱?�?��0���>!��w��m]���@R>Q�������)=ҋ�����<o�=ZQ�|���1��:?���>��>��4?�U��<��Y:��}?�	�քF>��>���>���>Wp��R�@\�Ӿ����\Ͻ'�>Q�s?�K?�Vr?�i�{3��;���7��D
>�F�s<CZ>��?F=��py��.�K��,.��%���'�3􋾛���݅=��6?�B>N��>ٍ�?4T�>�ľ�P���˾r�3��z�=�?�ދ?��?P�^>*��[�1�O��>��l??��>��>���W_!���{���ʽ�&�>�>��>��o>r�,��$\�xm������9���=��h?߃����`��҅>�R?�:q�H<gw�>\Fv�^�!�B���(���>��?�Ȫ=l�;>�rž�Ƞ{�J��N�)?�`?f���^Z'�%�g>'} ?�[�>���>�ȃ?�˖>'��x� <?�?U^?R^J?��>?�8�>�(0=�x���xнW'���;=b��>�]>��=u�="a#���i�Z; �[&'=E �=�� �SսǿP<�F���e<u�%=Z�I>��ֿ��J��?�~y"��O�|�߾p��?+i�MGz�ŨO���������bp�0�"��}Ƚ�{��|�-s��ܫY���?+��?m=��@ז�)L����|�b�ھ2�>�>������ʾ,񰽥�����󾱍���W�J�8���`���a��?�ޛ�ͿaI��������>��?��?!�羝��\#_��P�>�w�=�H��uX��޿��^���]?���>1��_��;��>x�?�f�:��=!B��Tf��>�_�>$�J?Z��>A���Zƿ]6¿�V	=��?~�@�zA?��(����rYV=4��>��	?R@>1�0�i?�����r�>':�?Y��?�N=�W��	�Yze?�a<��F��?ڻ�=Mڤ=:x=��/oJ>Bd�>�\�>NA���ܽ��4>'݅>X�"�8���`^��m�<�]>�ս�	��HՄ?X{\��f���/�U��kR>!�T?t)�>%8�=i�,?�7H��}Ͽ��\�o)a?�0�?L��?��(?Zٿ�Qٚ>"�ܾ݊M?&E6?���>�e&���t�E��=L*�~������'V����=#��>��>�~,���W�O�zO�����=�� ���¿p�)���0�ӑE���=�哽c�۽�.Ž��i�����fW�[[��zo=0^m= �>P�>�t>�M2>��j?B�r?��>�L�;�'��6�S�޾�sp2�R���W�z68��b�p&�D�	��վ���I
�b<��Q�9�A�]<v�Q��Ø�9�W��>��s(���;?08>B��C^��8�=�翾]j��_���4�n=F�˾�W6��yj�\��?4�K?5���\�U�;���,&��<c<�jh?N2_�|= �f�;s��=�9����=���>ݞ�=Ę���w5��V�}�/?�&(?�ࣾᎾ�U�=�"� ]�;?-?�	?r��=3A�>x3(?cĽF��$��>Z�*>���>y��>(�&>����s����"?�+Z?����́�'��>�E�������N�F�$><�PȨ;�
>��;?{���2ϼyݎ��X�=�(W?���>-�)���b��� ��W==��x?!�?m.�>�zk?��B?#�<�f����S�j�"hw=��W?�)i?t�>䈁�	о�����5?ӣe?�N>�bh�
��G�.��T��$?��n?@^?~���v}�1�����po6?1��?W-v�켪�����^�$o�=f�?�ա>��:��?��?������(�ȿv,�O%�?��@� �?���==2�nӥ=��?5�>����Đ��a>@� �Ә���?ٷ���,��?�������N?��?[?�iľ���`��=#���ͣ?t�b?�`��Ω4��6���m�!�Xܢ=�v�= 'G=�4&�)�y�f���Ⱦqh	�N_���4����@>%@����=�>�������ѿȤ��sI㾪��{��>p��>�w�v � J��;r����d�:a��m���K�>~�>��������"�{��p;��#���>a����>h�S�O#��f���Ο5<��>հ�>��>�;���꽾ř?w^���?ο����t��ǸX?mg�?So�?sq?�M9<+�v���{�?��	/G?��s?�Z?:�%��=]�z�7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?��>*6�?���=��>q�=m����{��*>�'�=�:-���?��M?d��>\v�=�M-�uf-���B�4P�N�P<C��w�>��c?T�O?�h>$淽�O%��� ��\ݽn59�R���@��Q%���ؽ��2>I<>�Z>�HE���Ҿ̾'?�6�������#�w>\��>n�U>8j�>H����߽j�����x?��0>e�+��s�����������?�&@E�?�7��~L��v��>���>���=�lݽ]8>�~v�a@B>�<?�@��֩���>���H�>R!�?�@��?�9P���?���d&��!�q�^碾� ���@	>q-.?Y7�,�>h��>9�{= �{�<֬��pm����>C�?z��?�?�,i?��e�W�&��>�Jh>�[?y&$?�8��m��2�>5H?P�0�Њ��L�)�X?��@�@D?O?�P���Pѿ�Ж��_������U��=��=s >Ɠ��ͣ=���<pR�Z��H]	>�q�>c�q>�ps>�9.>�Z:>�h&>_���~�!�8���4��h;�a�V:�#���c5
���\�������u츾��ٽ�F���q� �T�S�����7�=�CY?S�W?�yu?���>i�^��==�x
�k3L=d���<�!G>��)?Y:I?k}%?�}�<(C��pAz�Ql���އ��u����>9�&>��>}e�>�Α>tϔ��~*<�=�>䶴>Cf">�}�<~�D=��=c�[>1ܗ>kκ>=Ď>.�>X�>�X��B���`|�F^�A��׮?�!\��(c�6Ú� �b�$'��=��=@�?A>�E��aȿ<���P?g&}��1��������>y�?`�F?=�d>$���������=�K�e����v>'��O˾=`G�fД>Ђ?r�f>u>ʛ3�/e8��P�2|���i|>�36?�鶾SE9�|�u�̲H��cݾ{GM>wľ>�D��k�Q�����0vi�E�{=nx:?��?b8���ⰾ6�u��B���QR>s;\>�R= j�=5XM>*cc�'�ƽH�rh.=���=X�^><?w*>$[�=M,�>ݔ����M���>�4D>!|->��??�9%?8 	�����ꢂ�~�,�^�w>���>X�>k�>�wI��j�=_��>9�a>��@ჽ�����A���T>��}���^�OYm���z=蜽P��=ٮ�=W{��_=�R+=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿki�>_���[��w����u���#=���>�9H?R���O��>�{
?7?b^򾳩��r�ȿM�v�!��>�?���?Y�m��A��
@�p��>	��?bY?�Ti>�_۾�LZ����>�@?6R?H
�>�:��'�]�?��?#��?��=zu�?�Nm?]��>-A{<�gN�?�¿�����i�B騻\R�>�ax>-:��;h����y���>��$s8�Ȕ�>�8�O{�>����4��<ցR��搾?Z2���>��o>\�C>߭r>�?�{�>���>G�&�R�= ���L���M?�v�?�Q ��f���Q�s�W�����p?��P?ƞ�=��ھ�8�>v�Y?��?�]^?��>��ց�������������s�%>�3�>�	�>819=���>�ľ�O��xl>�>�h�<tmھ�������О�><#$?�v	?�lg>ՙ ?��#?��j>�(�><aE��9��d�E����>Ԣ�>�H?�~?��?�Թ��Z3�����桿��[�D;N>��x?V?lʕ>_���胝��kE�-BI�@���[��?�tg?qS�?82�?��??_�A?�)f>ԇ�ؾ������>*�!?��C:A�)�%��F���?��?2��>=\���ڽ�\ļxa�b����"?�\?�.&?� ��`�����\?�<v$���U��<�=��F>ӣ>�h�����=
.>�߫=��n�
�7��{`<
"�=�w�>u��=n�5�����?<;?Ͽ��eα��(�e��� `��l�>�2�=��'��?����y��ʼ��n����;2֣?��?<��?�<�����t?1#�?S�2?���>�P��E9���t���Ѿ��� �۾L�>U�>4�M>�㾲������y�z���.�R�S�Pq�>�*>�P?�?R�s>ɦ>\��W_n���3�B땾�x�l�� =���&����M�\��~T꽐�Ѿ�1��		�>X,��$F@>�[�>�V[>�>�?�ɔ=Q�.>�X)>+Mw>���>��w=	'*>^�3>�*�=���$KR?-���o�'�Z�辞����6B?:vd?IF�>��h�S������$�?6��?�q�?Fv>,sh��!+��i?a9�><��Il
?A :=o��͈<P����EA���
����>�n׽t:��M�Eff��j
?�.?���d~̾(׽ɠ�����=~τ?d&?.i%���S��\t�jKY��P�9�*�ee�z�����%��s��Ɠ�pj��U���ݑ(��>6=U�%?�o�?���!\��/����m�3?�	�U>��>^��>Cc�>��F>
�b}0���`��+��Q����>�W|?�*�>ЂW?��L?D�L?@� ?�O�=��M>�@����>�c�<��>��?Q�H?�#?��@?��>�~+?MY>�j��*����Ӿ�}+?��I?`�?7�?��	?� �W�g��gG�:>��h���в>\E<�?6�a���� �=���=�d?f��t8�(���S'j>��7?��>�E�>�ȏ������/�<��>ү
?���>6v���'r��+��3�>���?���C,=]�)>��=����Bk���d�=��ȼH��=����?���<��=���=�`V��1����:�ʓ;a��<t�>�?ǒ�>�C�>�?��ة ���`e�=�Y>�S>Y>�Fپ�}���$��i�g�	^y>�w�?�z�?F�f=��=q��=b{��rU�����������<�?�J#?XT?畒?g�=?�i#?U�>6+�"M��p^������?w!,?��>�����ʾ��։3�ڝ?i[?�<a����;)�ސ¾��Խұ>�[/�h/~����=D��텻���W��6��?�?IA�W�6��x�ۿ���[��{�C?"�>Y�>��>U�)�~�g�s%��1;>���>lR?j�>��O?;{?�[?7UT>љ8��0���Й�1���!>J@?j��?��?>y?�R�>q>��)�;�e�����<I�@ڂ�Q�W=C�Y>@��>�>ݩ>C��=��ǽ����~�>��?�=o�b>���>���>=�>H_w>N��<�ZH?�i�>�E��l��(F��o���΂���)u?�V�?��.?4Q�<���=����>�>K�?���?R�'?��^��a�=M���1���wb��
�>�s�>�%�>���=��<��>4_�>~�>]�����SQ5���^��j?5�J?~N>X>ƿbr���{�:>���1X�w���׊d��9����Y���`=�ݙ�F���觾�][��,��df��b���rѝ�^�t�P{?���=��=C��=:�;Gռ�<N�r=Nd�<l'=������<�8��ɼ�ޣ�+q%;g�j<A�5=��v˾�y}?��H?��+?V�C?��y>��>\ 8��|�>W\��Y8?��T>P>Q�P���;�{�����-�ؾؾ�d�������>1NI�1>�j3>gt�=���<�=ut=L~�=
pW�գ=���=Q�=.��=.�=Pv>�->C�|?P���j>��-�S�(��hU&?G��>�Η<7ɾ�
R?;!�=R2��ݺ�\��-�x?���?�p�?2�?�FE�rN�>q����e=n�S=�P�xI!>�*�=_j'�Y۴>��V>/H"�����n�����?0Q@��:?8����ɿ��6>�7>Lv>��R�.L1�fY[��b��Z��[!?q�;�$�̾3��>�P�=�C߾��ƾ1�,=g�6>G�c=�'��C\��Ϙ=��|���>=ϡk=�h�>�^C>+��=Vo��7��=?OK=���=+�O>񫑻=�7�
�.��	4=�{�=R�b>�i&>B��>B�?�_0?oSd?�'�>��m�Ͼ�'��P�>��=O�>��=�B>k��>��7?��D?��K?�~�>Ϟ�=	�>��>�,��m�4q徃ɧ�&_�<=��?_ʆ?���>��Q<�{A�����c>��ŽUu?oR1?�l?��>�	�ٿ�s�)�.�܇���=IѪ=fn���f���K���ʅH�oZ �>7�>���>�wO>~�F>�=NG�=JC�>�,=V����������=6�=[�i>L�P����ۆǽm�p�֢��4��<f������<'n��_W���ͽ^��=�>��6��q�>TkS>�	��#�=Mm��d���y`=����EJM�����X������ڽ)	X>?�u>ɐ��E���$?Kdg<!>�X�?͗�?0��=�z�(=�8ÿ�al>�н׊u>� L>����%	?���U��f����@��>�ߎ><�>��l>�,�]#?���w=��Bb5�l�>�|��~��)��9q�3@�����li��ҺՠD?�F��a��=>"~?�I?M�?͍�>����ؾ~;0>�H��#�=Y�*)q�2h����?'?��>�쾣�D��H̾���g޷>f@I���O�}�'�0���ͷ����>����,�оv$3��g��������B�ALr�R��>��O?~�?3;b�W��LUO�����(��xq?�|g?��>$K?�@?!$��z�8r��Kv�=��n?���?6=�?>>~?�=���>��>T\	?� �?�ϑ?�Ms?��8�k�>��^;�'>V����*�=�>A�=P�=��?�	??

?�����	��B�B�ɗb�� �<��=��>7w�>��j>ú�=�z=0B�=�[>8{�>�_�>��f>::�>�c�>�'��$9����>���=���>� ?�vK>���=�,��פ�$=fᅾ?ݦ�ˉ0��Ni�,�=��=�>w��i��>3�Ϳ*;�?�m#�
u�B�?���\o�����>7\�>O�8�QA?���=�>�>��>�,�>L�=�}>�/�=BӾ�}>'��/n!�(.C�AR��Ѿަz>����c%&���k��eBI�Qf��ed�{j�#1���<=��?�<�G�?������k�O�)��x��_�?Y�>Y6?*݌��戽 �>&��>�̍>qC������5ˍ�#p�^�?���?�9c>��>E�W?�?e�1�j3�luZ���u��(A�oe���`��፿����-�
��
����_?��x?�xA?�N�<9z>���?��%�Zӏ�;(�>�/��&;�wK<=�-�>�'����`�n�Ӿ��þ�7�~FF>�o?%�?�Y?�RV�e0�=���=c 9?��Q?
�:?� W?�(?�
:=�?��=_<?�5�>�+?�L?���>���<b��=a�=��K>T���y�a��DR��b+��<C>���=��.>����n�< q;=]��+#f<���<��Y?�w���{R�ō(=�C�>2�]?�#�>S݅>��6?�o�7d8�@b��t�/?�{C=,悾�����v������>�oj?a۫?�Z?��c>��B�3C�Z�>��>e'>L,^>�)�>@�7I�*_�=��>�o>�&�=�'\�ѵ����	�'�����<��#>���>&t|>�э��'>�����Zz��ed>|�Q�d����S�I�G�4�1�Dv��c�>��K?��?��=�B龼N���Cf��)?�T<?�KM?�?���=a�۾��9�S�J�Z^��'�>�ȫ<I���Ģ�G����:��A�:��s>ڞ��k��	'8>�k�y�޾�Es���I��⾻O�=���=�
�Y�Ѿ��i�72>���=:x�����0�������L?4�=7*���l�l�þ��>��>dͽ>�S/�S�˽��>�3����r=@��>d7>�M;:�꾘I���
�W��>�I?�`d?<\�?r���t�-[F�4#�.��kmW;�j?V��>0�?6�b>W��=������d�ܽK��!�>�r�>���V]K��b�������)�P��>-r?�(J> �?*xB?n?6)V?9L"?L�?��>�;��Y����"?y��?QG>�K�������M�-yg�)��>�K?�=���>d�>ק?��#?��Z?��<?��]>h�.�K�_��>wۓ>�9U�:o��NPA>NX<?y�b>"u?u^�?W#�>��%�1������n��&>�59?�,?�/?���>`�>g¹�Ʒ$>���>��R?��?7~_?9'>��?y�E>��>]��=�ԉ><�?�,?	B?`T`?��;?���>@��;�H������������E���7=�����=F��<aٜ<{���P��=�f�<�y�����vt�;at�;J0�������_�>_�s>v
���0>"�ľ�O����@>b���P��[ڊ���:��޷=���>��?���>�X#�ⷒ=1��>eI�>E���6(?��?�?��!;�b�I�ھ;�K��>8	B?m��=��l�������u��g=��m?��^?N�W�l&��O�b?��]??h��=��þ{�b����f�O?<�
?2�G���>��~?f�q?U��>�e�+:n�*��Db���j�&Ѷ=[r�>LX�R�d��?�>o�7?�N�>/�b>&%�=iu۾�w��q��i?��?�?���?+*>��n�Z4࿌������Fa?�>�>P���|*?Ь�F!ξք�D���'�u֤�}N��y���xK����N�l�2޷�>"�=p�?\Hq?-�q?Z{e?���q�c��^`��ҁ��J�W��(���8�.�6��gL�ȹq�\�qZ�fc�����=w�w��+A�^�?�]"?��8�%�>R���_�Iž�;>�̠�2��u=����*Z�<�kf=�P�.��Ư���?@3�>�6�>C?~�K�x�>���4�=����G>�T�>qp�>e��>^vT��qN�4��(/׾r+��S��� l>�i?�:N?g�j?	7�.�0�H��[�*�����>&����H>�i>k��>k�E�h�4��-,��N>���t�#��K���X����=j�4?�Bp>ݢ�>��?��?��������B��h�*�Ͷ�=�a�>0n?,��>,8�>���-�#����>x�l?>��>��>Q����Z!���{�X�ʽ�!�>�ޭ>Ƹ�>y�o>��,�6"\�Tk��Ǆ��V9��\�=��h?�����`�$�>�R?�C�:jH<��>L�v�+�!�E��p�'���>�|?���=��;>/}ž�"���{�I:���R*?��?6	��^I(���p>��?͡�>�!�>{�?���>�B���	 <�?W7Y?�&K?tKG?A��>�\=�����gʽm|*���8=۫�>'Z>��=�>Ѧ��}�k&�֡=���=�OS��ֶ�\h�;���]9�D<:�?>�ٿ[*N���ھ������
��������h��R/�������`�}5�?�4��FH��[Y�rD����{����?d��?��͍�k���/������z�>�k������Q�����]n��)�Ѿ2���zy�y�G���h��`i��B?�jF�hƿ�~��&�ž� �>��<?���?�e���M?�l�S��|�>�>Ŏ)��BӾ<���[׿=�����Z?��>@쾙dS=�TA>4�L?Prd=h�q=u���i����>�-�>=A?�%�>�����տuB��u��<���?<�@�|A?��(����BV=T��>&�	?7�?>�S1�5I������S�>�<�?��?�|M=�W���	�e?��<��F��ݻ��=�;�='D=�����J>T�>����QA��<ܽص4>)م>��"���R�^�g��<|�]>A�ս�4��5Մ?,{\��f���/��T��U>��T?�*�>T:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�����{���&V�}��=[��>c�>,������O��I��U��=�o��#ƿf|$�V0�l��<��I�?�^�Nܽ�����N����{�p�`�ѽVt�=sz�=��R>,i�>�VF>޾L>t�X?Lh?�Ѻ>/U>i3 �W0����ʾ��Y<	�}�����]������&��`��A侲�������Wξ�7��3���BN��d����@�%a��71���G?�c`=�$�^�(��0<�2��`�V����]��<�ܫ���E�_6�����?v=?^���a�Q ��;<V�漷�[?�ڽ�$���¾��8>����J� ��l�>�C>�h��=���a�}�1?��(?�7���z���>���0_�<TV2?�?W�a=@g�>�?)?}��:�8h{>[x>ǽ�>���>L�>
%�����i�?Og`?����"ኾ �>����㭾O�=K��=}Z��9˻g�f>Cw�<o���Rټ��뽕_0=�(W?婍>��)���c��"/���<=��x?�?�9�>�vk?��B??ޤ<�d����S���ww=C�W?r%i?��>6���$о�l��ݽ5?��e?��N>q[h���k�.�?U��+?��n?�Z?~���Tt}�O������o6?_ʄ?��J�N�����5I���U�=�
?��>>*���>Y�?ߺ�,���p}ȿ� .�h��?�@9"�?���=���Y3>�+?��>х�C�����<� ��{ӼE,?�����1z�Vx5��e��"?��?;3?jc���C%��x=Я;��j�?��|?&9@�l��=��5�Y j�?���ҳ��|޼���=a]7=��)��b�<�ʾ����F��H�=&H.>�@�YH���?���������ؿ^�v�䐼�G�����>��>8u�=�ǽ����q��C5\��OY�in"��5�>I�>��������{��p;�%���k6�>����Ԉ>�S�u������ܦ7<�ߒ>���>c��>L诽������?O:���?ο쪞�ĝ� �X?Qc�?�i�?ul?}3<�w�^a{�l=��G?o�s?Z?�N&��f]�ݓ8�ſj?'`���U`���4��EE�U>�"3?�@�>h�-���|=>O��>v`>%/�эĿٶ�t������?���?�m����>G��?�t+?�j��7��PV��l�*��30�=A?e2>/����!�0=��ђ���
?�0?�y��/�[�_?(�a�O�p���-���ƽ�ۡ>��0��e\��M��)���Xe����@y����?M^�?h�?��� #�b6%?�>^����8Ǿ��<���>�(�>*N>>H_���u>����:�i	>���?�~�?Oj?���� ����U>�}?1$�>2�?�u�=�a�>�a�=�񰾱+-�Ii#>� �=��>�ݠ?��M?�L�>�V�=��8�%/��ZF��GR�@$���C���>$�a?[�L?#Jb>n���2�!�r}ͽ�c1�Y鼖V@���,�ݕ߽4+5>t�=>V>��D��ӾH1?���&oѿ-���v�>r
�>	�!>�-�>$L��(5��4h��)8?۳�>�J(����M���Y.˾Q�?��@�9?1�׾ �P��>��>��
<���*��dk�Z��=�6?:N˾�ȡ�7��&_�>��?.� @���?$AY�:&?~��Zn���z��Q��fv���>*�$?��۾�e>?F�>ЉT=�G|��C��l^i�	��>Z��?[{�?}�?'�d?0�Z�Kr(�Ǆ*>0�\>vN?�%?�W̼T��IHg>�6	?�lҐ��>�YY?�7
@��@��U?�H��	H��<��������̽I�>�Bj�2H3>a����7��ڼoc�=׽ʢ�=���>irg>C`*>l�W>RB>���=��|��Q ������u�b�9�Z@1�x��ˇk�tS��㙾����Ҵ��)�0�=��� ���`�=�"���l����=ˣU?�R?�p?g� ?Ow�i�>����0W=X-#�'�=�6�>�o2?�L?Т*?��=����~�d�2V���(��߇�hi�>1�I>W��>�O�>��>�<�+�I>��>>�f�>-N>�Y(== ��Q�
=��N>TA�>��>sq�>�>��@=j縿����w�����s)�=x��?����/E���؄��B��W�}�>��8?�"�>,����ҿ�����7?�7���7��ǁ��L�=i4=?��^?�?>J?��O�������!I���ͽ-��=Y]�=9f��I�L��R�>*?��f>�u>#�3�j8���P��m��	�|>p;6?�ڶ���9���u�C�H��TݾxPM>�Ҿ>sZC��u�����+�rci��|=<r:?$?���{䰾�u�<,��orR>�:\>��=�T�=�lM>�~c�0�ƽJKH���-=�0�=Q�^>HU?NH,>Cˏ=p̣>�`���O�)_�>{�B>�,>�@?�%?b����������-���w>�K�>5�>^O>JJ��r�=�o�>~�b>��v\���:���?���V>E$~���_���r�<}z=�P���O�=�P�=�� �xk=��'=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾT��>�h��j��xE��1�t�GV#=5=�>��G?�P���O�Z_?�@x?;�?{�񾜟���ɿ��v����>��?{Ŕ?E�m�&ؚ�@%@�e�>��?�ZX?�-c>|�ھiuV�.7�>@?BBQ?�<�>o��2&�q�?�̶?;�?�ג=�p�?'Bw?Pq�>��μ�v9�)¿kߖ�CP$��a�=H�>Y%{>7��i;�����锿Bhj���.���=Z�=mh�>�@P��^��
}��
��@��ʿL�Ք>0ܙ>V��>��F> �>}�0?��?�B����;�J��hھ��K?���?[���0n�s8�<~��=\�^�((?OK4?��Z���Ͼ�ר>��\?(��?�[?�i�>����=���濿�}�����<R�K>�9�>	G�>+���PK>_�Ծ�ED�}m�>'Η>�ǣ�,<ھG*��E.��g=�>�c!?ڍ�>(ٮ=ۙ ?��#?��j>�(�>CaE��9��X�E����>٢�>�H?�~?��?�Թ��Z3�����桿��[�t;N>��x?V?sʕ>b���񃝿{kE�>BI�<���^��?�tg?rS�0?<2�?�??`�A?{)f>؇�)ؾp�����>��!?���A��M&�T��~?�P?���>�5����ս]Hּ���z�� ?)\?�A&?��
,a���¾`:�<F�"�4�U�r��;I�D���>�>����
��=�>pհ=Om��E6�T�f<�j�=K�>��=�-7�s��#�3?�WQ<¬������Oh�:�O�ڣ�>��N��D˾v��?3"�F�������^����V�+@�?���?��?0���G�u��8E?a�?���>En�>�Z8����Q���þ�1��vc.��l�=�}�>/Z0>赾�����z�������q9�<Zn�v?�n]>�I�>as�>t4�>��>0g���F���߾���������=��3�ڄ5��k"�m���ڼ2p��Dʾ�>����>"E^����>h�?��>��>��>�r4�I�?���>���>#B�>��H>���>��>��<����� R?\����f(�#�߈��~A?�Ld?���>��b�n񄿰�� ?���?"ۛ?�zp>�i�}<,��.?� ?�}�,	?��;=�~?�V��<�`���~�6���-Տ>�Fٽ��:��%M��g�s-	?�i?A���Fɾ�UȽ����z�w=�C�?j)?�(�,�Q� �p��W�|�R�7��*+i�/񟾪�#�Z#q��K���Z���*��t�(���.=��)?�R�?#��V�����Nl���?���e>��>�ޔ>��>�H>G{	�"�0��N^���'����4��>7�z?���>�L?�y@?p/O?��>?�V�>���>&��w��>kn�=p��>��>{%8?��$?�3?t�?��#?�;>oƽ-W𾏸��?��'?��?�[?`:?�Z��$-�*y_��t��f^9��;߼�B�=��<"����;s�<=�[>8J?ei�Ӫ8�T����j>��7?���>���>�+��a)����<l��>�
?V6�>� �yr��T�Y�>f��?���G= �)>��=�a��ԺʺII�=g������=BC��8i;���!<!߿=��=�o�	�����:eA�;��<`t�>;�?^��>gC�>u@��Ʃ ���/e�=)Y>�S>�>�Fپ ~���$��o�g��\y>�w�?�z�?T�f=��=j��=�|��U��i������J��<�?J#?�WT?���?��=?�j#?ִ>�*� M���^�������?_!,?���>���7�ʾ�񨿣�3��?�[?/<a�N���;)��¾��Խ��>�[/��/~����D��ۅ���������?���?�A�F�6��x�鿘��[����C?�!�>�Y�>��>D�)���g��%��1;>���>�R?,��>�lR?�{?b�Z?�\O>�L8�dܭ��������=">��>?�&�?��?F6w?�-�>3>HT0��o�!��]C�������~��Y�=i1T>�֒>(��>�]�>T�=�Ƚ�n���;���=�p>r��>o��>��>}�w>I7"<��I?��?���*q�m_��e)��*�]�.{y?Oj�?0�B?��=��!���:�%㾧��>�?�?J�?׼?�}v�) >�mf�լ��A]�m��>�G�> ��>髾=c�=��=~��>,6�>!����')����z��>��<?Ǟ8>�ƿTu��H~����J��A����\���z���q����=bN�����xU����=��������Tð�ZǦ��҄�s[?D:�=��=$��=
����� �<�Y�=�n�<���<w�'�v� ;���'�<z�ս��<`�=a��<��(�uTݾ��|?D-?6?[p6?`��>bg>�z�e�,>�:���L'?�
>㰽ο���Y�����b�P�~
��4��E�]�x"���G>����;>�BA>z|=�^=L� >�� =��=|%F=&�=֎>�t�=5*�=Y�=���=6�>�6w?L�������4Q�VZ�m�:?9�>Cz�=o�ƾ�@?��>>�2��ė���b��-?���?U�?m�?�si��d�>���Ꮍ3q�=繜��=2>���=�2���>V�J>у��J��D���u4�?��@��??�ዿˢϿ�`/>�
2>\�	>}hR��*1�$X[��<\�i�Q��- ?�u<��f˾�|�>jή=��ؒǾ�=+�1>wFt=���ԔZ��o�=�F~���G=�Bj=/�>K�E>��=�ۋ�=T�K=g5�=\�V>��x;��/�Ǫ�6�B=���=�;`>�h(>���>��?^�7?DGb?cN�>�
���	�g}ľd��>�/>���>��=X��>�7�>5�<?PJ?��G?Hʑ>S-��6�>��>�j0���x�TM�=ط��:���?���?���>^[s<�����#���<���½�s?��/?��?(�>���t�׿���Ҿ�/B�y�e�W<)UK����;���������0u=
N�>���>R�>��>�N�jG�=<��>�'H> �I<�5I����_��=ݐ��=[&>�D==���=վ(>Χ<��A>��ؽ�$H����=�����̽���օ�=�v�>���=�B�>}�=����;��=4��
\��4�=���'Bq�㑄�I�o���(�}���8Rv>* �>Խ��Ǖ��?�E�=�ƍ>"��??��?Q��=���=�ݾ8T���dL=����w4>ȗ�>&����P���n�^�N������>�ߎ>��>�l>�,�#?�*�w=��wb5�-�>�|�����y*��9q�@�� ���/i�X+ҺѠD?�F����=#"~?�I?H�?B��>8�� �ؾ�:0>
I����=1��)q��h����?'?Η�>��o�D��H̾A���޷>�@I�'�O���P�0����0ͷ�/��>������оq$3��g�������B��Lr�k��>(�O?��?T:b��W��?UO����^(���q?�|g?"�>�J?�@?�%��z�r���v�=�n?̳�?Q=�?a> �=[^ýYG�>5�?��?��?W�r?T?>��{�>HԮ:�&>L���{�=�!>��=�Q�=�;
?O
?��?�Z���=
��>�*��]�Y<�<���=kA�>�o�>�1l>�_�=>�M=���=a�d>be�>&;�>P7b>˜�><T�>���*Ҿ�?�1=d#>VP?�kz>�H�=.h��Q�T��=�U��w�!���Z�L���׻��>���=��.��$�>\Vɿ�Q�?O�>_��f?�����D��¸>��=>9����>��>${>	�r>�+�>z��=_�Z>vp���EӾ~>���he!�y-C���R�O�ѾB�z>T���n&����_y��*@I��m��f�0j��.���<=�ݻ�<�G�?���9�k���)����{�?�[�>�6?Wٌ�"���>b��>�ȍ>�J��}����ȍ�h���?N��?�;c>g�>\�W? �?�1��3��uZ��u�G(A�e�A�`�n፿����
�����_?�x?"yA?VP�< :z>K��?��%��ҏ�(*�>�/�9';��;<=�+�>�)����`��Ӿ�þ(9��GF>g�o?%�?AY?�SV��h>�{��n�R?��|?��J?g��?��1?�s�<�?w8f>�`?�:?�!?Va?�-?��>�M>N%��-�9=v�;���������Jc��I=M�w=�=�=�'�c��BI�>;c=�K�` ��G��=�K�=V�;�W��=۞�=ɼ>i�l?r� ?��Z>�l ?�D>��L?� �e���P?�/>wuc��t��畾2D�mH>/�?# �?`.H?��P>��9�SuE��=>�@�>rU,>"�s>J��>(ɽ2ᗾ�{�<9/�=bO�>;Z�=��~��t{���\��/�?��]V>���>R+|>x�����'>*}���$z���d>K�Q��ɺ�W�S���G�.�1���v��U�>}�K?:�?���=p\�A1��rGf� 0)?$^<?�PM?�?�=�۾��9���J�8���>���<���V����#����:�j�:�s>q.��
k8��>���hо�n�ܝ7�J弾�&>�U�]����#���:�=]��=�������aN�����UES?��3=-Ρ�r�e�Z��	�>~�>5$�>7�����ڽ�9�����-2��C�>'�i>�������� \E��?���>��-?Iha?��s?=V���a���b�\��3���qD�=��6?���>(�)?�#�>�[> �������}��c��1�>�M�>��
�z&J���ھ4"9��09�M��>��?�9�>U�?��&?��?:S?
9?��?`�>Mv��ـ���?ײ�?�
>�e;��ɾ{�|���z��?�}r?[�0����>v/?�0.?�?h�]?p ?�=T>��ܾed�v��>}c�>>V������y)>)D,?���>���?�$�?�3>%�g���ƾZ<M����*B=?�ZD?�`Y?o	�>jW?<�;��K>N��>�+I?DY�?��e?Ų�=t�?'ne>���>,s�>��>�`?&?�t9?��b?	�-?��?���� �j�^���������
V=|�Q>sEv=��1�b4��4&���e'�@z���*>yGD=R	νYY̼C"���s=���>��w>���;
5>�fľ0���GA>��8*��F�����7���=�P�>��?hٕ>�~"��3�=Uܻ>�?�>��bb'?��?�?@g�:�Ia���ܾd�K� ��>�9B?�o�=�1j�ꝓ�I u�O�{=�*m?C�]?88Q�"���O�b?��]?5h��=��þi�b����c�O?:�
?0�G���>��~?a�q?R��>��e�$:n�&���Cb���j�Ѷ=Zr�>GX�O�d��?�>q�7?�N�>-�b>>%�=_u۾�w��q��c?��?�?���?+*>��n�T4࿧����L��J']?��>hY��$1$?�.��ǐξɗ�'팾j�\X��eq��f�������y��C�r���˽�p�=��?�vr?��o?�]?����=Pf�K�W�Z<v�)�O��j�����8��J2��G�B�p�^Q��P��=���B=R���8I��Ӳ?�?Ӑ-��I�>s������׾*C>�����7�C�=�8��,��<g�=�eQ�&�%�����_�?
޵>���>��<?�TW�,>?��.�Y�3�aW���#>��>Ct�>���>d-���>��v��޾�������->�P?��K?��M?�H�J-�; ���jA� jV�����U'�>���=���>ˬ��m�?�]e7�2A�6���o�!�ލ���!���zE=��I?�R�>�g�>Օ�?"�?�ͻ���L׃��h�� >�߼>�Fn?�y?6{>�x����2��>�l?���>���>Ť���^!���{��0˽��>dܭ>0��>��o>y�,�\��n������L 9����=z�h?�p����`�H�>�R?Ew�:�>H<�o�>�kw�غ!����Ϩ'���>zi?1ͪ=P�;>�rž��k�{��Q��6h#?��?�C"�n,��>ԓ?�`�>��>�<�?�-�>�/����I���?�gQ?>�W?յ7?���>��;�}<�-m��=17�X��=ѧ�>=0V>;�=|�>W`�׵c��;�	\�=�A�=�Mc��C�M$Ż���'�����a[�>7�ֿ��W��z쾷;����,;˾V���b0�	c8��1 �9ľ¯I�����ә�k+���r��"������,L��0�?��?�6�ң6����Q�J��-⾒�>�׽���z���v��Y\�T����پ����ܾ��+�]\���M�o��>����Rٿ���c�a�>��F?���?����,Y�ٻ4��wy>N9=}�h=]��i䚿�ٿ��[�Zg??x�>�n �#>⽡��>aa�>B��9��s>�S�xν�;#c>���>�B?>�4?�a;Tۿ����hm�=��?�@bA?$U)����h�U=ut�>��
?2�C>3�0��I�����[��>|�?~��?��`=�JV������d?�#<&�D�E��X��=U�=&M=1�>RH>�ғ>�?���F�&��"/>�T�>�8���fh`�5ۘ<Y>�u׽���4Մ?({\��f���/��T��U>��T?+�>Z:�=��,?W7H�`}Ͽ�\��*a?�0�?���?#�(?:ۿ��ؚ>��ܾ��M?_D6?���>�d&��t�օ�=M6Ἑ���{���&V����=Z��>_�>Ƃ,������O��I��a��=�����ȿ��`��IO�<{ �<?���
����{�?��7��w7���:$� eM=��=w�m>·>r�N>�\U>z�R?�a?T�>�h>G�
�Kv���ɾH���Ɩw��>�+$��,u��m�)��C�)���&��k �B��SC4���t=9�`��^��ظD��g7��*G���;?�T�>���z�B��S$=k蛾�������;8�=�ؾ�_=���a�"%�?�TK??ᗿ@�i������
=���e}?�&=,PF�f�þ��,>��i��y�3��>�Q�=v�6b2�h�i���Q?ȁ3?󛇾��A���$<(Z���r:��?kS?��n=�i.>0n"?�΅�A�7=H�>��>��>D߲>�.9>�ľPd%�_P?�;??������e�>aɾ�Ɖ����=�^>咽���>���=��L�γ��P����
>� W?��>�)���|o���s�f�<=��x?m�?@�>>gk?��B?KȦ<�\��4�S�H�91x=3�W?Si?V�>T���7�Ͼ�l��V�5?��e?O>H�h������.�IV��"?��n?tY?�����p}�������w6?�_?�ǉ��m����!�(�e��}�<��?�^>]�7��,?�y�>Z�þ�J����̿6B��ͼ?ʐ@�@�`��O\�2WN>�'?��>AM��<�C�=��<S�=�?�����m���t߾׮���4?l��?5�?;��D�b��<�����ͦ?�3v?���N�1�/R!�/�`�E	�M&��]�ȼm�}���G���Q����
��f���c<t�j>�`@�ӽ_��>�<_�]��obĿ�_z�%����k��J?���>��>���G|��a���q^��KZ��|���>�o/>pϣ���|�Uoq�s-��x�<��>QiL��|>S[H�f嶾z��06�<�"�>7/�>���>����7��F��?��ɾ��ӿ16����� O?׺�?��?;?�p:�/����щ��jf�Ç7?*a?�cP?�uM��%m�^���#�j?�_��oU`��4�kHE��U>�"3?�B�>S�-���|=�>���>g>�#/�t�Ŀ�ٶ�7���V��?��?�o� ��>l��?hs+?�i�8���[����*�.�+��<A?�2>���O�!�H0=�[Ғ���
?K~0?&{�d.�\�_?&�a�J�p���-���ƽ�ۡ>��0��e\�N�����Xe����@y����?N^�?i�?ӵ�� #�f6%?�>e����8Ǿ��<���>�(�>*N>8H_���u>����:�i	>���?�~�?Qj?���� ����U>�}?���>�t�? ��= ? 5>�喾�)<�%>s�y=��v� �?�E?�R�>�T�=}'$��}&�ϙ?�	M����FtA��>H�\?��F?��a>Խc������˽��,��%�<-���b/���h,>^>>C> yC��ƾ�0�>\W��㿸��<"�>XI�>b�`>"�?˹`�/���Q����?B>��,� b���T\���Ǿ?�O
@c�?R���.>?�>�#?V�� ����<�1��Ѷ	?W�>���Iح��d����><��?9�	@�?�_�c?�3.�o�����y�>�������g>J�)?�sᾙ�>�ln>lr=Mn�����A�v����>��?�u�?D?I�a?�`�R �!��=5*>KKT?�?y�����YX>n?��8��ǋ�;��~B?Q�@*�@�mE?����q�Ө�H婾Ӊ7�q�g>&�d=J��=r��&<_�,�4��=n#>r�q>S�f>�ǃ>|n�=Zs'>'�c>����0�t0������U�6�0r��I'��2��"��X%{��$���������
B�)e��[���3���\����ٽA9�=��D?�,I?�Eo?ô�>e� <:�)=zF�:�)��	U��F.>[a>$ 0?��@?͇?�V<�O��c�j�,k�������u�!w�>��>�r�>�շ>�{>���<L�=:��>��N>4�>��=�s�4E>�e�>At�>*[�>�b>��P�A��=�¿�̿8�������)�C�?A�n�: ��R�������վE�=~�,?��p>�á�_ǿ��6NZ?��B�"9�UP<�>?q�?Fb8>���^`��Xp8>=�E��l��8�>(ɂ��ɾ�j<��7�>�W?�3?}�>�)���@L7�V����>��Q?�>���X���k��iK�����H>��>���9+��S��Js�l���N;�0?�?RI6=1���}�� ��[�>�r>�>���;8>I֦>,�m=H�]�'�m��<�>��>��
?N>Ic�=+��>GB�=��(�>ʕD>�'>ƶ5?yX ?�ڝ�*�h�{�p����K^q>^��>^�>q�>�FV��6�=��>yT>.��������?���j>�N�E�R�,�3� �&=K@z�-�>k�=S�&�(�SBY=�~?���䈿���d���lD?Z+?O �=�F<��"�? ��|H��@�?o�@m�?��	�ҢV�?�?�@�?*�����=�|�>�֫>�ξ*�L��?��ŽSǢ�Ԕ	�X)#�XS�?��?T�/�Zʋ�Bl�O6>�^%?��ӾI+�>�1�%X���D���Rl��!��&u�>	mM?a�Ҿe�ѽ��R�'?p[?�x�ה��aK˿�ր����>�<�?��?�]{��v��$`;�E$"?Xe�?�/?Ɍ>SBӾۧu�H+M>��K?�}F?^�O>7R���
���?Xĸ?�2�?����(y?�g?��=��;5J�n�¿cf��^�۽�+�<�i�>��@>7(��K����Y���@|��G��|�=���=p-~>�O�ml���C�=��<������k��:j>�!�=ժ�>�9�=�v�>��?v�?%U�=���H����Ծ��K?!��?~��n#n��a�<���=�^�%?�A4?�\���ϾCԨ>0�\?���?h[?K`�>���!:��J῿E���SȖ<��K>l1�>�?�>���"8K>��Ծ�2D�;n�>Xؗ>쑣�X/ھR(��A���>�>Na!?Ñ�>N�=ڙ ?��#?��j>�(�>>aE��9��S�E�ò�>ۢ�>�H?�~?��?�Թ��Z3�����桿��[�s;N>��x?V?}ʕ>c�������YlE�6BI�+���]��?�tg?|S�,?92�?�??[�A?g)f>ԇ�%ؾj�����>~�"?�	�I�<�ڞ$�w	�h�?)	?��>�ȝ��;����C�����<�?�*Z?�
"?:���^�������<�j߻�����#�9�E�>5�>��W����=��>��=�nx�E��&":�f�=�؎>��=�?��f���R?o�4��n��]�m�)���qTb�%��>b���;	��*��?�c������M��������腾�Ĩ?P��?�C�?)�,�܋x�sj?�R�?<~D?'�>C���'�2���[J���þ������>˔6>b����<ɾiw��E�������X���螾��>���=Y��>0�"?&��>SB�>��ɾ��n�#��:-��q��rO��^u���8� ��{�P��[罭"3�=�;���7��>^q��ET�>S�>��>���>b��>��;���>��]>Pow>�7?��x>?F>�`C>���=O=H�N?ΡӾ�O�L۾#Ј��M?��h?7��>�B��*j��؅�E?j��?��?��m>��h����B�?�$?�y�	�?\G[;�H����<=_������xb�;�3��{:>�e�@�P���[��v��*K�>���>q�����Ҿk��㮾fF�=V�?� ?<i)��^V���y�2V� JJ���?�.({��Ղ�+��v�s����]����Z����-��I=^?�e�?f8�_ �帾ߜj�nFA���">���>��>��>�e�>��վcK-��t�v�4�荕���>�cj?(֮>�|T?�1?:�P?s��>�>6�>TxO��{�>0�.=?�r>�5>�?;)3?��D?���>��>'W>�9�=���r����'
?V[?�n�>F? ��>%߾�R��%w�ʥ=v��D�O�>k��=&`��&H+��+�0�8>7"?P �a3+�����- |>��>?�s�>�(�>��������`<�>!P�>qq�>����o~r�r���>m&�?����%t=�Y>��u=����᪮���=�9{<Te2=���Ԙ9�Xc(�+�<�]�;5d��M��E���Bмj�; u�>,�?ȓ�>�C�>v@�� � �T��lf�=�Y>S>u>�Eپ�}���$��j�g��]y>�w�?�z�?��f=��=��=�|���U�����7������<ۣ?AJ#?1XT?c��?��=?Xj#?��>+�aM���^�������?5�-?��>����~Ǿy���h2�q�?��?�m`��
���)���¾]Խ��>��.�d}��P���pC�Gܡ�Y��������?p��?>��6�������^����C?�C�>'��>b��>q8(���f�����j;>���>3�R?�`�>��N?~�z?��Y?j7N>�8��2���^����W�W�>�A?L��?�n�?(�x?�Z�>�>'C.����V�����$�����1N���Ks=frX>�Y�>��>^��>K�=�ĽM`���D<�Hǵ=?_h>��>*L�>~
�>�~r>�̺<0�<?���>����;��a���d�����㴂?� �?�e1?9�?��&��V#� ��o�>�,�?���?[�*?�M��D��=�Bb��o��p#V�)�>.��>�'�>��h=�n��w&>�>:l�>~w����{;��S��g3?N=?)>��ſ!�q���n�d�����r<�~��ڄb��9��A~Z���=P���������DIZ�m���gR��~����s����y��N�>�u�=���=ä�=圾<�&ͼ��<�0F=F��<��=�2n�P}N<��?�Qͻ~��M�����a<�I=�3޻x�e�d{?xR>?�A?��G?]�z>T�	>4�����=�2��N#"?z�a>n��������I�a���Q���վ�J��3]���Î�PQ*>���p�=0~�=���=��=0�=>[�=��=�.M;�<�U�<26 >�{�=;>;O>Z^=H6w?�������5Q��[罢�:?�:�>(s�=y�ƾ�@?��>>3�������c��,?��?uU�?��?�ti��c�>����؎��u�=XƜ�6>2>��=g�2����>��J>����J���~���3�?i�@r�??�ዿm�Ͽ@`/>��q>I4 >��Q�A,�L�p���J���7��Z)?��6���׾w��>�ґ=�`��6¾�QK=��,>�bN=���9[���=�����z|=�j=�ڊ>��<>��=<ﺽ�u�=hp=�H�=0D>�0��T3�6�����=뿤=�V>`	>m}�>S?�P0?��Z?��>k���ܾ�#���>Q�(><��>_��=�F�>��>U;?��9?�8?Թ�>�]<���>;?�>oG8�˂o����`׾���;�-�?� �?�w�>��ۻ�c����t?������?��4?�8?M��>�U�z�࿫X&�$�.�ň���e��+=zmr�cTU�����qk�����=�p�>���>�>�Ry>�9>�N>��>Ī>7�<�m�=���ĵ<f��,��=餑��/�<�sż<p��q�&�K�+�v����;Ե�;f�]<D��;�?3�x�>�������>���=`򞾖H>�ܾ,Ug�]�\>�����Ab�b㑿�ՠ�Z9� 7)�:&�>$~�>2���{��5?���h6	>R��?= �?�wP=[���{h�%P��pp�=�F��p>��=I���!|Q��������	nǾt��>���>��>޸l>�,�#?���w=��&b5���>�y��i��=&��7q�)@��2����i���պ��D?�E����=s!~?�I?��?���>���N�ؾN80>�I����=��3*q��b�� ?i'?n��>x쾤�D� G̾
��a޷>�<I���O�������0��o�f˷����>B���e�о'#3�g��F����B��Ir�U��>��O?$�?�1b�5X��	UO�/���)��}q?2}g?��>II?@??�+��Vz�Nr���l�=,�n?��?�<�?�>�>Ѡ+��o�>s��>д�?D��?8sd?����}�>��b=��>��P=�->6�>�˸=y{�= ��>0��>n�
?�s?� ���Rܾ 8��R}���=J[�=*!.>7>*��>���=�/�=�}I=�>r�>��>^>*S�>,͔>�׫��{���?鱨=��>f"?>�T=��$���=n�@>�2����־��+��n�`Џ="�I>��,>78ݻ��>%�˿u�?;����$�?N�����ŵ>Ў�>��"��Y�>��>�H�>�h>J��>�.�=)@>լW>.Ӿ�>.��IW!�k C��lR�߈Ѿ�z>�g��O&�׎��V��I�DP��}Y�`�i�'��})=����<�S�?��� �k�#�)�'���~?Xx�>�!6?w،��Y���x>���>���>2E��<���2Í��Q᾽
�?���?�;c>��>B�W?�?��1�3��uZ��u�l(A�"e�;�`��፿����
�-���_?	�x?(yA?�R�<:z>F��?��%�_ӏ��)�>�/�';�7@<=~+�>*��-�`�x�Ӿ��þ�7��HF>��o?5%�?oY?$TV���=�A>��*?vU<?t�,?Ҍ+?�?�/c<,�O=����#�>��1>�?�B.?�}'?�p�=�m�=����sCQ>u���D���=��a���Zc >�#*�����R>�]�=X��D�<S|�=]Q�=�<¼0!���:��=k�Q=��Z��R�>��\?(��>9�E>�B?�`��Q>�۸N�a�K?��>����"���C�Fj�K�>S�]?Ɦ?4R?:�>��:���T���4>P��>��>�6�>���>�*F��ك��9O=��=��B>=h����}��`	����> �� "�>���>A�>ÎK�9�8>ۚ��Ec���m>Q�7�Rk���(]��B�.�1�W�l����>�{M?�$?�܊=�9�*~X��b�T$?��<?lM?��|?��=��辗`;���G�<��p�>W�A=�|�>ơ������;�Z��;��>*@���8��z�_>q�����m��1I�yP�iT=-����2=���u�Ѿw"�����= �>1����!�h���J?x�=h�����e��j��vs>a|�>�+�>�EJ�u��ȳ?�k���i�=E��>�6A>Br��n[��I����,�y>�7;?��b?�#�?8خ�XQf��R�����I��Fѽ�<?��>�-?z+�>��t>�/i��� �[h��b����>��>�m&�$�a�/ľ��P�7�F��>�?3���>C�I?*�?d�B?2?��?뿍>s��:\�k�1?}��?���=p>�����:b��Od�mC?�^?���h�>��?Z6?�'?^�h?��)?��>�9��_��q�>�
�>��T�����#>2�0?���>@f?���?Ƅ�>,�@��G��������]�6�=s4?=G:?��3?`��>,?Q0��-��>��>Q2?o~?u��?t�>�m->��>�;?l�=�O�>ls"?<\D?@CM?�e?�?x�>
�Z��6ݽ�c�����׫C�h�=9?>�af>f�0>U�%>LZ�4ˡ=��=MR��1�0��ES��!,���4,��_�>��s>�����0>��ľ%K����@>�j��P���؊���:�Nܷ=r��>��?謕>S#����=��>�I�>����4(?��?�?%> ;��b���ھ��K�U�>�	B?V��=�l�0�����u���g=��m?�^?�W��&��I�b?��]?"h��=���þ��b�܉�T�O?3�
?]�G���>��~?e�q?I��>R�e�4:n�(��Db��j�2Ѷ=cr�>LX�K�d��?�>_�7?�N�>)�b>J%�=Ru۾�w��q��c?��?�?���?+*>��n�U4�P�����2U?���>=ڝ�Z�0?��!�	�ྡi��Do�+b辮9��+��mb�2��1�3���_��櫽�">{I?��j?�g�?�X?�A�3�e��^b�����7k�w��c���[/�?�1���L��j��I#�S��(Q�����;�~�ګA��u�?]�'?��/��.�>Θ�Y��̾�dC>�������9��=�s��p�>=�Y=��g�.��í�7 ?m�>g��>M�<?G�[��:>���1���7��z��:u2>ƚ�>���>zF�>?0:8�-��d�~!ʾs���!Խ�d>Ko?yiR?jh?W���kC�i����=����/;'��=nC�=��>%�G�DY<�~Y3��6E����8e��g��[
�ڨA>Z�3?�o�=,�>�<�?>�?�����(l�[�h=��-�渄�x6�>�?{)?q�z>*�f��J��ܷ�>��l?��>L�>%����Y!���{���ʽl$�>?߭>��>��o>`�,��#\��j��M���d9��v�=y�h? �����`��>NR?a�:�G<�{�>ͨv�`�!�����'���>�|?癪=��;>�~ž�$���{�17����,?��?�{���.��C=>�:?���>���>O��?*c�>������=*?snX?�%G?vF?_��>rCt=����̽��%��x=�:�>�m�>�)�=��>�mཌq����%��=&ӵ=��a1ýȼ���h�E�:7t<C?Z>�Dѿ7X�Az�1��,�������L��v(�9�P�`s��ҩ��'�i�m�r��6	2�L����7t�ˌ��R���s�?&�?�|��ž���yJ������>I�.�e�½��+��������Ⱦd�����#�=�C��K�BNe�p�?�R�9ӿC~��g�f=���>aQ?h?N?�����$�W�L��>���,C���۾BF��C⿻԰�C�f?7��>w�����^����>��>�@�=�t¼Ծ��H�zcd>&�>��H?�	?0ܾAuҿ	鳿EÞ==��?�@�|A?4�(����g(V=���>I�	?��?>�P1��K�����W�>V;�?���?1�M=Y�W���	���e?��<��F���ݻ��=K�=�.=���ؔJ>�W�>�|��UA�z@ܽ��4>�օ>͖"���&�^�R��<��]>J�ս�6��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=�� ��<ǿ��$�����Y<d��;����ֽ ���sF��#Ւ��N��>нS�N=���=��g>�w>l�:>k�H>U�Z?��k?p��>vP>|��Euξ�6����l�i{�������߽Qc���徆�վ[L�@s�	��ҳž�7��p	=�{`�����5�$�8�]��z4���$?x4.>��޾�\U��n�= ɾ�w����<rh���߾�1��rw�e;�?ϴV?�Ѐ�;:x�Ի�&fN=7ཪX>?�(���?[Ǿ8��<��#�%��:���>��B=�0�?xL��sP�?{4?b"0?aN������8�=OR&��d;��A?��?³�<�I�>]�'?�%������|~>�f>/��>Z��>���=j���-۽��?�g?������t�*��>�վ2�ھ=�>�N$� #9=U>2�k=\a��e��=�����=�(W?���>Q�)���c��k/��$==K�x?�?�,�>Syk?��B?��<!`��j�S�����w=K�W?�"i?ϲ>7�����Ͼdj��b�5?T�e?��N>Chh�����.�Q�"?k�n?�[?�3��u}����W���q6?��~?�]��<��ж�<ჾ��>"��>:F�>��&�Α�>��!?��Ծ�ܡ�s�ȿ�;��`�? �@a@��>�$�����=��.?Y��>K9����x��T�)4ƽ�?�tƾ�G����Z����-�?�^�?�?����A�.�:��=VS��R�?ǲh?�܏��(�=�V&��2��n^'�:���C=91����伱$徴�I����b��x��k�H<�G�>�r@m�=��?\ 
����yο�y���_�$-?���>�t�=�d�'ċ�$���!h�0�P�jo���M�>��>����:���J�{��q;��&����>c�k	�>L�S�-&��q�����5<�>��>��>Z,��R轾3ř?�b���?οs���͝��X?h�?�n�?q?��9< �v�^�{����-G?��s?MZ?�p%�#>]���7�h�j?S`���U`�u�4��GE��U>�"3?�@�>��-� �|=p>݆�>�a>�$/�0�Ŀ�ض��������?݉�?$o�}��>���?�s+?�k�8��XZ����*�S�/�=A?�2>�����!��0=�7Ӓ�{�
?)0?&z��/�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\� N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>eH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?x$�>�?�s�=yb�>�`�=P�u-�Sk#>u!�=m�>��?)�M?GL�>�Y�=~�8��/��ZF��GR�5$���C���>G�a?�L?Lb>[��2��!�?}ͽd1��>�DW@���,�m�߽�)5>~�=>>U�D�Ӿ=�*?8���߿�����o>	�>��$>Z-�>����P�uY��q?,W>�?�*Ǥ�yK����q�4��?`�@�.?#��<��=���>�:	>t�=@�<�f)�s�׽��m>�N?�9Ⱦ4��i�q���>M��?�{
@��?�K��+?L<��o���t�B�Ӿ��a�6�
>&�#?(�Ǿ�1�>�%�>Ӕh=~�u����k����>���?�H�?��?m�c?��g�1r��G>+@>aT?}�?s?��AA��/>G<?C�B�*��S�Q�M?V�
@y�@lh?�:��D�տj���̧���-���>$4O=!��>��=�.�=R,:�I8/�	>���>X#�>~�> �2>cA0>L��=Q��=�������U���HL�����܈���5<��ھMG��Q��:֛�c�����͠h��ɽ+&�
�I�4��E:�=��R?%Y?�w?���>`_��ΰ�=^}��F�J<o�-�T��=��Q>�=.?�G?'?�q�=�ݯ�y�j�]��o����
��b��>��{>��>���>�>��.=Y�B>��[>��>��&>'�=��=+��=}qk>��>J��>�¬>�� >��$>a���P޿��RI�]b��p���Ք?�q���zZ��䔿v�k�8��$=n{6?&|>�H���Uпu!��4P?(?���#�Lk��|:�>3~#?��Z?��>�S����p���>܏2��ӌ���=��ѽ���Q�E�B>�,,?�f>�u>֛3�e8�v�P�}|��j|>�36?h鶾=D9���u���H��cݾJHM>�ľ>�D�l�~�����vi�;�{=\x:?ل?�6���ⰾb�u��C���PR>w:\>U=Li�=�XM>ibc���ƽXH�g.=��=�^>O?�+>�V�=�0�>�0��N��a�>C�C>�d,>8	@?�|%?����)H���H,��w>��>3߀>i�>��I���=5U�>��_>���ł�{��U�=���V>�x�~�_� �v� v=����=��=���=����x�=�Y� =�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�h�>�x��Z�����;�u���#=@��>8H?CV��K�O��>��w
?r?�_�թ����ȿ�|v����>��?l��?F�m�7A��_@����>|��?�eY?�ki>�e۾�[Z�ъ�>��@?5	R? �>�9�m�'�1�?M߶?m��?V�]>9{�?�8o?\��>^��<a>���ǿ�d��r�
��ו�$��=�C>�eӽ|�/�2ǰ�`���Y�u�!
9�ɬf=#�[=��> ��/Zs�;p=E1d�(�q)Z����>�e�>�t<�V�>SU�>v�>Ӗ�>�m>>�����e���?¾�K?0��?i���;n��w�<�ӛ=��^��7?��4?�vW�ìϾ8�>֭\?���?�[?���>����*���࿿�s����<��K>��>�S�>�:��%K>4�Ծ��C�B��>���>J,���rھx)��5t���)�>�m!?L��>�4�=ԙ ?��#?��j>�(�>8aE��9��f�E����>���>�H?�~?��?�Թ��Z3�����桿��[�A;N>��x?V?�ʕ>W���䃝��kE�wCI�����\��?�tg?�S�$?:2�?�??Z�A?)f>��ؾ����>s�!?�l��jA���%�9�(�?��?R�>����ӽ�Ǽ����d��k,?m(\?�7&?�L�\�`�n�¾���<����U�LU�;2�K���>�o>C��@�=�>��=wEm��O6�;Te<з�=�>҂�="�7�(落�2?O��n����P�=�����i�N��>2����о�B�?\8޾99��˙ȿn��G���u��?���?���?|���Q�u���^?U��?���>�"�>�a�r@Ⱦ����ہ��Uݽ'�C�~��=k�>J��=����ԭ�CS��&����;��A� �?�
�>���>nZ�>K<�>М�>`P̾��,�A@���ɾ]zr� z8��T�R<�&��	�>��zK=� 	=��ƾ����>*˖<$\�>y�?#4>/[>�6�> ���!��>;��>���>�O�>��>�т>��=TS��7|�uKR?������'�������x4B?�rd?2�>�i�"������?���?qs�?B@v>�}h�,+��m?/>�>��p
?D:=���G�<lW��Z��A��%#�8��>�=׽�:��M��gf�2j
?�-?/1��u�̾;׽�B��&;r=J�?��(?�)���Q�G�o�0�W��PS�V����g�����=|$�ҙp�1������6��ޚ(���*=�n*?-�?B�v��)ꬾd_k��O?�.�f>�I�>�s�>@��>uQJ>�Q	���1��X^�	U'������]�>b�z?�®>�R?�*G?�(S?��$?���>�>�ky���@>a���B�>���>6K<?k�??0Y=?J%?'�(?e�I>�۽��پ�����.?
?�k?��?Q9?H����ԾI�P�/S=OZ��я��՝
>c»��	�j=�n�=�>�X?̙�v�8������k>��7?���>���>���-����<}�>�
?}G�>�  ��}r��b�nV�>���?���ς=5�)>#��=�����Ӻ0Y�=�����=�9���x;��e<{��=���=�@t����b7�:���;k�<�s�>U�?[��>�B�>x?��� ���[_�=�Y>+S>1>Hپ'~���$����g��[y>�w�?�z�?��f=��=���=�z��(T��#���������<|�?�I#?�VT?�?��=?�j#?�>�)��L��{^�����d�?w!,?��>�����ʾ��։3�۝?i[?�<a����;)�ߐ¾��Խб>�[/�i/~����>D��텻���W��6��?�?IA�W�6��x�ۿ���[��{�C?"�>Y�>��>U�)�~�g�s%��1;>���>lR?r��>��O?�D{?"\?]�S>s8����j���*s9��c!>hX@?ݒ�?t�?��x?6s�>I>̌*��������o��W��T(��o�V=�Y>�>���>P�>F��=��Ƚ�
����:�x�=%'c>���>�ѥ>�K�>��w>0��<BMK?�	?�Z��9��F�־%������{?pH�?�J+?o�/=�c�z.�.aҾ'�>���?�ת?2#?7����=W��.����C��]�>���>�!�>���=5Q�=�NA>2�>���>�{���
�N&;�����e?�q@?�]>��ʿ��{��f��d��2eF=�~�2E�ߧ�u�H��"�=��p��������G�*��;�l/��~��������>�(=��=]ߔ=��C=��<�s�;G�Y<Ļ�<LЅ=��(�IS�<9	e���E< ����=�;�<#��<4�<�!y˾7�}??DI?��+?�C?m�y>Q>2�3����>�����D?
�U>TP�Cg��oS;�����Z8����ؾ�׾�c��ӟ��L>�H���>Y3>n�=�܉<��=��s=�~�=�gF���=���=���=���=��=��>P>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>I�7>D&>��R�ڈ1���\�;�b��{Z�O�!?5I;��G̾�9�>���=�.߾�ƾ�m.=�6>�pb=�]��S\����=V{��;=�l=jՉ>��C>zu�=�,����==�I=I��=R�O>�4��Jn7�9,�8�3=���=�b>�&>��>�.?�g0?�d? ��>��i�"�˾X���׾�>�o�=4�>�P�=m�B>��>�8?�D?%rK?���>�%�=i��>&]�>l+���m��G�X0��f��<ˈ?`�?�˹>Z/O<�XC����(�=���½�3?6�1?�?�9�>�_��P�K/�Œ��F=�ڔ>��t>qX>`�<2
;���;W�����=��>�B�>�O�>�W&>C��������>���=��B�����'����'�ս`<��啽�����$�=��=}�=���g�>���=Y��V��<靔<�t�=�Z?�=H��R�>Z�;=XӍ�4[J>+ƾQG��®>8�D����X��W�V�P��𚾲!�>��>{p�ё�$�?%�=>�H�=2��?�Β?�Ӽ<I[���4ɾ�5��e��=|�8�6d>2�G>L�M���3�=�O�Q�A�Mդ����>]�>J��>Q�l>�,��?���w=��b5���>�����P�C�R<q��@��m���Si���ȺZ�D?�E��B��=%"~?��I?��?5��>x4��J�ؾ�40>�R����=X�nq�qi��u�?]'?��>��D��H̾U���޷>�@I�-�O���U�0�X��+ͷ�9��>������оm$3��g��������B��Lr�c��>+�O?��?a:b��W��EUO����h(���q?�|g?/�>�J?�@?=&��z�r���v�=�n?ͳ�?U=�?l>��=�(Ͻȍ�>;�?k�?߬�?x�u?��,��n�>�@�<Eu]>����m3�=**(>�#�=�|�=��?�?m�?�����z���������������<�>�̩>4�>⸑>���=0c=>�\=�^>�2�>��>bڀ>�?�>�Dq>����>t�L�?�m=�h>UCP?ͺA>8��pC�W">d�*<����fQ��.0�L�S����;�U�=��#>3�=�k�>��ſ�ɗ?u��= 8����?aD���7��7�>	�A>35��m��>�8�>��?�Ӳ>���>���=B�=�\>�;Ӿ��>����s!�QC�	R�N�Ѿ�z>�����"&�}���q���VI��l���]�wj�f3��wA=��v�< G�?�����k�-�)��O��x�?
[�>�6?Hڌ�9݈�)�><��>ż�>uK������]ˍ�ip��?���?�;c>��>H�W?�?ג1�-3�vZ�,�u�n(A�+e�U�`��፿�����
����-�_?�x?2yA?�R�<+:z>Q��?��%�Zӏ��)�>�/�'';��?<=t+�> *��*�`��Ӿ��þ�7��HF>��o?;%�?vY?>TV����=!��=Y3?R�K?�qc?�_?��]?�{?=���>��>ng? �?�r=?dH?n�?v�s>cl>����>�輽�S��! :����f��X=�=$�v�Ȼ�<��ϼEr�=�Q6��ｽt�=���;���+���<d�q=�*�>d?̎�>�d>A*?mP.��y8��ⅾ<�C?5�[=M�f���n������ᾤ�>��k?�ȫ?rU?�f?>G@�A��n%>=�>��>>p�b>+�>��ѽ���W�K=��> >�*�=�bc��sw�%�
��}���z;zB>���>�/|>P����'>~|���/z��d>M�Q�x̺���S�V�G���1���v��Y�>�K?��?ƞ�=_龽+��!If�0)?
^<?�NM?��?��=��۾��9�M�J��?���>aZ�<��������#����:�Û�:~�s>2���8��z�_>q�����m��1I�yP�iT=-����2=���u�Ѿw"�����= �>1����!�h���J?x�=h�����e��j��vs>a|�>�+�>�EJ�u��ȳ?�k���i�=E��>�6A>Br��n[��I����,�y>�7;?��b?�#�?8خ�XQf��R�����I��Fѽ�<?��>�-?z+�>��t>�/i��� �[h��b����>��>�m&�$�a�/ľ��P�7�F��>�?3���>C�I?*�?d�B?2?��?뿍>s��:\�k�1?}��?���=p>�����:b��Od�mC?�^?���h�>��?Z6?�'?^�h?��)?��>�9��_��q�>�
�>��T�����#>2�0?���>@f?���?Ƅ�>,�@��G��������]�6�=s4?=G:?��3?`��>,?Q0��-��>��>Q2?o~?u��?t�>�m->��>�;?l�=�O�>ls"?<\D?@CM?�e?�?x�>
�Z��6ݽ�c�����׫C�h�=9?>�af>f�0>U�%>LZ�4ˡ=��=MR��1�0��ES��!,���4,��_�>��s>�����0>��ľ%K����@>�j��P���؊���:�Nܷ=r��>��?謕>S#����=��>�I�>����4(?��?�?%> ;��b���ھ��K�U�>�	B?V��=�l�0�����u���g=��m?�^?�W��&��I�b?��]?"h��=���þ��b�܉�T�O?3�
?]�G���>��~?e�q?I��>R�e�4:n�(��Db��j�2Ѷ=cr�>LX�K�d��?�>_�7?�N�>)�b>J%�=Ru۾�w��q��c?��?�?���?+*>��n�U4�P�����2U?���>=ڝ�Z�0?��!�	�ྡi��Do�+b辮9��+��mb�2��1�3���_��櫽�">{I?��j?�g�?�X?�A�3�e��^b�����7k�w��c���[/�?�1���L��j��I#�S��(Q�����;�~�ګA��u�?]�'?��/��.�>Θ�Y��̾�dC>�������9��=�s��p�>=�Y=��g�.��í�7 ?m�>g��>M�<?G�[��:>���1���7��z��:u2>ƚ�>���>zF�>?0:8�-��d�~!ʾs���!Խ�d>Ko?yiR?jh?W���kC�i����=����/;'��=nC�=��>%�G�DY<�~Y3��6E����8e��g��[
�ڨA>Z�3?�o�=,�>�<�?>�?�����(l�[�h=��-�渄�x6�>�?{)?q�z>*�f��J��ܷ�>��l?��>L�>%����Y!���{���ʽl$�>?߭>��>��o>`�,��#\��j��M���d9��v�=y�h? �����`��>NR?a�:�G<�{�>ͨv�`�!�����'���>�|?癪=��;>�~ž�$���{�17����,?��?�{���.��C=>�:?���>���>O��?*c�>������=*?snX?�%G?vF?_��>rCt=����̽��%��x=�:�>�m�>�)�=��>�mཌq����%��=&ӵ=��a1ýȼ���h�E�:7t<C?Z>�Dѿ7X�Az�1��,�������L��v(�9�P�`s��ҩ��'�i�m�r��6	2�L����7t�ˌ��R���s�?&�?�|��ž���yJ������>I�.�e�½��+��������Ⱦd�����#�=�C��K�BNe�p�?�R�9ӿC~��g�f=���>aQ?h?N?�����$�W�L��>���,C���۾BF��C⿻԰�C�f?7��>w�����^����>��>�@�=�t¼Ծ��H�zcd>&�>��H?�	?0ܾAuҿ	鳿EÞ==��?�@�|A?4�(����g(V=���>I�	?��?>�P1��K�����W�>V;�?���?1�M=Y�W���	���e?��<��F���ݻ��=K�=�.=���ؔJ>�W�>�|��UA�z@ܽ��4>�օ>͖"���&�^�R��<��]>J�ս�6��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=�� ��<ǿ��$�����Y<d��;����ֽ ���sF��#Ւ��N��>нS�N=���=��g>�w>l�:>k�H>U�Z?��k?p��>vP>|��Euξ�6����l�i{�������߽Qc���徆�վ[L�@s�	��ҳž�7��p	=�{`�����5�$�8�]��z4���$?x4.>��޾�\U��n�= ɾ�w����<rh���߾�1��rw�e;�?ϴV?�Ѐ�;:x�Ի�&fN=7ཪX>?�(���?[Ǿ8��<��#�%��:���>��B=�0�?xL��sP�?{4?b"0?aN������8�=OR&��d;��A?��?³�<�I�>]�'?�%������|~>�f>/��>Z��>���=j���-۽��?�g?������t�*��>�վ2�ھ=�>�N$� #9=U>2�k=\a��e��=�����=�(W?���>Q�)���c��k/��$==K�x?�?�,�>Syk?��B?��<!`��j�S�����w=K�W?�"i?ϲ>7�����Ͼdj��b�5?T�e?��N>Chh�����.�Q�"?k�n?�[?�3��u}����W���q6?��~?�]��<��ж�<ჾ��>"��>:F�>��&�Α�>��!?��Ծ�ܡ�s�ȿ�;��`�? �@a@��>�$�����=��.?Y��>K9����x��T�)4ƽ�?�tƾ�G����Z����-�?�^�?�?����A�.�:��=VS��R�?ǲh?�܏��(�=�V&��2��n^'�:���C=91����伱$徴�I����b��x��k�H<�G�>�r@m�=��?\ 
����yο�y���_�$-?���>�t�=�d�'ċ�$���!h�0�P�jo���M�>��>����:���J�{��q;��&����>c�k	�>L�S�-&��q�����5<�>��>��>Z,��R轾3ř?�b���?οs���͝��X?h�?�n�?q?��9< �v�^�{����-G?��s?MZ?�p%�#>]���7�h�j?S`���U`�u�4��GE��U>�"3?�@�>��-� �|=p>݆�>�a>�$/�0�Ŀ�ض��������?݉�?$o�}��>���?�s+?�k�8��XZ����*�S�/�=A?�2>�����!��0=�7Ӓ�{�
?)0?&z��/�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\� N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>eH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?x$�>�?�s�=yb�>�`�=P�u-�Sk#>u!�=m�>��?)�M?GL�>�Y�=~�8��/��ZF��GR�5$���C���>G�a?�L?Lb>[��2��!�?}ͽd1��>�DW@���,�m�߽�)5>~�=>>U�D�Ӿ=�*?8���߿�����o>	�>��$>Z-�>����P�uY��q?,W>�?�*Ǥ�yK����q�4��?`�@�.?#��<��=���>�:	>t�=@�<�f)�s�׽��m>�N?�9Ⱦ4��i�q���>M��?�{
@��?�K��+?L<��o���t�B�Ӿ��a�6�
>&�#?(�Ǿ�1�>�%�>Ӕh=~�u����k����>���?�H�?��?m�c?��g�1r��G>+@>aT?}�?s?��AA��/>G<?C�B�*��S�Q�M?V�
@y�@lh?�:��D�տj���̧���-���>$4O=!��>��=�.�=R,:�I8/�	>���>X#�>~�> �2>cA0>L��=Q��=�������U���HL�����܈���5<��ھMG��Q��:֛�c�����͠h��ɽ+&�
�I�4��E:�=��R?%Y?�w?���>`_��ΰ�=^}��F�J<o�-�T��=��Q>�=.?�G?'?�q�=�ݯ�y�j�]��o����
��b��>��{>��>���>�>��.=Y�B>��[>��>��&>'�=��=+��=}qk>��>J��>�¬>�� >��$>a���P޿��RI�]b��p���Ք?�q���zZ��䔿v�k�8��$=n{6?&|>�H���Uпu!��4P?(?���#�Lk��|:�>3~#?��Z?��>�S����p���>܏2��ӌ���=��ѽ���Q�E�B>�,,?�f>�u>֛3�e8�v�P�}|��j|>�36?h鶾=D9���u���H��cݾJHM>�ľ>�D�l�~�����vi�;�{=\x:?ل?�6���ⰾb�u��C���PR>w:\>U=Li�=�XM>ibc���ƽXH�g.=��=�^>O?�+>�V�=�0�>�0��N��a�>C�C>�d,>8	@?�|%?����)H���H,��w>��>3߀>i�>��I���=5U�>��_>���ł�{��U�=���V>�x�~�_� �v� v=����=��=���=����x�=�Y� =�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�h�>�x��Z�����;�u���#=@��>8H?CV��K�O��>��w
?r?�_�թ����ȿ�|v����>��?l��?F�m�7A��_@����>|��?�eY?�ki>�e۾�[Z�ъ�>��@?5	R? �>�9�m�'�1�?M߶?m��?V�]>9{�?�8o?\��>^��<a>���ǿ�d��r�
��ו�$��=�C>�eӽ|�/�2ǰ�`���Y�u�!
9�ɬf=#�[=��> ��/Zs�;p=E1d�(�q)Z����>�e�>�t<�V�>SU�>v�>Ӗ�>�m>>�����e���?¾�K?0��?i���;n��w�<�ӛ=��^��7?��4?�vW�ìϾ8�>֭\?���?�[?���>����*���࿿�s����<��K>��>�S�>�:��%K>4�Ծ��C�B��>���>J,���rھx)��5t���)�>�m!?L��>�4�=ԙ ?��#?��j>�(�>8aE��9��f�E����>���>�H?�~?��?�Թ��Z3�����桿��[�A;N>��x?V?�ʕ>W���䃝��kE�wCI�����\��?�tg?�S�$?:2�?�??Z�A?)f>��ؾ����>s�!?�l��jA���%�9�(�?��?R�>����ӽ�Ǽ����d��k,?m(\?�7&?�L�\�`�n�¾���<����U�LU�;2�K���>�o>C��@�=�>��=wEm��O6�;Te<з�=�>҂�="�7�(落�2?O��n����P�=�����i�N��>2����о�B�?\8޾99��˙ȿn��G���u��?���?���?|���Q�u���^?U��?���>�"�>�a�r@Ⱦ����ہ��Uݽ'�C�~��=k�>J��=����ԭ�CS��&����;��A� �?�
�>���>nZ�>K<�>М�>`P̾��,�A@���ɾ]zr� z8��T�R<�&��	�>��zK=� 	=��ƾ����>*˖<$\�>y�?#4>/[>�6�> ���!��>;��>���>�O�>��>�т>��=TS��7|�uKR?������'�������x4B?�rd?2�>�i�"������?���?qs�?B@v>�}h�,+��m?/>�>��p
?D:=���G�<lW��Z��A��%#�8��>�=׽�:��M��gf�2j
?�-?/1��u�̾;׽�B��&;r=J�?��(?�)���Q�G�o�0�W��PS�V����g�����=|$�ҙp�1������6��ޚ(���*=�n*?-�?B�v��)ꬾd_k��O?�.�f>�I�>�s�>@��>uQJ>�Q	���1��X^�	U'������]�>b�z?�®>�R?�*G?�(S?��$?���>�>�ky���@>a���B�>���>6K<?k�??0Y=?J%?'�(?e�I>�۽��پ�����.?
?�k?��?Q9?H����ԾI�P�/S=OZ��я��՝
>c»��	�j=�n�=�>�X?̙�v�8������k>��7?���>���>���-����<}�>�
?}G�>�  ��}r��b�nV�>���?���ς=5�)>#��=�����Ӻ0Y�=�����=�9���x;��e<{��=���=�@t����b7�:���;k�<�s�>U�?[��>�B�>x?��� ���[_�=�Y>+S>1>Hپ'~���$����g��[y>�w�?�z�?��f=��=���=�z��(T��#���������<|�?�I#?�VT?�?��=?�j#?�>�)��L��{^�����d�?w!,?��>�����ʾ��։3�۝?i[?�<a����;)�ߐ¾��Խб>�[/�i/~����>D��텻���W��6��?�?IA�W�6��x�ۿ���[��{�C?"�>Y�>��>U�)�~�g�s%��1;>���>lR?r��>��O?�D{?"\?]�S>s8����j���*s9��c!>hX@?ݒ�?t�?��x?6s�>I>̌*��������o��W��T(��o�V=�Y>�>���>P�>F��=��Ƚ�
����:�x�=%'c>���>�ѥ>�K�>��w>0��<BMK?�	?�Z��9��F�־%������{?pH�?�J+?o�/=�c�z.�.aҾ'�>���?�ת?2#?7����=W��.����C��]�>���>�!�>���=5Q�=�NA>2�>���>�{���
�N&;�����e?�q@?�]>��ʿ��{��f��d��2eF=�~�2E�ߧ�u�H��"�=��p��������G�*��;�l/��~��������>�(=��=]ߔ=��C=��<�s�;G�Y<Ļ�<LЅ=��(�IS�<9	e���E< ����=�;�<#��<4�<�!y˾7�}??DI?��+?�C?m�y>Q>2�3����>�����D?
�U>TP�Cg��oS;�����Z8����ؾ�׾�c��ӟ��L>�H���>Y3>n�=�܉<��=��s=�~�=�gF���=���=���=���=��=��>P>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>I�7>D&>��R�ڈ1���\�;�b��{Z�O�!?5I;��G̾�9�>���=�.߾�ƾ�m.=�6>�pb=�]��S\����=V{��;=�l=jՉ>��C>zu�=�,����==�I=I��=R�O>�4��Jn7�9,�8�3=���=�b>�&>��>�.?�g0?�d? ��>��i�"�˾X���׾�>�o�=4�>�P�=m�B>��>�8?�D?%rK?���>�%�=i��>&]�>l+���m��G�X0��f��<ˈ?`�?�˹>Z/O<�XC����(�=���½�3?6�1?�?�9�>�_��P�K/�Œ��F=�ڔ>��t>qX>`�<2
;���;W�����=��>�B�>�O�>�W&>C��������>���=��B�����'����'�ս`<��啽�����$�=��=}�=���g�>���=Y��V��<靔<�t�=�Z?�=H��R�>Z�;=XӍ�4[J>+ƾQG��®>8�D����X��W�V�P��𚾲!�>��>{p�ё�$�?%�=>�H�=2��?�Β?�Ӽ<I[���4ɾ�5��e��=|�8�6d>2�G>L�M���3�=�O�Q�A�Mդ����>]�>J��>Q�l>�,��?���w=��b5���>�����P�C�R<q��@��m���Si���ȺZ�D?�E��B��=%"~?��I?��?5��>x4��J�ؾ�40>�R����=X�nq�qi��u�?]'?��>��D��H̾U���޷>�@I�-�O���U�0�X��+ͷ�9��>������оm$3��g��������B��Lr�c��>+�O?��?a:b��W��EUO����h(���q?�|g?/�>�J?�@?=&��z�r���v�=�n?ͳ�?U=�?l>��=�(Ͻȍ�>;�?k�?߬�?x�u?��,��n�>�@�<Eu]>����m3�=**(>�#�=�|�=��?�?m�?�����z���������������<�>�̩>4�>⸑>���=0c=>�\=�^>�2�>��>bڀ>�?�>�Dq>����>t�L�?�m=�h>UCP?ͺA>8��pC�W">d�*<����fQ��.0�L�S����;�U�=��#>3�=�k�>��ſ�ɗ?u��= 8����?aD���7��7�>	�A>35��m��>�8�>��?�Ӳ>���>���=B�=�\>�;Ӿ��>����s!�QC�	R�N�Ѿ�z>�����"&�}���q���VI��l���]�wj�f3��wA=��v�< G�?�����k�-�)��O��x�?
[�>�6?Hڌ�9݈�)�><��>ż�>uK������]ˍ�ip��?���?�;c>��>H�W?�?ג1�-3�vZ�,�u�n(A�+e�U�`��፿�����
����-�_?�x?2yA?�R�<+:z>Q��?��%�Zӏ��)�>�/�'';��?<=t+�> *��*�`��Ӿ��þ�7��HF>��o?;%�?vY?>TV����=!��=Y3?R�K?�qc?�_?��]?�{?=���>��>ng? �?�r=?dH?n�?v�s>cl>����>�輽�S��! :����f��X=�=$�v�Ȼ�<��ϼEr�=�Q6��ｽt�=���;���+���<d�q=�*�>d?̎�>�d>A*?mP.��y8��ⅾ<�C?5�[=M�f���n������ᾤ�>��k?�ȫ?rU?�f?>G@�A��n%>=�>��>>p�b>+�>��ѽ���W�K=��> >�*�=�bc��sw�%�
��}���z;zB>���>�/|>P����'>~|���/z��d>M�Q�x̺���S�V�G���1���v��Y�>�K?��?ƞ�=_龽+��!If�0)?
^<?�NM?��?��=��۾��9�M�J��?���>aZ�<��������#����:�Û�:~�s>2���`��4�y>E�������S�`P�-��}E>"�!�sj�<ap!��.��鵈�	u=��=�¾^�������ܳ��GK?��=�h��/��0s׾kC�=��>)7�>��U����n=�dγ��H�=��>�A>��������Q����Ո>]�8?(�L?�"�?~��W��y�Q���j�����>/��>�w>��N?�>ޔ�=J���{0���p��ha�BP�>qk?�.)��p�􇩾����d4�^�	>l25?"�,>䩃>�_?��>��D?dL<?���>Ą>ر�1렾$�%?���?U{=
�.��-��5/3���c�9��>�C?Z0���=Iy�>�\P??^8?��c?��?�o#<{K2�3�V����>cf�>��6�*#���L>	[?�"�>�K?P��?�&>B�<����������>0�>��?z
?)E�>�>��>�~ξ�Z����>�a?�|?�Ј?�D�=��?ŹV��S*?�>A�<ś??��.?�E?P�S?+�!?��>��==�2N�D��W壽�F���<X��=��e>Gã�Ψ��}��rˋ�P��s�M�3U=�X�	@���a�+:��u_�>��s>�
����0>0�ľ�N��w�@>����4O��8ڊ�M�:�C�=���>�?Z��>W#�K��=N��><I�>���6(?��?�?�l!;	�b�Q�ھ��K���>p	B?m��=��l����� �u�eh=��m?�^?k�W�G%��3�b?�(^?G�򾊗<��{ľ<�d��@���N?�(?��D��H�>�\~?�r?���>VSb�*vm�(✿��b���n��'�=��>�,�E�e�Ԗ�> �7?e��>n�b>Ϯ�=	"۾l'x� ���=�?��?-f�?ˣ�?��)>��n��q߿���U*����i?��>�_����$?ۓE�N��z��	�y��Ҿ5��Ǎ��A���=���d��j���ݽG)�=:6?1)q?�oi?5�c?�� 2h���]�^��bP���I��JD�t�8��=E���n�7������˲�2d=t
h��M�ܗ�?1�$?S:ܽo��>����n;qUܾdkd>�j���ֽo �=L���m=��y=KX?���'�߀��t=?&E�>=��>l�D?�i���C�<�2��HD�w.�->�I�>t{�>�a�>[��;j+�%�3�ھ�ͣ�~�۽f�>��Z?q�[?V �?<f��
�A�����D7������辆au>���=���>��n�.�}�s��\h�2ǒ��s�?ʞ��(���{�_7?HH�>��>���?[I?=�%��l�R��Wa��>lf�>���?�e�>��>|f���yJ����>$m?E��>X�>񍍾Ç!�s�}��Xཛ��>���>���>%s>Z�*�n�[�0���H��>�9�>��=�g?.˃� Fb��̅>+bR?i�ݺW9<�]�>�ec��!�z����9+���>�i?8S�==F?>�o��gR�8|�%����[!?W.?_�r��6B�AA>��;?1c�>S'7>�i�?SR?�~h��ط���?��J?��S?7N?���>�m�NT>���
�5��Y >{��>(��>���<�K>+re�:͑�����>p�>,S!<�< (��G����>:s�=��?>�ӿ9�U��/���e6��K��)M����N�=a�V�@eD�7�پ$傾0��@�ý�J�<.-�r�o����T��?E�?=���&�@���t�C4�v?�,��l��=8���L���YD��Q���;?�#��U=�!F�SDY�T,?T��9¿���v�ן�>W�?G�?r�)���)�FC�|yl>bw�	lB���ϾwԬ�|�ۿ�?���Nf?��?����4�Jx�>��>j�k>t�R>�dʽ6� ���=|?eh\?��?NJL�\`ſ��ѿ������?9�@ }A?%�(�q���V=d��>'�	?3�?>8S1��I������T�>b<�?���?F{M=d�W��	��e?j~<��F��ݻ��=�;�=NH=i��J�J>TU�>b���SA��?ܽ��4>څ>�}"������^�E��<�]>T�ս>;��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=u6�����{���&V�}��=[��>c�>,������O��I��U��=-��cUſ�#��1!�=��<��Լp\d��c���?���0�ɷ����n�O1�잛=N>��r>�E�>��&>yB>�H]?t?Xơ>�k��JY�SQ���uƾ���=ST���4�������N���kv����7�3��H	����e¾(�&�xt�=�<]�SY��_�񾚂^�Z�<��BX?�����ݾR)i���=Mݾ����Ɠf��Խ���&��w�S�?�Z?�`����H�& ��[�b�Ƚ��^?�݂����j������=R��;�Nɽ�B>*@�d�/c?��v��{a0?�?�<��̸��i�)>V}��`�=�s+?��?Zox<�m�>?#%?M*�&�⽓\>�W4>�*�>r�>�J>w/��x�۽��?��T?��(�����>�I����z�.�[=��>fd4�`��?a\>�?�<K���zV��Í���<i'W?4��>z�)���9]�����=k==v�x?�?J)�>Z{k?��B?���<�g��?�S�< �zzw=��W?�(i?��>�����о0���=�5?�e?�N>"_h�1���.�S�P%?+�n?�`?e���v}������tm6?20?�qQ�K盿����[���qZ>3�>���>R�D�r�>a�?J!�xa���T���uC�|��?�C@���?:�F=��½�:�=�L?� �>Yo~���$���$e����`�	/	?t���#���I�L�7�SE-?)�l?ҁ?���Ѧ�E�#>�����۱?�9�?0��DG;�m�f�Y�L����<����#H=�=�<�]���A���ݾ�$��Ѿf�c=��~>v<@�|��a��>CyǾJ��,K��L����a�3���{>�d�>�ҽ��ھ�.��SX���{`�s�H��c��IN�>��>	���������{�r;�i[����>! �'�>�S��%��^���4�5<��>��>��>D9��d꽾�ę?�_��e?ο꫞�����X?g�?En�?s?�w9<o�v��{���O0G?F�s?�Z?�n%�aA]���7�Z �?�9��7u��=%��O���>ie*?	�>۬?��>�k��II?5�D�;,V�b�ſ陿y7;��?w��?jU辴"?�¨?��'?k�6��G��3C��h,�����G�?�Z>��ރ���/������e(?&`�?��<�p�<�]�_?*�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?ֵ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>cH_���u>����:�i	>���?�~�?Qj?���� ����U>
�}?W$�>��?�o�=�a�>�c�=+񰾦-�5k#>�"�=)�>��?m�M?7L�>�W�=.�8�`/�[F��GR�r$�3�C���>��a?��L?�Kb>����2��!��uͽ�c1��N鼑W@���,���߽(5>��=>�>��D��Ӿ��G?G��޿�׌�/_S���'?뵏>h&?9�!�6�ʼ�O����~?0��>�!��z��~Ø��ʳ��ս?R��?�I?�7پ e�<��=�`�>�i}>�Q��0쪾aH���">�I$?���+��/����&X>�|�?@��?I��?B�b��	?���P��y`~���7����=��7?2���z>���>�=pv������s����>�B�?�{�?���>��l?�o���B�O�1=|I�>��k?.s?�wo�t�e�B>5�?�������K��f?��
@�u@Ŝ^?}<Uڿ���������W����>�׾=�_D>����<+�,<�$p=h���Z�=b��>��N>EJ{>S�>/�G>u�#>�h��z�!��Л�fK��=�$�,�������N���8��=��}�2=������j3�F�S��;L��q���k�Ty�;��=O�G?e/R?Q�?5��>�;�>�=�+㾗���N<ڽx��=h �=�GO??B?�B?A�h=�����dn�����q��B�>4�=)�>�(�>r�>���;@�P>u��>�1\>B��=���='�<?y1=�.!>�׷>�>��>��G><F0>Y\��m���R6e��ێ�W˽S��?���o�J������>��E�ƾ�)�<�'?S�=�t�� eͿ<﮿1C?�����"��f齖�j=��(?IU?�c�=Q���(~��?�'>�����{�8=�=����������1���F>�$?_v�>��>�-K���0��ZG��#��1N>tI?<Ӿ�]��+��;�1��;����J=H_�>���\&������T��P:Q����= oH?��?ư��,���K�D�ھCB�>۫�=ђ=��*;0��=ѕ�fb���]u��/ͽ��=��>�U?"�+>���=ϣ>�W��8P�/��>�^B>9,>�@?D.%?�u�p���n����-�?3w>�[�>b�><>ZJ�ǯ=�i�>��a>�	��񃽚����?��cW>�k~�Ib_�x9u��x=����=:�=�� ���<�~�%=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�)?#�н����j��av��=���m�>��y?��6�=e:�qZ��&�Y?�\�>�Q�Is���>���% ?� �?$�?�@��7|���^2�@�?Ö�?#�B?��>5�����=9��=��:?�܆?���>�Y�ѵ�t5?w(�?nz?W��>�\�?�F�?�y�>�o��(�(tͿϬ��ޤ=�
.=y��>���>O�G���`�x���擿�!p���#��ٲ>T�2=�;>N���a���f= }M���о,�S����>���=��>��C>k��>M�?2��>^�g>�1�y���������??���?��Ѿ�q���t�p�X>�Z�
U�>�#k?<��>�þ�j�&�k?�ބ?���?�E�>ɒ�J����������J=%>	$�>��>վ[>_��>⥿�'���j��>C+?���!����n��׽��>�5?��?�3�=�� ?�#?�j>�)�>aE��9����E�Y��>Q��>�H?W�~?��?�ӹ�v[3�	��#硿��[��7N>��x?�U?�̕>���������KE�>I����"��?�tg?�P��?+2�?~�??��A?&f>���xؾ������>e�!?���p�A�jH&����C�?�>?���>���{�ԽK�ҼX���V��Q?_4\?�F&?�|�a�þA�<i�#�bU��I�;�A�:�>��>�W���ǳ=y�>T��=
m�+r6���b<��=��>��=f�6��@��$�;?l�;��}��*�;���5�n�bYw>�W9>�<
��ju?h�����n�������Ӿ��G�q?w��?~�?]mνܽ|�H�4?�?u-�>Kg?�}����������:�h��q���$��4g�ض�> �����׾����������[C3��R����>6�>;`�>��?X��>�p�>�Ȅ��~&����e꿾.~�Y�� �-��QS�E7"�+�$�I��j`�˾֓z�{S�>��%����>�J?���>�f�>׆>O�=ٴ>Bm�>��>���>dT>i�=�CI>��==7���KR?�����'�h�辖���h3B?�qd?51�>�i�4��������?���?Rs�?;=v>�~h��,+��n?�>�>$��<q
?yR:=o7�9�<1V������3����V��>�D׽� :��M�1nf�{j
?�/?�����̾);׽*����5�=��?�`/?,)���T��X~�r]\�"�L��8üP�����l�X���y�Ԧ���������^,��$�=K�?8/�?ǳ�a�쾭��_?c��b�$��=ȅ ?x��>���>9"�>T���X�+�t�f�.F3�������>�v?xD}>ݻb?x�H?\*?Ca=?���>~G�>t����?���>�?�L�>��3?(�:?uH7?4�+?�$#?	�j>ፆ�PN��i�߾��9?�bh?&�$?�q�>8�?�����Xd���V����=�Je��Ƚ�(>D���F1�--��� >�41>�X?���Ϭ8�5���yk>W�7?���>��>���-��?&�<q�>;�
?�G�>Y  ��|r�Jb�\V�>)��?b �k�=v�)>B��=j�����Һ�[�=4���4�=�M���|;�_P<��=|��=�!t�|с�S�:
Ї;�i�<�t�>6�?���>�C�>�@��(� �]��f�=�Y>S>�>Fپ�}���$��{�g��]y>�w�?�z�?ϻf=��=��=�|���U�����)������<�?8J#?)XT?`��?|�=?cj#?�>	+�iM���^�������?[,?ߑ>�I���ʾ�Ө�T�3��V?&�?"a�PH��)��[¾�Rؽ��>��.���}�G񯿂ND����&��������?��?�)O�]6��^�=���� ����B?JW�>���>���>�m)�؈g� @�tw8>�a�>��R?�׻>��O?�#{?�:\?dR>2-9�����q��o6=���">N�??�?�1�?�8x?L�>�A>�=-����8����0�`������RP=Z>�[�>���>���>��=#5������K->���=-�b>�S�>�*�>j��>,x>B�<�G?ұ�>ރ���� ��<����G�a<t?���?�,?��=����lD�W ��fx�>�5�?�Y�?��(?��W�mw�=?�ܼ�ϵ���o�m�>�Ժ>�-�>뮈=�.=�> >��>F�>>��l���8�C;�;?�jE?��=`�̿��o�����Hs��J���A־C�Y��<��LN�^G{>�d��Y1��6��<�i�i_i�r>/�����1Gx�3t���g�>��=n�@>5N;>'f������.����W<���<���=������=Ë�~�K���j�<�o4<°>>z.�=4{˾߅}?�<I?��+?�C?
ky>�>=�3����>�6��@??��U>7	O�r���r;�ʡ���*��`�ؾ�׾��c�$ß��&>��I���>�(3>�=v��<�0�=t=S��=��L��m=-��= N�=EG�=�=t�>�T>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>5�7>}.>��R�i�1�S�\�&�b��yZ��!?Q;��F̾k�>��=�/߾��ƾt�.=Vt6>��a=&��Bg\���=�z���;=xDm=Q��>�C>:��=�y���?�=�/I=��=b�O>�v���8���+���3=ǎ�=�}b>� &>G��>��?�a0?�Yd?�9�>�
n�dϾF=���K�>�=:I�>
օ=�yB>l��>��7?�D?��K?���>���=0�>!�>�,��m�}m徵ǧ����<1��?�͆?�и>W2Q<��A�v��:d>��"Ž�u?~P1?�j?�>���ӿb���k�Y�N��w����a�v�j��=P��[@�V��(yf�<:�>���>���>��P>��z>ܐ>�M�>Hܝ=)�}�ʥL=��W=�2S��y��li5>�<ȑ��_�0���>=���Fٽ3�n=ap�<q`!<���D��|*>�.�>13�=6��>�K�=����>f�T�;U�6\�Eɸ�U�b�O������a_�B�j��
�>��>�_������k�>S�=)k>[1�?���?nއ>� �TҮ���rN>Ǯ��>D�>��3Q,�Kk��M��������> ��>��>�l>%	,� "?�^�w=g�*b5�c�>�z����'6�m:q� A��.���i��4к��D?�F�����=�~?x�I?b�?5��>����҄ؾ�@0>4M���4=���q��8��f�?�'?���>���D��H̾R���޷> BI�`�O���>�0�����̷�Z��>������о^$3��g������̍B��Lr�.��>�O?��?�9b��W��FUO�����(���q?�|g?�>K?�@?�%�� z��r��nv�=��n?���?J=�?�>(۵=�㱽L6�>�+?�z�?x��?ϻt?X@9����>�/���5>�@��>C�=$�,>�=��>Q?�?"�?o�����
��z������h�d�1=�j�=��>Oh�>��t>;r�=^\=�h=/nf>)؞>p��>X�W>z(�>�"�>�a����5;4?��<dK ?�ya?ٮ�>�P�>������=p�s=�VϽ���P2(��(��m~���N>�~>���=��>Igٿ��?{�>�ؾ܄�>������=]/�=AC�>0f)��,?���>���=ѽ4?Z	�>w7���7=Y��>�U���2J>������VQ�2�U�S�� ��>+ڪ�IKi�S����^f����Ͼ����,l�z����W?��g�;Y�?�r��]�V��`��,����> �>�2?(���sK�ؓi>�N?��u>+������u��h����?���?�;c>��>I�W?�?ْ1�33�vZ�,�u�n(A�-e�V�`��፿�����
����.�_?�x?2yA?�R�<-:z>R��?��%�[ӏ��)�>�/�'';��?<=u+�>*��/�`���Ӿ��þ�7��HF>��o?<%�?wY?@TV��6K��J>��G?��Q?ӈ�?�P?i�g?#�����5?o�W��n;?�J�>�?	hY?��?���>��>Ej>iA���wK�	���<�G��Aӽn��;LL�<�:�9�Z2�L����G�����q��=���;�e{��/��E���>4��=��>�Ʀ>�]?.�>&F�>vh7?�;��98��7��Y:/?�J=������gġ����>k?��?�Y?Lb>.�B�fNC��>�h�>4s'>?�Z>5��>�:�$F����=N�>��>���=��E����u�	�: ���\�<�'>��>�3|>���ó'>�|��K-z�=�d>)�Q��ʺ���S���G�B�1��v��Y�>��K?��?���=l_�D2��If��/)?�]<?�NM?~�?c�=t�۾��9��J��<���>;p�<��������#���:�$��:��s>�0��<���4jY>?�3�sKھ֟}��Q���� �=���������*��뚾�}�=ue:><о��E�KL������VR?�$=�W���P(�@>�.=�;�>c��>�@��θ��@��ѥ�_�<	:�>�cs>A���j����JZ�
��w~V>
01?��]?�Ƙ?���vy���7�k�־���p+<;�@?��}>Y�??�pO>r�H=9�ɾ�i2���T��6'�d��>���>}a
��c�T����\���p<���>B?(?n�{>���>ǔ�?ʾ?
�g?/7-?�X�>��>�����De'?!y?c��=q�)��bD�S���xU���>��1?wh��^<�>��6?w�A?p�e?v�b?o?�U���M%��N=��>��~>f}K�ae��7�>�P?Ӱ>S�e?�σ?N�&���C�U+��F��R>�(f>�',?*E?�B�>���>f��>̄��G4�=���>8c?�5�?�o?H"�=�?2>`��>�Q�=���>]��>Q?_RO? �s?I�J?o��>_J�<�~���<���r���O����;J<Iy=7�St�����x�<v�;���<��U��
�D�������;d_�>9�s>�	��a�0>��ľ�O���@>���P���ڊ��:�Oܷ=���>��?��>'Y#����=M��>�H�>���6(?��?�?�";ߡb���ھ��K�Y�>T	B?���=��l�$���Q�u�M�g=^�m?~�^?��W�>&��?b?|�]?;��+Y;�>�ľG�d����M?{�
?YF���>�S�?Cs??�?)�Z�hVl��e��c�C`n��!�=jl�>YT�"h�߇�>��8?���>�zh>�"�=��0Hv��,��?�?jߍ?���?���?[�(>An���޿��������e?�7�>5����#?��)<#Y̾�㕾Tq���hܾ�Z��&������,��r|$���w����Ϟ=Kn?�u?�[j?�f?!	��&c�~3_��~��PJ�D'��g�r9@��B�^a;���p��x�F��2ȝ��t�=0�����S�Jk�?�'?���,&�>yh��'Ҿ�澔#>Pۚ������=�h��7���(=W�1��;��繾22?YV�>Ee�>�zH?��f��g4��G1��ze��kԾ��+>N�>�Ɉ>��>���;+l�N���ȵ��*u��T�!>�Y?E�H?�s�?z�"����y��,%���=�w䛾���>	�>(��>�^n���O�q/�}JS���[��.������ь
�*y8�\J>?�>ê�>�6�?�U?RI�7?"�١�=��U�i�\>R��>V%Q?���>�=�������>1�l?6@�>.�>U��U;!��/|�'VϽm6�>�7�>(c�>S�p>�B+�l�[�]7���_���09����=@�g?�O��Ima�u��>��Q?���8��W<w9�>n��\"����xb#���>��?��=��=>�ž6���z�M뉾�I#?I�(?2v�!%�?]�>ܡ,?�^�>\c�>���?K*�> -־��=�0?��S?!D?:11?z��>�m�<Zu��
��y�y��<ݕ�>�Oo>���=R�:>�ӛ�p5�+%��=Ȗ>�r=�U���׽˛<�S>�*>���=�ؿ��1��)��8��?ؾ~Tپc���ͻ.���V�g����"�nCv��i+�ł2�q=1�,rt�8t3�%I�s��?���?�� �3�������E�����>�F��&�D�������?ܾ��о%vZ�����A9�˘\���p�A�%?(�����ƿʞ���S���?A}'?v#v?�3��,�/�8�V�)>�z<�A9�/
׾R읿��˿�+����g?z7�>1w��|!��=�>���>I_r>s9>��j�@˟��X�=�H?�%??�O���@ǿ�i���KR=MM�?�	@}A?�(���쾄V=E��>*�	? �?>�S1��I������T�>p<�?��?�{M=�W�O�	�/�e?7<��F�p�ݻ�=�;�=4F=���ҔJ>~U�>G���SA�I?ܽ[�4>Qڅ>[~"�f�� �^���<��]>.�ս;��_#�?�+a�na�z�F�g2��#�"= g?o��>j<�=$,&?�w�J޿�u���N?�:�?���?@�>?_M�E��>�^���P?L7;?r�?>�Q+�x���mB>��м�Շ���jH�֍���C�>��,>r�u�e-��0�ðB�^޸=;A�Q�¿��%��v1�竃=�>a�(}��$�ý*1�O���WE�|Mǽ��c=ʦ�=�T>�z>"_^>~#�>4�c?��v?�Gr> �=�(�eު�������6=y}�d׽���r��5���P��`������/Z$��_���ƾhY=����=�S������� ��lb�DD�Yg.?�">V�˾!M�P�k<��ʾ�Ȫ�<�l�"�����˾6X0���m���?ńA?���S�?���.��/���V?�[���� 묾sb�=B0�+c=c�>]͚=`���4�b�S��50?��?޾�䙑�W�+>����A�
=-b+?�w?��u<��>p"%?p5%�ὁ	\>�4>�o�>l�>[X>D����۽u ?8T?�+ ��D����>�4����z���b=�&
>�1���漜�Y>��<����<�m]���a�<�(W?s��>��)��{a��~��0Y==��x?��?$.�>o{k?��B?�դ<'h���S����aw=�W?4*i?��>����	о_���E�5?�e?��N>�bh���=�.�^U��$?�n?5_?`~��)w}����o���n6?�W�?��m��"��R2�(�P�'��>N_�>\��>��L�͓�>��*?� �4����dĿl�0��X�?M\@pa @���f��)�1=��>���>z	��򼾹��8������=_o�>Z1ƾ�z��")�}�ĻE?�ܐ?��?�6���<�に=�.��#��?���?�i�Q�Z�1�w�>��d�<Ik�=��k�j�� ��GH���ξ������h�5<�:|>�l@f$i�\?/#���A޿d[ӿM��$�t���
l!?lH�>��q��}��!�p��4q���Z�z 6�I���M�>��>����`���_�{��q;�v"����>���	�>-�S��&��隟�Ƒ5<��>��>F��>n+���罾;ř?�c���?οD�����R�X?2h�?�n�?q?#�9<��v�͐{���<.G?��s?IZ?�p%�S>]�_�7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�i	>���?�~�?Qj?���� ����U>
�}?-�>X�?u��=t}�>�I�=.ﰾ&�,��K#>?��=}�?��?�M?�R�>�Q�=�8�& /��`F�xER�� �y�C�r�>d�a?�L?pRb>�s����1��� �y�ͽ�F1���輢r@��+��q߽�5>p�=>�>��D�RӾAG(? 3(�*�ѿT{����i��I,?T�p>�?,.	�Q"ý�Y<�V? 5x>S+�L'���p��!�����?�_�?5?Т��XD����=�v�>��>3G��gh�G꫾��V>п9?���s)���u��}$>?�?�@���?Λv��k? ?��l���Mz��2�
|��Y�=4�>?����1�>IG�>���="�m��鵿��o�S�> �?(V�?�?*La?V�n�Ĳ=��p�=|��>ETX?$:�>�v�� f�V�>0��>�N��O��*�����M?V�@[�@ZJp?u2���<�Q#��?���!S��=>m�n>yY&>�#��J�=F��K�ռ��:���=��>�I>8O3>��@>��e>�Rw>�����$!��.���񒿢3�������sp���D�h3���%�n�پ!� ���	�n���ؽ.����/A�/¡��V�=ZS?2YQ?.�s?���>�����>�}��N�T<Qs0����=z>�*3?�7J?�J'?9/v=Z7���d���������A�>��J>���>}��>%R�>ލ�;/�9>�K>?�>t@�=y�=��Q;���<��O>f"�>Q^�>�U�>ڎ7>��>�����ͬ���p��]��������?')��7�H�e/��V���")���Ɛ=#�/?�5�=_���7Ͽq���(I?WG��ڍ�g����=@�*?<V?�$>r���)�����>�J�sTR���=G����T�)���E>+�!?�Wb>��r>F�7�5��*V��������>be4?xO���>�#Mv��D���߾��F>���>̑���������~��uW���Y=�;?�*?�Fӽ0᰾��g��x���@M>u%f>�=D�=9�U>J���伽c\_��5=F�=��}>�S?��+>b��=-�>_���@P�{�>�oB>�,>�@?U+%?���8���4���@�-��w>|B�>��>�P>[J�x�=�l�>G�a>��� �������?�o_W>��}��n_��ku��=y=�%�����=�-�=v� ���<���%=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�B�>�=��m��D���rU��X�.��0�>�0I?���+=b�A�ƪ?/q�>�
�ْ��ҿx�i��>���?���?�Pw�lł��lM��1?K)�?�t?�a�>ߡ�Ce>�?��>TV+?��K?�Z>>P�.��y�=�3?��?��?ݭ�=�ņ?�x?��>V~��\q&����t��!�>���>^3?>B��>6澺"6�@P���u���m��e�`�>+�=���>$нx����&=证�Jʾ���=���>Em>�����+�>��?�
�>�[�> 1L=�v�<����(߲�|RF?ǘ�?U"�2d�$D�=�%>4���+???9P?m����+�>�i?���?N�i?�R�>k
�����FΤ��L���Ȭ=�0&>qd�>���>��<�eb>mۮ�h���d�>gj�=�{��þtLϾ����qBu>��0?΃�>F��=�� ?�#?Ǜj>D,�>�_E��9����E����>���>�I?`�~?�?�ӹ�!Z3����x桿ג[�66N>�x?YU?�͕>'���`���MuE�x6I�������?5vg?A彖?�2�?s�??.�A?*&f>I��Hؾ����a�>��!?����VA�#P&��(��?�?n��>q���3ؽ�ݼ6V�O�����?�^\?�&?8���7a�u�¾D
�<6X��Z���;�<���>��>sކ���=]J>���=��n��p6��,B<^��=��>��=�x5�r�����,?�#��.��Ƀ<�y�z��P�t �>��l>��Ⱦ�^T?(����f������3���lS����?�+�?cx�?�3��n�MGC?���?��?�]?�����㾿�ؾ�̝�_��������">`�>ʎ�����ԧ�����N�����"�G�>�>d�>�d?�,?�NR>!��>ܨq��H/�� ��";){o�>�&�'�*}-�<� �f�c�A�[��Q.�9�ɾ�M���&�>/(���:�>���>�Q>Kx�>fl�>{t��pZ�>�H�>�h�>��>B�>��>���=�<��
��KR?����'����e���R3B?Zqd?�1�>�i�7��������?���?ls�?^>v>�~h��,+�
n?B>�>1��Tq
?T:=�:�_=�<�U����k1����e��>tH׽� :��M�(of�Ej
?u/?���+�̾D:׽k��j�r=�&�?��0?N���R��m�a1h��5C��t<���{#��ρ&�b{o�}��ry���タ5D#�/�=![ ?�~�?x��x]Ӿ����l9e�O`V��#>�?[��>�C�>v�q>����K"��^��O"��P��'��>��v?�q�>r�S?"�'?��1?.�K?x��>l��>u���{�?��=�>=�?�N?�#?,�%?�l?R�(?���>M!��B���ľ�??h ?�?HX�>,�?OlѾ��3�����0>a��w��]�>_E�<�罔x�~Ϙ=?�`>�X?j��۫8������k>|�7?}�>��>���-�����<��>ڶ
?I�>�����|r��b�<T�>��?y��=��)>���=������Ѻ�]�=&���-�=P���;�(;<���=�=�(u�������:(�;�l�<�t�>6�?���>�C�>�@��/� �c���e�=�Y>?S>~>�Eپ�}���$��w�g��]y>�w�?�z�?ڻf=��=���=}���U�����H������<�?@J#?)XT?`��?{�=?^j#?е>+�jM���^�������? ,?y��>t�� �ʾ����U�3�W�?�X?�6a�%���@)�l�¾�+ս��>�K/�D.~���*D�鈻����������?���?�A�d�6�<g辕���IX����C?��>4Q�>� �>��)���g�!1�O;>\��>NR?ܻ>��O?^{?�M[?�S>��8��L���������Fa$>	�??���?���?κx?[U�>&�>��*�:���z��(�y��];����S=^�Y>#�>c�>�Ǫ>���=��νw����?����=Y�b>s��>kG�>}N�>Պv>'�<�G?���>�X��H���᤾X���hD=�.�u?]��?��+?��=0~���E�8:��
N�>l�?���?!/*?��S�M��=��ּ�߶���q�h&�>�׹>�7�>u~�=X�F=�r>��>8��>��yd��s8��/M�g�?^F?��=�\ƿ}�q���q����wXt<u��h1c�I�b[�<��=�ߘ�����r��8�Z�蕠������O�������y�o��>iL�=ԣ�=W*�=\�<m�ҼS(�<�PQ=�<ϛ=�r��Pu<>5��������	��6<�GI=t����ʾ�F{?jH?��.?��A?�ms>�p>�9G�v��>�?���?��E>5�o_��	 =�3����=ھYJ׾{c�K���>�7�OP>F�!>c#�=���<�p�=si�=���=�3���_=m_�=I��=O_�=���=��>yB>���?�!��ޝ��L��~�-?8m�>�aB>3���1B?�E�����`j�����?�z?: @5��?:�D?�i���w>�Q7���<~�Z��LD�é	>���>�(���?iz�=z�'��	���NK��+�?u2@Gm]?�����ҿ��>,>0�>(�R�^]-��-C�@\��L��z!?X�;�־�P�>/+�=��A����=	f;>a0�='��F�^��C�=Ya��a�X=�\l=�p�>��>>i*�=�|����=��M="X�=�uZ>��;�JF�)<�y%=��=�c>T�>���>��?ma0?�Wd?B6�>n��Ͼ�=���J�>��=IE�>,�=uB>b��>��7?R�D?��K?Ä�>g��=��>��> �,���m��l徝˧�嘬<q��?wΆ?�Ҹ>��Q<L�A�����g>��0Ž�v?pS1?�k?��>�!��߿�(%�5�3��i�)�=d|]=Z�i���p�?$���1#�liν�D�=��>d��>�X�>�z>x�;>te>.2�>4|->���AcC=|���4�<�@��oH�=$��^	=v�ia�;�+<l��U��4<���b�</{<TN�=p��>
l�=>D�>7O�=MSž"7x>%�i���S�/;ಾ�s^���r�9�\�_#�Խ;�>"$>������ ?�>d'�>h4�?{׃?�t�=����վ�J��Ğ�<�0���=
�$>�m��3x=���\���S��~�����>Eߎ>f�>{�l>�,�+#?���w=�⾛b5�G�>r{������'�l9q��?�������i�8�Һ��D?lF����=:"~?װI?=�?\��>���'�ؾR90>�G��Q�=���'q�Hg����?�'?���>��l�D��=̾z+���ҷ>�JI��P�d���ܪ0����η�}��>|����о8!3�`h��q���H�B��Lr�q��>�O?z�?{Nb�T��IWO�J���腽�e?�{g?m�>"O?C?H(���t�^}���>�=��n?\��?x@�?[>�=�鳽�2�>�;	?�?u��?y�s?B�?�^�>�FW;��!>�z��K]�=k>���=ґ�=b?��
?��
?[����	���y���]�7/�<��=ᶒ>I1�>�sr>�_�=� h=���=��[>v��>C�>�d>�'�>�c�>����lM?�,�<�:?F�?��>.�>y�q�W5����佅x���Ƌ�y��1E��N=��Y>�?=� ��J��>6�ɿC#�?���<�׾P�?�Ӿ��c���=��>��)���
?�E�>��ǽT��>"�(>[.�=T`�>$�D>63>�t����z`��v\�@����[�>	���1�&����|���mb�췾\�ھ��p�g���D��k3=���?+�+�QKG�q?&������?^�>zM5?���%�<� >1��>�.�>cC��^��'h���Ծ�*�?f��?�;c>��>H�W?�?Ւ1�23�vZ�+�u�n(A�-e�U�`��፿�����
����.�_?�x?1yA?�R�<,:z>Q��?��%�[ӏ��)�>�/�'';�@<=u+�>*��/�`���Ӿ��þ�7��HF>��o?<%�?wY?@TV��Խ.�>y\E?�B?K�?.5l?�P?J�Ⱦ�H0?(q��ظC?�?,-;?h|N?m?�>>*��=��>6y=n�μ�����s5�opw�ㄽ�=9->�}�=a����f=F�＞�/�y���ڒ��U0���m=�=�/�>�
;>���>S�]?��>�>�>�7?"���W8�z���b/?�x;=���۵��Eϡ����>��j?��?T5Z?xc>�3B�=%C��>�s�>��&>��[>���>v1�]�E���=$H>�P>ץ=��N�\큾c�	�O(��.��<��>ہ�>�p>xA���{>��=ފ�Pz>��=�oS��B�V��uK��:��F���T�>�H?�R?kd�=�=�[W���.i��i,?�f7?x+R?�ޅ?*��=�?�18�7aL�gx?��X�>�a,=0��Q��E(���V>�a|�{�P>b쩾Ϯ���^>%7�����t��E�?߾���=l~���U=r�������p�4��={�>1���!�������LL??��=�{��D/�6�ʾJU�=�>8o�>��3�U��:�)���/�=���>��N> �!�^��E;I�]���o�>��U?�R_?���?��H�pQ:�lf���ž~�������T?��>��(?��#�-�<�۾37.���Q�*����>�Q�>h���<[d��k�����y��ݐ�����> �?��>:\?��X?�A?ڪ?z�?/#�>S���ـ��k�&?w��?���=����,B��r!�5�I�}	�>6w"?#��-�>vr	?�)?�*?�zO?0?"}�=�o ���E��Ѝ>�>�]��;���zQ>�M?�3�>�YX?B%�?jxE>�c4�Lɶ�������>�B>p�+?L?��?�3�>.��>=줾���=���>AVc?/��?�zp?Ȯ�=z�>��$>&�>U��=+��>׭�>8�?zM?]|t?ǐH?a�>څ�<�"��/#���WR��Ќ����:�C<ٳC=��
���g��+����<��;ͨ�6�������a�T����%�j<`�>�s>A ����0>��ľ�E���@>E٣�4K��QԊ�\�:�e��=���>��?���>�\#����=:��>�G�>d��}7(?��?�? ~ ;R�b���ھ��K��>B?I��=��l�:���+�u���g=2�m? �^?��W�����'`?�e?��b�AYH��G���`=����?by�>m]+���>��a?��?���>��Q�M)X��r����\����(�=�w>[j#�����9T�>��h?#��>P�=>hN�=ڪ���'|��� �U?�ڟ?��?��g?`@>�uI��ο�u������8f?/��>:$��eq?�Jq=���Z����L������q��r����Ғ������+���S���Ӳ�=(?�w?)Sc?5�p?���cbb���d�D�����9�	1�����@�ƝB�ߎE��?v�7-����Q=�����=%Fc�``D�~��?�?���S��>@�_���վ��!W�=4����o"�yĠ=Z���_�=Zb*=b�%��9�����gY?�%�>�a�>�F?��Y���;�/��&E���\[=>���>�9�>�|�>4�.��GX�Y"��!�ھꃍ�s`[��o>��a?��5?]`�?�(�=I�������[�y�>�`��7�>C�><i�>��þ�ă��-���P���h�K�������Cݾ���=�=?K�n> �H>���?��?+�*�è$��B�������'=�n�>��l?
�>��>w�⼛F�E��>�Bi?g� ?��>*���!������{�w��d1?�8�>��?aI>�p��(`�WM���7���{J��M�f�{?�d�5���9=�~L?�Ԕ� �>�"�=���=�� �������=�7�>>B?�5��5�=��p������a����ξ%(?��?������1�ݎq>�0?�
�>tg�>Q��?Ĭ>�ó�ȇ���?�sg?��N?�6?�h�>�O3=7Q�4�ܽR[���=u��>��^>'J�<�$>{�B�3�5�i{%�u�o=��>�ϙ��,��G[��)<q�"=��=�g8>�>ҿ��B�2�ྣT�~&�4�⾉MX��
�]���#���¾�^��G���Sν�[K6��O<�L䐾�Y���<�?��?����������A�������_�>*��H`���s���hн�Hq��=��&��&�H�b�g�}�w�3/&?3����-ǿ���l��?e_?�hy?q���� ��7���)>>p�<��ɼ���ʚ��ο�W���^?wN�>7R�^���U��>Y��>7GR>^�j>
抾�Z��V�<*�	?�3,?��>	�}��ɿ	���r	�<�n�?�S@dvA?��(����+NU=���>�	?�@>$,1�Y�O��\�>V0�?���?V}M=J�W���	�2e?><��F�c8ܻ,�=X~�=�=���|J>:I�>���B?A��ܽE�4>(̅> �"�½�>�^��"�<yM]>��սh锽�\�?��U��a�d#�Q����?=^Cl?)�?��=�?.j}�%Rѿ̼j���]?��@���?�:?�P�� �>w���T?�L?X�E>�W+��m��s>�F�=��2�?�վ�B�a��5��><�=o���f8�ێD�yUݼ�B=]8��釻��#��]'�`�,=0�=IH<�;��Wl��L����������;��>L�=�� >�EE>m�g>��;>�}j> �H?? f?{H�>�*>�K���5���˾�����N�ԚB�}�V�]߾��������_˾#l�݉�����8m��6��{M=��Z����y�)���S�t84��A5?�c�=�z¾!�V����=����Dʚ�O:ٻ5���FL¾��5���y����?)�G?XՋ�4<<�1�&����*�����_?ʡ�����~Tʾ?Җ=q�<MH�9H)�>wVw=�6��4>��5Q�u0?5\?�����^��o.*>�� �*�=��+?'�?*Z<�&�>�I%?�*�u1�Z[>��3>ף>��>�3	>k���V۽J�?�T?�������[ܐ>�`��ȿz�]a=�7>275�R�鼑�[>�D�<����V��R���R�<�(W?{��>��)��ia������X==��x?��?7.�>h{k?��B?�Ԥ<!h���S���oaw=�W?7*i?��>����	оa���@�5?�e?d�N>�bh���2�.�SU��$?�n?*_?�~��"w}���w���n6?�?}?��g�ī��� ���@�>ɧ�>���>m�E����>�3?�Q��3(��Q���� 6����?u@@#tݼ�B����<��>�@�>�
��
��AL��F鲾�o&�P8�>�̾����"�d��A?�Ґ?=d?�ɝ����v�>������?��?`���#<���djc�������=į½�ce����:���ƾv��nM��|,�<���>)�@+���?�·���ڿS׿�^��r��.�����>8�>����\����s��]f�/cR��o=�OW��R�>��>d��������{�D^;�����>*���>��S�X.��sy���K7<9�>���>3��>ZA���������?\��%@ο1�������X?kh�?�m�?Pp?A*:<��v�.�{�-�4G?�s?AZ?�c%��$]�(�7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.���_?��a���p���-�
�ƽ'ۡ>��0��[\��Q������Ye����OMy�]�?g^�?�?Ǫ���"�]5%?�>`����,Ǿi��<�t�>�&�>1;N>&�^��u>6��:�WW	>���?0~�?Zn?���y����N>�}?��>��?���=���>8B�=:Ͱ�\j7�?�#>�%�=�JE���?�M?�>�>i�=��8��'/�ZsF��ER�����C���>
�a?.aL?��a>�a����0�T� ��#Ͻ�1��2��v@��,��B߽�J5> �=>�>��D���Ҿ�� ?�%�QLֿ����Nj�?Ҋj>՞ ?����-��}�<��`?Bu>`*#��H��>r���۽���?�D�?��?���/h#��q	>���>6�>,�Ž[F���<����.>��9?i������ev���z>��?a�@�>�?�Ch��*?5�������@Z�i
�c���2�=��(?�<˾�ŭ>���>�!i>*�u��Ź�(�y��{�>Z�?u-�?|�?��n?�����H����=?�Ra?�?[�7�j�$����=X��>G�������}�ВT?��@��@�I}?�����ɿ$����a�+ٌ�B�R<�]����>�讽�v=r�b= Kؽa��=�S+>	�>%�g>3Bh>ܛR>1��>���=��}��) �l<���猿
nZ�ɴV�H�
�A������)�m��K���s�������ֽ�Ӵ�n�g��� ?�p4�=	RV?��Q?�o?D�?��F�j�$>�W�[W"=B�%�=�x�>%3?�N?=�)?t�=-W���kc��A������ ㉾N�>�2R>��>[�>�L�>S�:��D>��6>St�>'�>Pe=�~�:��=��J>f��>J��>5ո>e�8>�x>=��������#o�%n�������j�?�U��dpF�+��Ӫ���������=�r.?��>�J���"ѿ�y���IH?2����]��0��{�=��%?�GO?�P!>ނ����J���>�%�`�f���=�.གr}��(*��9>a�?܉U>\^}>3�A�"�*�|fj��=žMmm>��C?Χ����9���x�b�'�\);&�F>nE�>ü�J���=����3��">��6?QD?�Aҽ�J̾ۊ�����@��>�xS>w8>��=N>H!����rQ������́�=�r�>C/?�
)>'<�=���>����p�N�p��>�C>�a'>��>?N%%?֐�\����1��rn,��)v>N'�>�h�>h�>�`I�� �=��>�md>t�
��ԅ����<C��LW>i�z���]��u��v=����x�=���=�W�]�=���,=�~?���(䈿��e���lD?S+?] �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��L��=}�>	׫>�ξ�L��?��Ž5Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿf��>���b���	��/d�"�W�>�aF?Zﾰ����t��?��>1/ �3T���ʿ�2s��k�>���?F�?,w���-�9�o/�>.��?��K?"J<>U����E�O��>M�5?I7H?W�>%~%�r8�?�o�?Ic�?�!x>N$�?܁?=��>r��<�qB�c﮿VɄ����>�u����=��0���@������E�|���R��2��?�W@=���>��}�ӾW6>>ŏ��ҵ��������>��>��w>3~g>���>KҪ>qj�>_�&�� ���MQ����@?�/�?aK��.��U�;�"?|9Q�R�Q>��=?Bt>@�����:;=]�?^�?�r?��>��
�]�h�����v����=�`�<��
?��>�W��?
�����=�5A>��y>4$�=l8��-9�(4n<�̹>��?�R�>���=7x ?U�#?�*l>8�>iD��'��NF���>�C�>n�?�V~?�q?JW��*!3�����顿}�[���N>�Ry??�L�>�_���C����E��z=��#��9d�?��f?��ὡ=?G�?��??��@?$�d>�!�|ؾÍ��6��>��!?Mp��A�1u&�I��ɿ?�-?���>�o���ս�lԼ{��G����$?%\?�&?
��Pa�Mþ���<����zr�� <XDJ��{>��>�g�����=>���=pgm�V�6��m<s'�=�\�>��=�6�{荽J�,?N�~�u�����=c�t�[�D����>u�V>�þ=J\?��P����f��#���":�у�?U>�?H�?65��b6i��>?뫆?�?�%�>����P�����p���~��M�D>�,�>���!�!����U��( ����Ͻ�
�k6�>��>n�>�,?�>gZ�>�z@��**����*���n�����1�':� *����FU�����7��l���׺�>߁ý�s�>��?��l>2k�>ET�>JeY���>�O@>���>�Ķ>�_>�3�=�2 >р��k�н8R?�B���T'�m>��,��\8C?��c?�>��f���d�ˆ?�ʒ?旜?��x>5Wh�:/+��5?�K�>2���h
?+f/=s���|<�Q��K��؅�Q�����>)�ؽ� :��HM�;,d��
?:�?�����j˾;�սU�\��F�=>�?�>?�L*��bL�uF[���W��3������s�W갾� �	Wk��m��q�o��Lq��(��p�>�?{��?�ᾔn˾�'���i�������=��?��>|�>�/>�(����[TP�ق�����q?���?	̊><>a?�-?X�=?i�[?,��>	��>a�,���?�e�<��>I5?�G?��U?h�"?��?�?Σ&>R����9��y�ɽ3?�w@?ש.?�l�>���>}���	-��?T��^�=���<�ڶ�\(�=����ɽ�v�����;��O>sX?���_�8�����k>�7?���>���>����.����<r
�>��
?�G�>c �A}r�<b��S�>M��?y�1}=	�)>(��=.����)Һ�_�=����s�=C���p;�8S<%��=���=;t�ݹ�����:F��;�j�<�P�>�?淋>j�>�o��U4���{G�=��\>��S>�>'Rھ2���@���
�g�C)v>��?4��?\(t=���=j��=hݠ�a��������+��<�S?�f#?��T?[}�?�=?[�#?3>��L���7��C���K?=�+?�'�>r���ɾ,8����3��?��?3@`����� )��࿾`vֽ~�>+".��~��ï�6�D��Ӕ�������!�?@b�?M;���6�ݷ�-�������mC?���>�(�>��>_*�3/h�Un���9>���>^�S?[I�>�>P?Q�z?��X?�U>!�4��%���{����H�i�%>��??���?Aɏ?n�x?QZ�>,d>��-��ྒྷq�����f��
q����6=|�W>�1�>
,�>1ϩ>���=�t��5���E��Ť=��j>�q�>�d�>�8�>T�y>���<��G?���>�]��6���줾�Ń�\=�5�u?ɛ�?��+?�Q=k��)�E�lG���J�>ko�?���?4*?��S�J��=��ּ6ⶾ��q��%�>�ڹ>�1�>aƓ=�vF=b>��>���>')�@a��q8�iTM�l�?�F?���=�*˿����o�J��EVs�D������0mi=����=�ڱ���������v�=�
k����e�nQ���Z�x�0����>���=��<5.=HD=��)=�8o;�-=!{�<K2=�z����<�j��rn
���W�7ǩ;Ӽv�Ƌ=�}=��¾]c}?<G?�!5?�RC?St>���=��ļ��>d����?i�P>6�3�j.ž)�8�tY��	��u;߾Vpվ��T���� �>X=k���=4�'>���=�K=�ŉ=0�s=+ڣ=hr���%=���=	�=
��=���=��>iL>���?2e���׭�)(�q#�\?U�>�	�=4��;�7?G`�<��i�?������So?�*@��?�o%?�T��Ӄ>ȘC�\�='p���(����>�K�>�W�<�U�>		>��=������}����?�E@kn?NL��eԿ�t>��5>�>|�R�i�/��wL�ūd��L��,"?s`;���Ҿ�%�>P�=��߾O_¾���<?D3>�g=��$�b�]��=i����d=6`="��>XI>��=���G��=y�)=���=�K>���;@�H�)��=Yn�=�X\>�B!>��>?�?`0?{>d?�)�>ǭm�k+Ͼ�I��TG�>M]�=49�>f�=�B>���>��7?ˢD?��K?�|�>;��=,��>��>9�,�M�m�g徙ǧ����<ܐ�?�φ?�˸>��O<��A����dO>���Ľ6o?�K1?�s?D�>�0�C5ʿ����:����@x�!Sr>��>������=�竾A�>�yX=s�>>��>�Z�>�=��e>�=z>{#�>�)q>���������=ȌW>�����=7��<;\	����;�Y{=ƫ[��󸽗�����<�J�<�Q9�R	�<�M>��>�߂=ë>p�">⥻�z�s>��O���R�ϔ�;�����S�o�d���k�3�,�'K���ek>O�=^�	�����n�?am>i�P>x��?-i?~�>5���I���T��;�L�B�y�>N�,> �Ծ�N���a���S���ﾄ��>��>��>u�l>�,��#?��w=r��\5���>E���L��m7��8q�t@����3i��ZѺ5�D?kD�����=�~?�I?���?���>bQ��w�ؾ}K0>pJ��ĭ=���Cq��S����?�'?���>���D����������>��9�0-]�ࣖ�6�*��ݡ<��4L�> ���x��ߒ+��\��ͤ��Y,L���{���>�6c?;�?rC��I�x���E�(�B�H���>�Q?��>��	?�2?т��]뾮p����=��u?
f�?���?f4>�=�䵽r�>�?���?���?z�s?��>�3��>0�o;�� >j=�����=C�>)�=���=�?�t
?Z�
?b����	��P𾞳��5^�'��<��=< �>�A�>�r>��=�h=]��=6�[>0ʞ>�͏>��d>���>7s�>��}�' �K� ?ѥ��܈�>��"?�	�>Z3a>_f��M�M�� ���ͧ�Ӕ3�주�����m�*F>�h����*f�>#MĿb��?�T�=@��>?�e��=���r�8=�^>�O���	?��>�
>�)�>u��>�br>-t�>Ǔ>/����G>�`��V�l�]�rU^�2�ž�z�>���a�!���cw<�\�;þ�O��4u��}�N��=8-�?$����K����!P����>D�{>�x
?$�v��}5=�X�>���>"�S>d��ܿ������>�ľ���?���?%�h>��>�?[?�L?�6���J�ٝ\�1�v�\�5�r5`��'`�E����r��[��O�yX?��n?^�>?�6�=�Kq>'E�?���J��/��>�#,�}O@�
�=V�>Hm��2�k��!ܾ�}پ�q���#E>h?���?�a?�N��0?��P�>;�P?:.X?�ą?��:?��M?�ž�/?ֳ�;(U+?�'?��;?�Oa?+v ?�/+>$w>��E��{����Ϛ�D׼=��������G>�09>� ��r��<	"�=[��;3|���<M�n��\,;�N=��=�X�=�Ʀ>2�]?��>�ن>n�7?�F�T�8��Z��[s/?�8=�"���֋�x������(>�pj?��?��Z?jf>��A�x|B��x>�щ>}O'>I[>j�>t��C���=&v>��>���=[J��^��
�Bp����<\>��?�T>�|ҽ2t�=�Z��D|��j�>�:۽��Ѿ)�O�K[�RPN�E����$�>ä^?Q+?k�(>C�ҾE���7m�T52?7)'?x�:?��?���=����[*>�GhQ�2^�Q$�>�7�=����[��������U�r�i�ӈ�=j⭾*u��_b>�/�(�rp�Z�H�Eb�:�u=��f�=R�z;�}����=2>�����"��ޗ�詿�M?SP�=M���O��b���
	>/,�>���>��:��{F��D��������=px�>�hI>�|��]ﾲ�I�֛�+��>͚<?�V?>Ek?[��ѠN��i�FQ��'P���2=?�b`>OI+?�s!=k� ��iﾶ����a�+[=�g�?�>g�� ]z�����<�� ��s;�=�2?g�>)�>�2?4��>?�:@?ZY?���>�>��;q��zA&?��?3��=��Խ��T��8��F�~��>!�)?�B����>��?^�?`�&?�Q?T�?>�>� ��C@����>RX�>��W�ob����_>!�J?ꚳ>�<Y?Rԃ?��=>P�5��颾sة�}b�=*>v�2?5#?į?���>��>s���)[�=J_�>�mq?T*�?��x?	!�=���>I�=�?�0>��>��?� ?�&B?NUd?g�@?^~�>��-i���Kt�'-𼰪ڼ�>�<J�<<}P=�!����	�����2=�8������(�\�
i��>;��<G^�>A�s>����c1>m�ľh;����@>+�+S���݊�4l:���=���>��?H��>�V#����==��> P�>����6(?Y�?;?ִ;�b�۾$�K��"�>	B?ݦ�=+�l�������u���g=d�m?r�^?~�W������n?��O?;����t�wL��۪��_�(�g-:?`"?�3�����>�u?C�?��>�A���^�����l�j�����>�,�>f��.k����=W�7?9�(?��>`}q�R*ؾo�Q�άd����>�ݝ?Jo�?D�x?���=~�]�ցϿ�ݾ�Ǌ��o?i��>i���{E?ݼ"���imb���Y�S�þ�о�v��T���G˾�K*��U����v�1>]�?.�z?}r?��l?!���bv���c��Ǒ��k(�&߾=L5�
�L��U��{8��E{�r���>����j��*�O>�[~�[�A��s�?�.&?��,�Հ�>ů��hO��U;wsD>����¼��=���Ǒ0=�GP=��b�	�.�g7���} ?�(�>��>��<?&b]�z�>�1�1�X8�����7>T�>���>�O�>Ps;�4�0��a˾`A��^C����u>��c?�	G? /q?/���f,2����L�A����q��!�L>��=�Ӗ>.l|�@�G�U�-��B�j�o�����鑾��	�:q=��3?	�>�y�>�?�?��~����p��6�9I=���>*	[?���>���>Ep��;�/�9��>Ñs?���>n>����>���̔���YU?� ?�y�>��<�=�ǀL�&��WD��0 Q���<��?{}��[~{��fW=��k?ӊ>�c彂�9>7��>�[�tM6���^=�Xy>�(^?��g�<H>?>��R0�b*�����
T)?\L?˒�}�*�f.~>�3"?gu�>��>@ �?N�>=Uþ.�?���?��^?7BJ?z:A?��>U`=�沽�aȽ��&���+=2��>��Z>xal=6��=U��y\�ɋ�ѽD=�K�=�ͼ���<f���j�J<+��<�3>�տ��N�s���'����H���[����#��:%h�Fd�^����I�AaR�y���x�G������@Ë��Rq��$�?�"�?�y���g������O	h��T��3q�>�.W�Q����վ|噽ϛ���qP���>
��0[�pZx���O��-&?p5��eͿ�H��V���u�>ǣ*?��{?e���k�U���Q>S���yL��ݹ��,���tͿ����O?:�>ʳᾏ���'�>jO>ʙ�=�kd>ň�������b>;3?*?���>�Ԥ��ȿ>�ſ_=��?uZ@�|A?��(�p�쾘V=���>2�	?U�?>QS1��I�����,V�>�<�?���?��M=8�W���	��e?��<��F���ݻg�= ?�=O=���L�J>�T�>��RA�"<ܽA�4>{څ>��"���6�^�4|�<��]>��սv9��eՄ?�r\�f�ϟ/��T��Y�>*�T?�>�=u�,?KFH�xzϿa�\�0a?'�?���?��(?I���vؚ>$�ܾ	�M?bM6?�ؘ>,c&���t�:u�=p�߼)������'V�-��=ˤ�>�>�=,�ǐ��O����] �=���ƿ��$�i��,��<>�Ǣ^�)?ܽcu��ڦf�߈���g�	���g=)��=��Q>{`�>m@V>�V>��X?&�k?�>�I>S��>f��3,;|���ۀ��C!�?ދ��}�Z��[��e�ܾ����^���?cɾ�6��z=��k�pS��cg1��P�s1���2?O$>g��Q�j��=�X��Hƞ�k�X</@p�<ﾋ;?���c�(�?W�Y?�`��8oF��K*��IýY�=��S?���f�߾]
���*>�琽�Q6=vܾ>�N�=�Q��J��u0?R]?K~��^��g*>N� ���=�+?��?�Y<V&�>�K%?ݼ*���㽮v[>̥3>ã>̥�>�	>����S۽�?y�T?��������>�c��\�z��Da=�B>
5�z��[>i�<�錾��U��S��~*�<�(W?���>��)��ia��Z��W==��x?Ӓ?�.�>T{k?��B?�Ӥ<h����S���x`w=�W?Q*i?��>1����	оH���8�5?ףe?B�N>�ah���#�.�9U��$?9�n?_?:~��)w}��������n6?��?�Ra�����C�뾞f*�⊈>�&�>�U�>�t�c��>|.?��L��O��_�ſ^3��5�?��	@x#�?��,�M��>���>���>����m���='�����S>�Y�>�-��#Ј�Hz1�+4�=JK?�s�?��,?mA���)����=(C���?�w�?J��0`�;.}��k��[�����<6�=ꍽ��S�I��F<���þ�6�C?��̢<z:�>.�@?,����>]E8�Xk῔�Ͽ2e���sľ�b��<? ��>I"�rƤ��ij��4l�j�A��;=�Pz��W�>��>�֔������{�>^;��l����>����	�>��S������U���R3<㴒>���>Bz�>a���<Qə?�;���1οg���6����X?ta�?�Y�?�u?To=<@�v��z��2��HG?��s?JZ?U�%��t]��a8�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�g�|=�>���>g>�#/�y�Ŀ�ٶ�>���Z��?��?�o���>r��?ts+?�i�8���[����*�m�+��<A?�2>���I�!�C0=�UҒ�¼
?W~0?{�f.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�i�>���?A��=���>'��=*m����'� >���=�N@��v?BDM?k��>�/�=M�4��U.���F��R����B�C���>ʳa?��L?�$a>���y�)�Q� ��ʽg$0�^�׼�L>���2�Gٽ�M6>T\>>�>��E���Ѿ�c-?Õ!��ҿQ㓿}F�X")?��S>N�?w��p�9��ս��_?��b>r+3�����s:��k�U{�?!6�?/??�z���8��$.={�?|�>c�ٽʯ��b�����;�8?G�A��$���s���5>�k�?�=@���?Nr�yo?R^�煊��-~�{����#�9x�=�#;?Uf�Z��>��>��=�q�w𰿍.x�T;�>	H�?���?`��>�b?��i��;����=��>�TV?ud?~5u�������=*�?h"�(l{��^?�@b@g�\?UP�����8������ʕ��7�<�a��fL>|l�s��=x� >f�7�U�E�G=>>��>�L>L�:>w�U>aR>>�>aց�7J#�����좍��O�C���o�h�X3�E�_�|�	��Ɨ�&Eξ���y�;�?e�P`V�f�!�Y��A1�=Q�\?F�]?�{�?��\>�����C�>%�7�@�>���ܩ�>���>�pS?-Ew?{$O?��i>TGǾQGw�����K�����%��>�ߤ>i�>�h�>2>�>U�^��(.>��=���>��o> '��>�9��fs��p>խ�>J��>�1�>��H>��> V¿����:U���p��sj�;�M�?�}����?�]��v����x���N�=��=?+�0>�l����տq}��!_U?�c�8��a�s�ϼ���>�lr?*+>�렾�!>�u��io����Z'/=��P��ξ���*9N>��?��g>Rv>BM3�Ɠ8�8�P��ǯ���{>��5?!˶�Ն9�i�u���H�5�۾��M>.��>�BK�������]t�"�i�e{=_�9?��?B���mԱ�C�t�\Ȟ��@R>A�[>u=�3�=-�M>�a�@ƽ)�F�t�+=Q��=�^>�V?��+>A��=Wߣ>�[��(-P����>́B>�,>W@?L,%?�s��ۗ����V�-��w>�S�>��>`>�VJ���=at�>��a>����Ӄ������?�:�W>z�}���_���u��x=�3�����=��=�� ��=��&=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�c�>ph��Q��O�m��a���ݽ�$�>��P?^;޾��q>5Е��?���>���u���&)ҿ<�s����>�R�?�`�?W��Al�?�K���,?�W�?_��>��>������>�b.?~bH?eIX>�O>��V��T�?�	�?j!�?�C>sҋ?	f?1F�>G=U(�oI���[�9���R�{1�>����FE��9[�+������l����t,>C+=#N>�1��ھC�)=�W4=���mSU;"V�>�[�>t�!>J�>��?D}�>��<>Ҩ=�~����~�BD���XV?|��?�f����ص�9hu>��o��$�>�X�>�K��O���Y7>Y.�?l?SUQ?O�=w�*��ޛ�u-Ϳu�ƾ��
=e
;=?�'?��I>�A���s�>���0*���=_�>��c�������M�F=1<�>r��>OW�>���<�-!?�!#?�|>��>�+9�%���Z�Q���>���>H<?�w?��?�����0������Ӡ�t[���4>�>q?�!?q�>9���Gá�����%�h���y?�h?������?ⓐ?p�:?�GL?cۓ>+>��Aپ����u>��!?���L�A�#j&��)�e�?�:?���>\t����ս�ּ{���*���?�%\?E!&?���P:a��Kþ��<�t!�V�f���<6jG���>H�>k����_�=��>\+�=�m�76�Ufc<�#�=�v�>���=@7�L����2?ب���J���{Q��3h�OV|����>�=%>���Q�M?����/���"���Ԋ�3e�5ƪ?� �?���?�<�V�y�͉T?R6�?�-�>�n�>�2��:۾�i�iή�1���Ω����:���>�=�e���d��ӳ��@�r�[�1��==�N?>�>��?p��>2ŏ=s��>��N��5��u�L�¾4�i��t8��>4���0����8{��Z�� ��S]Ǿ�7���O�>:b��4�>>�.?�M>N�>7�>���=5�>a��>c��>.fH>�]>X�<>{>�����䜽�KR?����]�'�3��ܱ���3B?Dqd?'1�>�i�􉅿 ��q�?���?9s�?�>v>�~h��,+��m?�<�>n��!q
?pT:=�*�<�U��8��~4��2����>�G׽� :�}M�nf�:j
?A/?&��0�̾�=׽������m=ܽ�?��)?��)�rzQ�#Jo�^X��PQ�R(	��i�QU���!%� �p��>��b���{@����'��Q=x#*?	É?�&����#����k�_jA��<S>Q��>��>���>�C>�0�)1�R]�m1%�m���/�>2}z?�9�>3�H?�1=?�PR?b�M?*+�>*�>�;���T�>~{����>��>8?�2?�2?+�?o�&?�MX>:8�����Ծ��?:�?�[?�` ?2��>����਽�iK�+ݻ��x�}������=5��<�ܽ����<�W=j`>X?���z�8�]����'k>��7?`��>"��>8��P9��	�<��>��
?
Q�>�����vr�M^��U�>X��?� ���=)�)>��=�Ņ��lк�N�=	���;��=�����;�� <0S�=^ɔ=��v�g/���>�:�Ɉ;���<el�>�m7?��>V��=�,�Ͼy=���Hg?�>�Һ��-K�����F���l{���>d�?O��?���>I>|l>�P��Kžf:#�)b��<�	?3�?-
n?Mw�?��0?^�??d3�>�K"��ᕿ�ڥ�6*쾅EE?Y�)?}H�>�;8��i��fT��w�\�:!?�6?�xD�m�<P!O��������=�n��Ɏ�x����+>�ơI=+m���n�?{Ɩ?>"�ݠ*�
?�Im���_����d?j��>]}>x��>�>�����9��g>�4+?�<p?���>S�O?FD{?��[?hT>�v8���љ��V0��!>�+@?z��?��?�y?��>Y
>Ȝ)�N&ྯ�����~����7T=�)Z>���>��>��>T)�=��ǽ�����>����=z@c>ͣ�>cZ�>���>K�w>���<#�G?���>1[����餾RŃ��#=���u?��?��+?�4=�����E�cH���G�>o�?&��?o5*?ϹS�	��=��ּ�㶾��q�&�>Kܹ>!1�>��=��F=g`>��>���>�$��`��p8�UM���?>F?ˤ�=�4ƿ�Fr���q�P��)I<d5���Td�y����Z�e�=�:���_����h[�E���=钾FU�����?{����>�˄=���=lY�=6��<�忼˙�<�0K=n��<�=_3p��"�<��8�>ọ���Xֺ�`< kF=�`
��m˾�}?ANI?�+?��C?LIy>k�>ݣ6��x�>7ۃ��O?��V>�N�_;���;��h��*��]�ؾK�׾��c�A�����>�K�d�>�4>i��=��<��=9s=:��=��?� �=���=ð�={ث=�?�=ID>��>��{?;|��x��9ZB������$?C��>�Ec=4Vؾ�
F?%��=����S���E�m?�� @�	�?`�??r`����>�7a����<z=� ��?!=�>��Z�??�>G�G>�&��Q����
�?n�?��@TsF?(퇿[\̿\�]>n3>�]>U"R���/�\X�XTi�"�W��!?=
<��:Ҿ�ԇ>��=k�侨�ƾm�=��5>S�i=���(V\�E=�=23���aC=h<p=��>X�O>�Q�=������=6T=���=QW>��(;g�M�1�!�l:=L�=x^>��%>{��>f�?��0?�#f?d�>y�a��=ɾ�����>\k�=���>���=��B>�c�>
A9?�#C?��I?��>���=�`�>���>�;0��/n���澶L��bH�<���?���?/�>�]B;)kD�Y��8<��EýE?�1?e�?�Μ>�z�[)�X�*�J�)���vX=y�>��=sA=�������1�=:�J=�_)>�	�>��>q�J>0D>�Q>̮�>�5	>Ҭz�.;sȆ<�__�����!�G��<;�������0��=�ak=��\�)b�-*=^H��0�V�����=��>�N�=�ϲ>͔^=iI��L>#���8h���˽���0^Z��0��q���2���#��>�4�>�6��S��͔
?��C>�>NJ�?�p?Qj�<�c�������Tz�=��I��eڼ�/>��N�I��Us���J�N-�Q��>J�>|�>��l>,��"?��uw=�\`5�
�>w�����n��:q�\@��l���	i��Y׺�D?%E��_��=]~?:�I?l�?��>�����ؾf0>BR��c�=9��q�r�����?�'?��>�쾎�D�v5̾����׷>VI�4P�������0�>L��÷�ᨱ>�����о�#3��g��������B��Rr���>�O?'�?�+b�P���QO�����慽gT?�ig?��>K?B8?Z5����y��d�=�n?۰�?@�?�>�W�=��5��I�>�$?���?"�?T�r?��)��p�>1*ýPU�>H �<��=��>tW> ��=���>=��>o<?�P�<���q�'����a��� �=1��=J��>�0e>��X>��G�d�;���='�8>+j�>�
�>G��>�Ų>�,j>^��`���?��=���>e�+?ZD> X>�|��_Gp���*>v懾�Ds�5р��v0�x�;�>�!�=8���8��>��ɿO�?"��=	�
�y?���� ���>��>�`�O�><?��z>�؄>I@>m�=�
 >�>\Ӿ<�>� �Q!�&[C�V�R�EiѾ��z>C����q%��������^I�܇��lI�f)j��1���8=�V�<�<�?R����k���)�����N}?��>$6?Ќ�7N���>��>�ȍ>T�������Ѝ��2� �?6��?A�x>E�>��o?x�?�d��h͊��or��됿���E��3l��i��a͕���,���$�E?x�y?mH?�ue>d>*��?[02��t;�?�����_�i�G���>ॅ�*��	(�s�����In>��Y?�L�?I�a?2��e�Z=�3�>jL0?��k?���?17�?�n?s�/����>�����0M?Z�=?O�>yMd?Y>?�E>4 �=���<n�2>�5����S��i�OK���k>�Q+>A��=S��=�vr=*�=I0=�7սm+�ތ`��Vû��[��4�;�}�=�nF>�r�>��]?-E�>�c>�)@?���XD��a��B<?-��=�ֳ�Q����Gξ:K ����=�e?�I�?�Vl?�l>��7��y�=��=4�U>r�>�e|>U3�>�}��T���7=:->�w�=ɨ%>��S��
v���
��ϑ�O�=D>���>1|>S���'>r}���Tz���d>��Q��ݺ�-�S���G��1�s�v�mM�>��K?T�?=ڙ=R龁4��Mf�3)?�Z<?�NM?��?7�=$�۾F�9�T�J�el�t0�>�< �����~&��C�:�ə�:k�s>�<��^⛾��_>U,�Q`�1n�:�C�M�d�=U�s�v=��ubѾL�m��%�=��>�����!�P���;x��cuJ?�[=͌��8%P�q��n�>*�>j��>s���eY�7A�֭��pܐ=�^�>�>>����=�yE��g����>�RA?�4S?O`�?`jN�V�x�O[���'$���)�=�A?���>[�?!��%���{�/)��T�3�.���?4H�>d駾e�y��xM����7��)�>�c?E��>��?�[?=}?
_]?L"?�Y
?���>/`����9'?,��?��=&S�<b�40��QJ����>�5'?[�#�(Q�>I�?u�!?��,?�T?��?�+�=���A�B�P��>�6�>�EZ�qe���%Q><\I?�ζ>��Z?C�?��M>�7�\����|���>�=��->2?r!?Fp?6!�>�d�>V`��nj�=���>Dc?s1�?��o?�W�=?�u1>�5�>�=^��>ɧ�>�?p,O?Ƿs?��J?x�>��<�"��]/���r��N��
�;f�Q<e{=�����s�-��s8�<�+�;.���|I��iV���D�	����a�;�_�>��s>U
���0>V�ľ�O��K�@>H���P��ڊ�(�:�޷=��>��?��>�X#���=�>I�>?���6(?��?�?�!;�b�'�ھ��K�$�>	B?���=��l�����|�u�n�g=��m?��^?��W�V&���\e?�S?&�1�l�H�}��-�O�;���=?}��>�q�=���>�*b?���?d�?l��k�j�m閿2Eu�4�j�>��]>��ﾚݔ����=Bs?��z>��>e�=��{�1���c#"��F?Q�?�?؍�?�L�;8�U�TĿ����B��[$c?��>U��vH%?�<�X������@X��C*۾U
��!b���E������$0#�����.|#���=��?�3x?̂m?��b?H��r�k�]~^��ۅ�LwG�:��:
���4��xN��aG�?v�ٍ����P���x��=��f���D�״?��?q�#����>�p��7���	U�&�;>����rS��ex=?豽�Wl=�Y.=��a���q��s����?%Q�>�.�>�;=?�[V���C��).��>��,侺*>ު>�0�>]�>�ռ��b�Y���c!ξmh���m�y�u>�d?n�G?��p?fzҽ��2�n����U �ۏ�GS��	~>>�X>s�>/�d���*�S�*�]�A��q�������\�U�^=s^4?�>��>���?�??�*�D�%y���.���=���>�Ih?�A�>�{z>�-ѽܼ!�0��>��n?��>}{�>���W�U��ꏿ�I�_��>U�>���>u�.>6	����a�����ݝ�9Q]����=�no?,Ы�����Q;5�i?N�>(�=�Y�>y+=�t<���E��?,�0#�>Z?�7��}�>Bɹ���&�9}��m�ƾ/W)?T?�Ò���*�#
}>�;"?���>T��>�$�?v˜>�þ+W����?@_?UeJ?>.A?���>�=�v���]Ƚ@l&�?9*=2��>6�Z>�wj=^��=���P�[�����E=���=C=ҼSr��/�<1����O<Y�<��3>�׿mH�k������V��H����x�o����������c=��\]�����6Լ4���U��u���p\�as�?���?�[��g3��1q��Jj�[M�	i�>7�X�&�C��S��f'n�'���i�����5�G�4om���[��+?o}����ӿiϊ�w�5�Q��>�*?���?v���{m[�?L�>Zm������^
�����пJ���i�X?s��>� ¾:>�S�>5�$>�팽D�>:�t�~�m�'kO>�c�>"P?Z��>_U[��
����ο�s[;	��?ć@�|A?H�(����V=���>А	?��?>�R1��H�G����S�>I<�? ��? zM=��W�*�	��e?�v<��F���ݻ��=�<�=�U=z���J>V�>5��>SA��BܽҸ4>ۅ>v"������^�C��<%�]>m�ս8��=(�?�Q[���e��1�]��;�m�<I?�L?����?��w�_�ȿΨe�X&[?,K @��?��@?⽡�Y��>���knn?�??�w�>S#�3%��4">��B����@N�	�E�Uѽ�?�ò>l�|��G4��v������$�=��������P(��!"����<�<�<��ټȫϽ����sȽ�-����s�M�׽�'~=�D�=l�j>3��>:�L>��H>>�^?��s?�L�>R M=41���fD��վz_�=�Ę����yB���	�!zd��a�
rԾ�F ��r�]�ӭ��I�5�@<Pu�f���d���?$��;���E?~B�<X6Ҿ)\N���=�q���A̾k���!���Ū���9���R�k��?F�.?�Ֆ���?�������<��u�w�d?�c���ھ�=��h�>>.`<9r]��M[>��=�+�)jF�i�N�x.0?	P?ū������M%>O ����<f�*?��?z�<��>��$?���A 潒1\>gI:>�"�>��>���=,����Խ��?.�X?�v�������>��ƾ(w�#=v>��#��
j��xV>��<\̊��`:~⡽��<�(W?ϛ�>M�)����a�����P==S�x?ߒ?%/�>^{k?��B?9ɤ<9h����S� ��]w=(�W?d*i?�>�����	о򀧾��5?��e?�N>�`h�/��0�.��T�&%?n�n?�^?�~���v}��������n6?~?ˣk��h��!M�+*��d�>f��>��>�X����>&r(?Y���8��f�ÿR90�T`�?o�	@���?�8L����<�w�>���>�=B�e���J��֥�����=��>�۶�'k��sH �I�*V?��?z��>�Z��I���>x���h�?��?�꨾��<lk
�e\�{H
��,<?�=������������9�~��������@��:��>_@ ����>��d�#��GпՑ�{���/�e�ު?!d�>�\��ľ�<s��gf�g�=��/��r��]�>
�>�R���$��,�{�P;�]���*+�> �n4�>�S��)��H\��z<<W�>5��>��>������� ��?T���=ο2���ơ���X?�b�?q�?�m?��=<�+w��{�.��v/G?�s?Z?Aw%��]�~R7�Y�j?Tા� a�j=4� �F�n�O>xU3?Dw�>�D-��Z�=>Ǥ�>��> /���ĿsB��̣����?���?��1�>�@�?^�)?x��8ș��Ƭ���*��"��C?�5>�l��L�!��~=������	?\�1?My���=�i�_?�a���p���-�}�ƽܡ>8�0�?d\�^Q������Xe�����?y����?G^�?I�?h��� #��5%?��>����	9Ǿ��<��>�(�>A*N>QC_���u>_�&�:�og	>���?�~�?�j?ϕ�������U>��}?�D�>NY�?*�>�7�>�-�=J���:7&��	>��E>�7���>�K?R?�;�=)��W8��,5��}L��#�hH� �>�KU?�?a?۸�>oҽFh"=��;�`���\�K�Z= `�Oy<R�B���>�>��?>����2���(?u�!�P9ʿQđ���A�?���>Q�?f��r���O��{ir?av*>$�%����P�����;�?٭@�
?+m�1>w$D=[�?.*�>xH���E˾#ǔ>X�W?	�.�"����!t��w�>��?�i@�۶?��U�;-$?	�;���@Dy�ֿ��C.��E9>}K??$r*����>絵>�#S>I:��PV��V~���>aC�?i��?��?ц`?i�|�(�V��I=��>Rbd?�<?��(#9����<��>[�,�n��!��KZk?��@i�@�e?꾿�׿\z���9Ͼ'rʾ��@=�G�<�#>�I����>뇽J�'=l
�f��=���>,��>��l>h<>�.K>��(>N����{$�[Ө�hu���,� V3��":��qh�zc�@��� �ф���Uپh���ӽ<�̽Z�d����޴��=n0k?b!B?�Ԋ?� �>��H���[>��7���9>��;�iݘ>%v�>7�^?oTP?��?ኝ<�-r���s��~w�/��?���l�>i�A>�V�>~��>��>8[��=�=|Q�>�Ad=/��$�=��<��=I�>�>]��>K�O>�^=�ÿ�^���o�{yϽ�$��y�?n���=5C�Q�<bh�����)ᐼ�?�J>˜��Jѿ����x�b?b������ =r����>шv?ޚ>�m/�˗��3Q6='��������.>9�7��r���F�_F>M�?A�f>dhj>�/���7���N������	}>�8?3��%6���t��J���۾,�H>�`�>_�Z�,�.9��th~��(c�?q=��;?��?M5���ݲ�Q�t�����kfQ>s<[>:O,=�h�=��G>0�g��Խ��C���=k�=P`i>�R?A�+>iP�=nģ>gV���O��~�>�B>>�+>�	@?�%?N��-���҈��g�-�� w>�?�>�π>4>7J��ϯ=Q��>�	b>]J��0�����@��lW>�~�5_�תt��gx=l2���E�=�;�=*� �3=���'=�~?���$䈿��Ve���lD?G+?� �=u�F<��"�E ���H��G�?r�@m�?��	��V�7�?�@�?��Z��=�|�>׫>�ξ"�L��?��Ž*Ǣ�Ô	�.)#�eS�?��?��/�Wʋ�5l��6>�^%?��Ӿ��>\��ڒ��W���ubw��1=��>�'I?��� �B�ެF�F�?��?������Sjɿ�w��E�>wz�? q�?�m�~����O@��N�>�H�?�7V?��c>�u۾�bK��6�>�??�O?�R�>�O���'��?�(�?>|�?MVI>HÏ?�Ge?�k�>"�(;��4����������� =ck��lp�>�1>�䮾�
J�&��@����}�o�H{`>]�T=NØ>�|a��F��#�<#����⫾q袽.K�>��>E%b>��>��?g�>'�>D	R=2�u�\�a��M��e�N?}�?�����%��+9��`�>j���teU?m�*?�O?:i��	=A�?��?�z�?j�;>�1�)���'���]������=�v��m�?s��>�T��9l�>!�۾ e�=����;2�>>6�Ծ�m��9.�kg�>^�?��>�Ʊ�� ?tL$?=q>��>^=C�PĒ���H�x,�>���>W?�d}?\?�ݽ�ذ3�A���3���'[��X>��x?<�?�ԓ>�����v�������U7��C��z-�?i�c?�˽"�?��?h�A?�>?j�b>���tz۾�`ȽLK}>q�!?�&�j�A�&T&� ��?�D?���>�~��Ekս+�׼Q��Zb�� ?V+\?z5&?���0a�3þ���<?�"��6Q����;�F�	�>S�>7������=�>��=�;m��[6�Ҧe<A*�=���>���=�7����|=,?��G�܃�(�=��r�YyD���> JL>���۪^?6t=��{�k��w��RU�_�?ˠ�?�j�?v��Şh��%=?��?�	?b%�>=J���|޾O�ྺSw�Xx�u���>-��>��l�q����t���+F��ƽ�b����>��>\:?�$?�BU>�p�>?���>����La�Iwg�e�#���=���8��#�K��P�B��'�ƾF������>�㸽�o�>V?!�5>�$�>���>յ�<�;f>Lr�>,�>%�>E�h>%��=)��=�]�1�:��KR?*�����'����a����3B?�pd?2�>�i��������?Æ�?}s�?:?v>�~h�-+��m?�=�>E��>q
?�K:=�E��1�<�U��ӻ�0����ī�>cG׽� :�pM��mf��j
?�/?Y���̾�9׽���qن=ԩ�?��*?1�+�frR���e�FrX�O�K��r,���^��u���_/�ϕ��0��V�v�ר{��[.�8�>+&?�)�?���￾�p��j���9_�p�$=88(?\�>a�>o�>@#!��3��Y�����1�A�?v�?�>&BL?ۏ8?�R?��D?i<�>e=�>�o��#?Mɦ;��>:��>e�C?aG*?w�,?�?��$?x�6>e-���ʐǾ?��?@?��>��?좾��Žv�����<��p�Bk~��h�=(*�<����W���6<�w>�X?f����8�`����k>Y�7?��>h��>���I-��8�<m�>�
?�F�>K �.~r�c��V�>���?�����=��)>���=:�����Һ+Z�=G���R�=u4���y;��g<̂�=+��=�Jt�" ��)(�:Ǡ�;�m�<�n?u�'?H�>6^j>��K�AW3�%(8�U�>�")�>ܤ�>֨=�!3�qߖ��ω�ǽ���Z�=��?���?p�>��=e�=Vf��q���W�4��<$����?D�>?\n?��?�fR?�P?��>���������3z�D�?a�-?>�]��ʾ�J�� �6��s?`�?��\�RU��2��%��H�����=�8��f����_8�ћ=K}��f��z�?�[�?����3�~y���5��_F��@S?���>���>���>��,���e�;����}>:?�:^?���>C�O?12{?b�[?�T>;m8���Dԙ�l-�Ϗ!>�C@?���?[��?�y?b�>��>l)��-���V����.���x�S=��Y>���>�9�>N#�>�P�=N�ǽy����'?��P�=�b>Ky�>>��>>��>�x>�Į<w�G?���>\��e��줾�ǃ��=�B�u?��?n�+?�C=����E��G���G�>�n�?���?�4*?�S����=?�ּ㶾��q�q&�> ڹ>0�>;ē=��F=�c>��>��>v)��_��q8��WM���?.F?b��=��ÿ�Cs��d��ؚ���w<Ӯ���(a��ra�S�e�i��=�ԙ�9�&�Y2����]�j:���ߑ�o����ԡ��#��ř�>�y\=n>���=ߚ�<��	��<� =���<�V%=*�W�;�<�L��Ze�	���''����;��/=dl'<��ʾ��}?0I?�,?Z�C?�|z>��>�N��4�>Y����?-�W>w�5�#��޹9�
���盓��eپ�ؾ}Uc������	>��]���>��5>fV�=皳<�?�=�q=��=����
�
=W0�=8|�=���=��=��>�}>B�?�������Q\��P��/4?NE�>
6>�3�8fE?A2��su�$澿*�'�Ě�?��@�a�?��%?�?�>o>�a�~q�<���;�x���4i=�J�<s<=��?;x=�l4��͛�9\��c�?uJ@�M?�,���ڿ��>]�7>>��R�}�1�`�\�S�b��iZ���!?�P;�/O̾^3�>q��=�/߾"�ƾV.=��6>�Ub=��;W\���=	){�`<=�l=�ʉ>��C>�]�=.(��w��=��I=���=�O>د����7��:,�<�3=���=<�b>�&>׀�>�?�c0?�_d?@;�>��m���ξ�\��W�>|��=�n�>L�=b�B>���>�7?��D?r�K?0p�>�K�=���>�#�>��,���m�^����e@�<痈?Y͆?0ϸ>�N<I�A�¢�JQ>��Ž{p?�F1??z?՞>)��`�ο�w1��,������J�� '��Ǿ�?3>!�����$�(<Wd��oD>ϝ�>с>ܪ>�[�>F>�<�>ۃ(>��»\�<�]����=�{�=��=6�����3���ս��<� +=)j�<(i<��=8�=\���4��|��=T��>(�=�=�>�OK>���U>�ߋ�S�j����a����d�}t�4u�8�3���ԽqzF>��!>U*��E��k"?�>��8>f��?톇?I��=�����|������!)=�]��N�=����ӫ�#N�n�d�k�G�����>��>�>N�l>,��)?���v=~
�yT5���>q�����~*��<q�TA������i�(�ںt�D?nE����=�~?�I?G�?ю�>鷘���ؾ&0>�z���J=7	���p��{��?�'?ޅ�>�(�r�D���˾�߽��>gH���O�Ε�t�0�gT.��p��mq�>����#ѾdJ3�Jv������uB�Tr��ܺ>�O?ծ?w�`��R��_0O�����*����?�g?�9�>wG?��?�^��P��%&����=�n?e��?�T�?4]>���=����S�>�9	?�?���?�s?M�?�X|�>���;(!>D"�����=3�>q��=U��=�o?ȏ
?��
?�W����	�/�����^��G�<*�=���>�[�>1�r>t��=��g=�_�=�\>�˞>�؏>��d>��>�:�>;������!?�Tw=%�>�w=?AZ�>�1H>W����C�.��j/��GZ�JDH�'䦽ޅ�����<b$�n�k����>��пo�?�t�=�Z��?<�پ:>�ǎ>��>N�h��3�>z"�>�~�>?��>��r>N��=��>��Z>�Ҿ��>�Q��E!�ہC�#1R��VѾf�{>E���ӽ&�����6I�����wc�C�i�N<���m=�畺<`D�?�/��-gk�pk)��N ���?���>��5?�:���舽�K>�|�>��>+���5����������"�?���?�Ê>���>��X?�K?=�^���ƾ*2f��3���p��A�2Xb����ݞ���&�˔v�H7?Y=i?��@?Wbb>;)�>�Â?3�2��0��p'�>�K3���V�b1}�Gp"?^u�uʭ����)�׾m�;�
>�)??���?�hP?��:����?��d?�Y?�=�?�1U? ��?q���9�%?�k���?Zt?�Y?UU?�_�>��=u�R>�s>q��:�UB�uȪ���#��ʽ⦅=C�=��@=g_=�OY��젻�S/���<��
��l��N��'�;�!A=F��=��
>�*�>��]?���>!7�>)6?��)��:��ⴾ�1?O�C=7������[���3��2`�=7�g?p«?�[?n>�5>�]@���>�*�>*>��Y>��>����>�(i�=i>�>j��=k*��8���o
�3ސ�!=�$>�@?��N>/˺�yr>D���g�ξ��>�uQ����d^����[�C[�}_�����>CTN?�4?��E>��޾�à��{�L�C?/�5?�J?%��?��F>�oʾ�A�$IF���A���?�����������5���-T�*���A>Ԭ¾wj���q^>g���&���s�SW�6Ⱦ��m=����.�=�
��~Ծ%'�� ��=�(
>R�о�s�F�� ����O?B�=@x����.���ƾ4%�=��>ٽ�>����Ľ͆C�������=3D�>�->�*a��:پ�{>�=Q��q>��>?��a?{��?�΂��dh���G�Z���;۾y	�:c�?)��>�?�,�>�I=p���	��i�k�4�B�SG�>G�?�)�GwB�D|C������*���>�T�>٧�=S�?��5?���>�|]?2?۴�>���>�e�S����G%?ܖ�?ˇ=@ؽ&�P�bp8�v�F��V�>�(?@�A����>`�?�?R�&?��P?��?Zc>o����2>����>Rg�>�W�E��D�a>�I?�X�>��Y?�߃?m=>v�3�)Ǥ�"6����=�>�3?��#?A�?{��>��>&Ѡ���=�P�>l2c?]�?vko?���=�%?�l0>���>S��=;�>f��>)�?w�N?gs?x3J?s�>��<����ݹ�[ox��Q�/G�;#p5<j�|=�� ���q����F�<SM�;!���|����F�r����
<v�>%�s>(2��E�0>�ľDJ��E�@>%���'|������:�᰷=g�>��?[R�>�[#� ^�=��>7�>���j/(?F�?#�?��(;�b�?۾/lK�<�>o�A?��=��l�!|����u���h=��m?�r^?߉W�����6�b?�]?h�=���þ�b����g�O?B�
?��G���>��~?d�q?��>��e��9n����Cb��j�Ѷ=Pr�>X�K�d��?�>Y�7?ZN�>��b>�#�=;u۾�w��q��T?x�?�?���?J+*>W�n�44࿍���L��M^?[��>5@���"?i.���ϾDQ���"����K������@��?x��ɮ$�����׽��=��?�s?~Xq?c�_?� �ad��0^�I	���kV�@&�#���E�W(E���C�:�n�hc��0�������G=�-r�R�]�S��?�>?�/��M�?�������@���z�>��ľ��>��;}>�Ϝ<�[>9y�>L��ǳA���ȾW�?4��>���>�8>?�=7��,�y� ��(M�b)�,�=�S�>��>���>0*��,��`Z�ei��v��/7��O�u>6nc?�K?��n?�~ ���0��m��^�!��.,�$4��&kB>�7>F߉>O�W�����x&�� >���r�+��Y|����	����=��2?�j�>�>�w�?�#?�	�}����x��X1�`c�<�.�>I�h?���>�g�>��н=!�Ú�>��l?��>h%�>FS��uL!���{�)�˽�T�>I�>]��>4p>	{,��\�)L��C�����8���=�h?����pJa����>�R?
�:��P<]
�>b	v���!����(��N>��?��=�w;>��ž_>���{�!a���?6�?2M2�uE�|B�>.�/?��>�>��v?>�{Ǿ�p%=�??]M?�9?�]?Z��>�������==�ɽ�^1�k&�=w�K>��$>�Qz=��w=ݷ��;���=�X���̅r=�X���Tv<M�.>6�L=���=/>�)>��ܿ��O�G�a��"b��0e)�/$���+��o���=�*���T��X��!�Q���� z��*�t���o�9��R�?�w�?ڃݾ�X=ѵ��8��(ξ���>=�b���`=e�����=$�����f���.��e;�F:�&��Q�'?�����ǿ𰡿�:ܾ3! ?�A ?:�y?��<�"���8�� >JC�<�,����뾫����ο>�����^?���>��/��c��>᥂>�X>�Hq>����螾�1�<��?/�-?��>ێr�-�ɿ_���¤<���?/�@��??q�$�$")��J�>���>�P�>��>|�ܼ#�7���
��j�>GH�?�Q[?v��>NZ��Ғ|��;H?���=�a`���=�=�<��=�,�r6�=}��>zD�=0��=�s����.��>�\�=`ӗ�(/	�y���� +>��]=1RW��&�<5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=v6�ꉤ�{���&V�}��=[��>c�>,������O��I��U��=�h��ȿ��#�"�#�7Y=<�;� �꽈0�����\��In��w���}�=Z�=�O>l��>�(]>�b>[V?&&j?(K�>�3>'��:ɑ��IȾ�/��1������;���p��qj�����I��'>�0����������<�	�=�XR�h2���!�MGc�+�E���.?k�#>��ɾR�M���*<^�ʾ{
���N�������̾H1�^9n�(ܟ?��A?B���mV�&!�˳�����SlW?g�����iB�����=-��M=���>�=�1⾲�2�x�S��.?��?�������8S9>^?��A	=�,?:?&yL;*ة>��#?��������J>�=>]k�>,5�>��>/2��K�ӽW]?��N?׼ �ٚ��1�>�M��BN��R�|=���=V�9����@�a>+��<�����:�b�����<W4W?��>pA*�S��Bf���6��8A=��x?��?�-�>z�k?G�B?+G�<�|��yT���U�s=W?$sh?�	>�Ԁ�8ZϾ������5?��e?�L>��f�_|�I�.�8��y>?Uin?�g?�Ӛ�ݮ|��������\6?F�v?Qr^��s��j����V�(=�>K\�>���>��9��i�>Α>?s#��G�����QY4�q?��@ʍ�?��;<�6��=6;?t[�>̮O��>ƾ�q��G����q=%�>���lev����OT,��8?��?^��>����&���#�= ݩ����?�ʆ?7Ⱦ�[�=Q
�駇�������=n�=iߜ=��/>&���a ����;&��ؾ�ݽ\w>�
@��8����>1�=|��1�����x����O��4#?�N�>�Z��zW��~������w0	��#@�lm�:��>���=[)Q��Q���S���e�b�>���>9���Zx�>����[s��鷾O1=Y��>�M�>��>b�N=?������?����ʿ�0�� d�l?T?�?�I{?�P?��h�p>��I5�o�"=O�o?zE??�3?)��<��?�n?!��j?�^���V`�C�4��GE�DU>7#3?�G�>�-�h�|=.>���>�Y>�%/���Ŀ�ض�!�����?��?�m����>�?sq+?k�U7���W��u�*�I!+�>A?2>�����!��/=�Ғ���
?�~0?���-�Y�_?.�a�E�p���-���ƽ�ۡ>�0��e\��M������Xe�	���@y����?L^�?j�?��� #�a6%?�>d����8Ǿ��<���>�(�>*N>�H_���u>����:�i	>���?�~�?Sj?���������U>�}?�>��?���=��>Z>�=·���-���#>a��=L�?�ߚ?d�M?f�>���=49���.��AF��AR�|����C�Y�>�a?6cL?�Hb>�	��%3�q!��ν�?1����h`@�Hk,�>߽�]5>�U>>�R>��D���Ҿ��?Kp�7�ؿ�i��)p'��54?3��>!�?'���t�^���;_?=z�>�6�,���%���B�X��?�G�?;�?��׾R̼�>D�>�I�>��ԽS���G�����7>-�B?���D����o���>���? �@�ծ?Ui��	?���P��Va~����7�e��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=7M�>Μk?�s?dQo���k�B>��?"������L��f?�
@u@a�^?*�{�yҥ�Q�Ǿ���0�=�%�=�kp>�e��gd�=�˝�o�8�Z��[&�=�p�>�N>1*>���>��9>��>Ã�Mj%���� _��u�:�}D�4�	�%�\�| ��������µ���kž՝&��(�<*P=�S��^���,�)}�=AHU?�R?�p?D ?z�t�{Y>�����=�Z"�q�~=��>&2?�>L?��*?ᬓ=q����d�Z<��bi��Q2�����>t�H>���>?��>:�>��T:ױH>Ux?>(��>�%>��-=`����
	=ުO>��>��>�ƹ>�F<>��>Jϴ��1���h�>
w�̽W�?]���l�J�P1���:��#����a�=�`.?z>����>п%���72H?�����(��+���>�0?�bW?��>k�� �T�8>)����j��]>�+ ��~l��)�7!Q>�k?�g�>�A)>ϵ0�+�(�#�_����D�>
�-?j�m��d��w������e��VF��8>W�	����������t��ċ����n	?��	?[���:q����#m���n�>X��>`8���e�=��S>Q�=���UoڼGT�x�K�tV�=��?G2,>�މ=ul�>z����"N����>�E>E�,>�??��$?��������@�.�tv>�B�>e�>��>P�I�}ï=�u�>��_>���,փ�?��93@��~V>�hp�Qdb�DT{��{=uy���p�=A�=FS��ޗ>��Y%=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�h�>�|��[�����u��?#=x��>�5H?`X����O�>��{
?2?�K�٨��7�ȿwv����>� �?��?��m�|@��c@���>w��?zdY?h~i>�l۾�Z����>7�@?�R?�'�>�@�w�'���?�ڶ?���?�I>���?.�s?LP�>�w�L/�0��؏��o�=��U;�m�>d>^����eF��Փ��b���j�����b>��$=��>�J佷A���A�=�닽�K���7f����>'q>`�I>mS�>� ?�R�>���>u&=�[���܀�;����K?���?(���2n��O�<��=0�^��&?�I4?�k[�}�Ͼ�ը>�\?i?�[?d�>7��O>��?迿4~��)��<��K>"4�>�H�>�$���FK>��Ծ�4D�ap�>�ϗ>�����?ھ�,��CO��KB�>�e!?���>�Ү=�� ?��#?[�j>�(�>aE��9����E����>΢�>�H?��~?��?�Թ�iZ3�����桿Y�[��;N>j�x?/V?jʕ>a���ă���mE�~AI�����Q��?atg?�U��?@2�?܉??\�A?�'f>����ؾ鶴�T�>=�&?�E���F���#�����/?0�?�(�>2������q�N����wa����><,Q?X_?W~��2Y�ןþ��<�����"�:�':���S@>��.>Q���+�=h�D>��;=$���H�8�ƶ���=�Ņ>I�=��Q�����=,?ֽG��܃���= �r��wD��>sML>2���^?l=�:�{�����x���	U�t �?}��?�j�?�����h�a$=?��?�? �>�J���|޾����Ow�zx��w���>9��>9�l������/����F����Ž�����>�r�>d�?���>ԪW>$ç>)D��iK��޾�e���`�^5���7�ۆ'�3��9S���I��dZ��ʾ�劾���>��U�q�>��?��D>�m>���>���<,�>��y>���>��>�Q>�O>�}�=��=�ٽ�T?��ž�1�ۡ־%����5?�b?�?M���#��{@߾�H?���?��?���=�db�6'*�.?-�>6.b��&?��=�ý��E=^����g�]�üci��t>)�7���I�SpF�*��m�?X�?�E��0ľ�Z��\���v;o=gN�?M)?��)�S�Q�A�o�2�W��'S��.�kh�>0��״$��vp��鏿�T��!"����(��)=��*?�$�?��ώ�⬾:k�{?�F�f>���>��>e�>�HI>��	���1���]�hK'��]��+a�>~Y{?��\>p�H?��<?ݍK?��V?s��>*��>��ྪ�?l7=��>W<	?փ6?�N?+A?�)�><H*?�/d>�+����X��F�?	�?�"?�?�vC?�
��' �Jr��ӱo��"(��t�<�~�=�γ��#[�y2���A��y=�8?�� �+����ƫ>F??t��>���>P8o��Nz�Ss=4�>?g�>5��ŅU����HL�>C"�?"奺
��=��>3/<�dd=�W�<�r =yY���<�	e=@<:�����=>�zB=���;ق@��m��w�Z=�]�=�u�>��?9��>?C�>[@��� �����k�=�Y>�S>,>fFپ~���$��$�g�]y>yw�?�z�?��f=��=��=�|��@U�����&�����<��?(J#?yXT?ȕ�?��=?�i#?�>�*�PM��M^��f����? g,?4Ð>&o���ɾ��2��?�?3�_�?�r\*��ľ��ܽ��>/�.��K}�������D���໺��������?�ם?C�E�t�5�b��g������oC?��>I��>i��>�(���f���=5>���>��Q?R��>��O?�%{?�[?�S>��8��$���ə�qJZ�:Q">��??嫁?��?CGy?D��>�>+D)�qR��"��E��a��G���lP=�T[>�0�>D�>�"�>x��=�`Ƚ�;��Bt@�$v�=D�b>���>n��>{��>�Vy>��<�9F?aP�>�'��� �2����.���5x��Ct?�/�?��*?,`G=�
���F��A��+�>-F�?�Q�?<,?�-M����=��ļ4�����r���>LP�>�י>���=�}�=3�>2�>�N�>Q��G$�"�5��R�{?\�G?׵�=o�ſ��q�$�p�����Sh<�����d��s���)Z�.��=(���wM�4Y���[�
���Ղ���㵾@���0T{�ݷ�>6L�=�Y�=��=u��<��ȼQͻ<�pJ=R�<�a=Nn��l<D]6�kջ�懽�&7�n`W<�J=���#�˾�E}?juI?;,+?�bD?m�z>��>�t9���>[���A�?��X>wG�?N���b9���3���Hw׾�rվ�c��s���>�-I��4>�Q3>�r�=Q�<���=�Zl=�&�=���h=�=l��=Lܯ=u�="�>��>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>@��>�}<=ɣv�����E�#��?lԽf�c?&7H�Ȏ/�4��>�5��t(��? ��8d�F�=m�������'T�i��=��L<�&�<�W�mUC>i�>>�I>�ἣlj>h��>k�˽&iM�L�.�����>�9>}�ջ/U>�;�=^�o>��>�f.?��$?��9?���>+в��v�|跾Y�$=y�>��?E�%=�B>���>�3?��F?�3W?��>�U�=z>�>%��>zs1�4 w�~�p�Y켾�-���%�??��?,�>5�">�Ǿ�Y[��W=�0�=p�?b�V?��@?K��>�a�<A�o�#�,7��}��}c<}4�=�ip�{�g��'�4���"�i�>:�>��>jܜ>6��>�E>^z^>��>�	>��<���=]�2��P�e%�z=D�aIg=�4,��c�q� Xi������Y�#w$�'rJ=��<˝�=��>�m>��>GM�=�����.>?��ҒL�\7�=F1��-�A��d��=~���.���6��C>}jX>~��M)����?�Z>Ս?>.~�?*Mu?+!>�����վ�G��&xe���R�ֹ=��>|�<���;��l`�N�M�&�Ҿ���>�ώ>���>��l>�,�7?�H�w=�L5�"�>i������d�I3q�/8��*쟿\i�K��=�D?_D��E�=6.~?s�I?|ڏ?��>�b��I�ؾ�l0>n0��K+=b���q�{W����?�'?lm�>E����D�-�̾�]���ӳ>�?���P�\���g.�����f��F�>n'��j�оD�3��n��m$���C�*zr�S�>4=M?~L�?�M\�[����LL�2e�!��rv?�7f?r��>?z?>>?S�������y�C\�=T�k?_�?��?���=�xo=�+=[A�>X�>�(�?�?�AO?�1O�=?k#ӽ?h>)r�<�B>\w>���=�d�<��?���>��.?0�`��ξ}����0y�t\=�8<���>���>JdP>6��=�ʏ��>��=5O�=���>&�=�U>Ӭ>�ჾ�n��1?̈)>S6=ܢ;?~��=_H���c>�_>K���P�[(��Y��Y����@>��m�L\�}�*�3��>Hཿ?��?��k=�U��?Wv��~P<N�p=�i�>�D�=ٟ?ּ�>k��>��>��>�j�=��>��=FӾ�~>V���c!��,C���R��Ѿ�}z>����	&�����t��CI��m���g��j�.���;=�鸽<(H�?}���
�k���)�U���l�?�[�>�6?vڌ������>��>�Ǎ>�I��Y���ȍ��g�c�?���?~:c>�>��W?U�?�1��3�cwZ���u�2(A�fe�Ǹ`�+፿Ĝ��f�
�i�����_?��x?�yA?�c�<y8z>Ӣ�?H�%��ԏ�+�>8/��%;��T<=-/�>�(����`��Ӿp�þ�<�YKF>W�o?%�?a[?LV�"���|k>O?��?^�?t:2?xw8?��e�&2
?��<�>�y!?�A.?\}?�?'yɼ~5>A\Y=Ɇ#>�-���Ba����v��>]���=qA=� s���Qc�	��=	���E���P�=Ar��R�=��=q}�<��:=u�k>U߃?e��>���=� 4?������j��\��o�:?.�>U��9>������徰]�>K�f?w��?���?�!�>"Y'�#�k�H\.>E��>xWl>��>���>�}���>U=��=|��Cפ>�n>�t��@�2��%'�'��10
�F�i><��>R�{>-ٌ�U(>�飾��y��>d>9+R�;���>S�DH���1�_;w�,��>��K?��?K��=��龋$��Ff�D�(?C�<?�CM?��?^��=��۾��9��J��Q��ޟ> �<���<�������w:�1��:t,t>���&���˥l>�9�1i����k��`��gžh{{=���d��=����tȾ�^��)+=B>�+��G��"��T7����J?<��=�������MȾ��>n�>֧�>Q�
�+�����?������=n��>�g�>��r��Ͼ��*���{9�>h�=?[zW?D��?n-�c���V����������L�"?�� ?�A?�P�>p,�=�u���}$�&f���NQ�Hd�>PP?��4���7����~d�0t:�z��>��>���k9?K�c?���>�ve?;�4?�u�>�M�>��>x���j�$?w܃?�oz=�ݐ�-%��o5��_Z����>	?eΎ�+U�>�H"?6�?�z*?�AZ?E�?�(�=��޾�19�%��>!�>�mU�(��%d'>(8?9Ȫ>�YX?ք?��9>�"�Ǿ#�)���<�xF>��6?'�5?�0?`��>P�>�ń���=e��>:�j?9T�?x3t?�w>~�?r�>7�>2��=��>���>�?��G?�8y?K>?�U�>�p`<�]ν���:O��R4<]D�<��v<�~=#c����W�Nv��#.G=��7�ۼW���솽��B�/���H����>M�?>��V�>����������>�
>�3ž�ː�l��a��<���>�#?�i> �X�k�t�>��>w}��?n�?xN?d����%L�~���i���`�>�G?x��=խv�',����t��=��j?S�I?[kJ����Ͻb?�^?+��C=�Y�þd=b�!1���O?��
?�uG�┳>�~?��q?���>��e�(&n���b�P�i���=�e�>�7�V�d�@(�>J�7?WW�>$�b>�h�=V۾��w�XȠ�'$?�ٌ?���?��?@�)>.�n������ ����\?z>�>�֧�(h"?V]�F�ξ-�������^Eᾚ��~����&��6��C#$�'^����ٽ��=�?K}r?
�q?2y_?l� ��!c���]��ŀ���T����P��fHE��bE�X�B�Gn�I=�p�������K=d�:��F�u�?��!?����Z�?-��i�������>`�޾�U��2K��+��M[���o~>j0��q�������?7��>\��>!�J?��)��]/�u��w�4������R�=�3�>93�>���>��v=�2��{n��5ؾ�����8��[w>�gb?h�K?Bo?QH���/��s����"�ʾ!�����~}=>E	>���>��U��p�K�%���>���r����ꐾ��	���=".1?�K~>���>�?^$?H��Y����t���0�w�u<���>�qi?�@�>֙�>i�ɽ�!����>A�l?���>�ޠ>⃌�YI!�:�{�ڑʽa2�>F�>N��>��o>Ȟ,��\��c��7��9�q��=��h?Nw��-�`�F�>� R?�Jq:R�I<(|�>��v��!�Y��(�~�>�w?���=1�;>�Cž�&���{��6���\?�]?ʘ�ۧJ�|�>T�1?��	?ң�>L�t?�O�>ʳ�&� �U�?�a4?�~F?�N?��>���;F��=�֪���-��"|=%��>O>�>�>�|(>����u��JD��b��ߢ==3w�=͠���:�>j==Bҋ��xA=�ֿ�PD�)�ݾ���y۾c��(K����	����)<��6�SR��𧣾}ĺ���'�8����|�����)�ѥ�?�1�?YL��v:�����Ö����ĭ>�o���A=�Wf���5�oܾ�ؾ�툾Ў���=�!B=�88Y�k�'?����;�ǿ䫡��1ܾ] ?,& ?��y?��ٺ"��v8�4!>�b�<����1�뾷�����ο̏���^?���>�4�����>�ς>��X>u�p>��������<X�?2j-?���>A�r��ɿJ}�����<���?��@��@?��&��R��0@={��> $?��8>�!������~�>�H�?���?��=nX��zG�i�a?`�;<��F���}�==Nv=�7����P>8ۉ>Ww	��]G�s^罐�4>��>�䤼�C��i�"��<�:L>�ܽcAw���?��\�ưe���/��i���>o�T?���>+ݣ=��,?�9H��vϿ�\���`?M�?��?��(?Y��4s�>��ܾ�]M?'66?�
�>Y6&���t��D�=,2��枻<��V�C\�=z��>�*>TC-�Z��bO�d\��Z*�=���ƿ�� �[�%���=�9�D'=��Ƚ���!��eSw��+^�ه���;��2(8=�<9>��N>���=T�w>��Y?�Zv?�ٴ>�->�\���Ӿ����[�ɻ���d𼃋&�	�g�����[��Fܾ�����8��Z����N<�
5�=-QR��y��( ���n��?@��C+?���=ۿ��%?�_��3ܾ���������wξ.F-�k�f����?�D?5Ć�ڬC�������|8��iU?%'����E���ސ>2I��D�t=�K�>@��=	�Ծ/�"�X�W���/?5�?F ��}��qK+>�I�(�=�)+?��?Ţq<ҍ�>ҽ"??/��i��y[>�Q7>A��>&�>�>����K۽��?��R?h
���e�����>�w���^z��=e=� �=��5�z��K�Z>�ї<�Ӊ��Ǎ�4����i�<��I?��>��Q�B#�#��������O=Mac?���>e?8=jU?�d?�U;=��ս��I�˪%�ڣ=L�D?m!?�\A>xv��۵����о�K?�%u?Ɩ�� ��<��H�G�݇��*��>���?؍#?����!�f��l��(��ԧP?��v?�r^�ss�����D�V�W=�>�[�>���>��9��k�>�>?�#��G������pY4�%Þ?��@���?9�;<��O��=�;?h\�>��O��>ƾ�z��������q=�"�>���|ev����R,�Y�8?ܠ�?���>������>�������?�o�?����1=�N��}k�W�Ⱦ��=f��;����PФ�8J�kF;��%������v����>G�@`N`��O	?8X�=��ܿ�ſh^���0�z���9?cN?W�C=te��1QF��j����Y�3#A��+��.�>ԣ>>�d���A^�M��Vw���_>m�>��.�E]�>�� ����E�������F?���>�>m>���=�X��@�?"+�{e���9��V��9�q?rT�?+O?�))?�J�[����}��d{=ߓz?&^@?G�
?#�=w���b��j?W_���T`��4��GE��U> 3?G�>z�-��|=�>~�>�g>!!/��Ŀ#ض�i�����?
��?�l꾙��>^��?1q+?ek�R5��PZ����*����\>A?��1>�����!�a.=�,Ԓ�н
?�x0?���+�5�_?.�a���p�x�-�4�ƽ�ۡ>��0�`f\��B������Xe���?Ay�r��?/^�?v�?��� #�6%?
�>>����8Ǿ�
�<逧>�(�>*N>�H_�c�u>����:�~h	>���?�~�?�i?㕏�����U>�}?h6�>��?H��=��>~p�=�����0��$>��=z�?�<�?��M?�_�>;��=e9��'/�,]F��@R�")�o�C�]�>��a?2L?Hb>R���N1��!��Kͽf1��N�j�@��-�m#�W&5>(
>>�>;�D�~Ӿ��?Lp�9�ؿ�i��p'��54?+��>�?����t�����;_?Vz�>�6� ,���%���B�_��?�G�?>�?��׾�R̼�>=�>�I�>C�Խ����_�����7>/�B?_��D��u�o�z�>���?	�@�ծ?ii�=	?+��P��o`~�,��g7����=��7?�1��z>^��>��=&ov�㻪��s�S��>2B�?){�?X��>3�l?ɀo���B���1=�K�>Лk?�t?�#o���l�B>ϵ?)������%K�� f?��
@Cu@О^?Z[���5���Ҿİݾ`��=�W<>S�c>ߴ���n=Yr|�)!�lW=
S>�>�F�=�H�<T�=D�[>��^> y��%�{������C��n�ku%�X�q����~���о5q��ˍ�Q<v�V���d��?=��`����=U?X R?�|p?'(�>�r��>V��\O
=�� ���|=%i�>{�1?��L?7*?��=�!���e��H���q��	���զ�>j�G>���>!��>��>��4:�J>	�?>�ހ>[U>˼#=\�$�=O>s��>d/�>�y�>�C<>��>Iϴ��1��K�h� w��̽-�?����u�J��1��"9��V���:k�=�a.?{>����>пR����2H?,���R)���+�$�>n�0?bcW?��>@��[�T�:>���c�j��_> , �[l���)�l%Q>xl?q�w>��c>��1�7L.�,�O��髾[l>�f4?����+%-��Ao��8M�f�׾b�L><c�>m���V"�5e����}��Uc���w==�A?2?�T�{��>.s�0���`^p>'�u>%CG��=
�*>��e�>ؽ��+�Ig<cq�="�`>�?.>J�c=��>����TO2�f&�> �P>��>YF:?�"?]{��DN��?v��O�C�d>�$�>��V>?�=�a=�ڏ�=�c	?V�H>Ւ��}qۼ����m���t�>;�<(��źý2P�;�7����=�A
>^�#��@U��S=�~?���)䈿��e���lD?O+?} �=��F<��"�B ���H��F�?r�@m�?��	�ߢV�?�?�@�?��<��=}�>
׫>�ξ�L�ޱ?��Ž;Ǣ�Ȕ	�-)#�gS�?��?��/�Yʋ�;l�n6>�^%?��ӾWl�>o�]�������u��#=љ�>�7H?9P��+ Q���=���
??�!�e���w�ȿqv����>���?r�?��m��8���@�m��>��?IJY?_�i>�n۾(�Z����>
�@?ER?��>mD�ۑ'��?�Զ?���?�I>錑?p�s?]m�>;x�3Y/�66��<����y=bi\;ra�>`V>�����eF��ד��g���j������a>�$=��>U:��3���-�=WꋽNH��	�f���>,-q>��I>�V�>� ?u`�>5��>�}=�i������T�����K?���?5���2n�)P�<ݟ�=��^��&?>I4?{r[�0�Ͼ�ը>�\?k?�[?�c�>H��D>��<迿~��˪�<��K>4�>cH�>�$���FK>��Ծ�4D�pp�>З>$����?ھ-���J��NB�>�e!?���>�Ү=\� ?��#?�j>�&�>,`E�l9���E�b��>T��>0H?Q�~?�?QԹ��Y3�F���桿�[�/>N>_�x?V?�ʕ>���ă��P�E��>I�E���.��?tg?�V�X?�1�?��??3�A?�(f>m���ؾ1���t�>�u?�\X�<��!.)�	p��Z�?�y�>���>���=9�=�����!�:��x��>}Li?]�F?�W�>[�J�۾r8>;Bc���=F=���!��@�=�fR>���v��=�-G>`��<�Ǟ�ϰݽ����?�E=z �>�>[v� �;�,?B�N��ꂾ�F�=$�r�P�C�^>M>K>�o����^?��=�|�l𬿷n���fT��&�?�x�?�+�?�괽�Mh���<?P�?�+?Փ�>����lrݾ��ྍ�w�s�x����>8c�>� `�#��ol������FH����ĽW����>y��>�'?��>��>&�s>|f�2� �2E������&W���$�����*�bl����{�Z;��L]ɾQ�w����>����.^>�?��t>烃>\��>�7�<��>~�X>.OC>��[>�m�>uG>�Ћ>~�=5�%�Q?A滾>kO�a?���8��t�?}o?� D?[����t��//ȾR�?Qb�?�)�?D�<�y��3�\3�>�8�>R�,�9;�>o>	�e>F	=´������U=OH����>P����[N���=�"ֳ���?�l ?�㵽^fܾ�K�4��z�k=�]�?��'?�w)��R��Bo�9W���R������Ta�L��D�%���q�Ǐ�;ۃ�����(�#�.=n+?���?������h��7�l�O>���g>���>�N�>�q�>�iH>��
���0�sG\��&�7*���>`yy?�s�>�LO?�?I?��5?��Q?��>;N�>�Ӑ��f�>l.��$�>N��>1=??f?�+?�C?zr/?@��>V]�<U���0�5)?'�?�=:?1?��%?�1Y�zWW��ҽW#��<N��m:>�+�=|�5;Ί���ȫ�����h�=��?ܫ��??9�F\�a�l>f2?�k�>� �>�팾���H�<�9�>�=?��>�����s�k�{�>�5?˼��(��<z{">T�=G�K��Cʲ=��<��:=�R�:?z����㼎�=��4=Xtf<�q�<� �{żr��<�s�>��?^��>5�>y1��� �B���z�=51Y>S>4!>Aپ�|��C!���g��hy>ly�?�{�?,�g=��=��=�q���S�����(콾P	�<"�?�F#?�RT?P��?��=?Hi#?�>�%��H��e\������?�0?��k>���N璾������"���>�:�>7�O��A��N�&�&<�|m���|$>/�>�K7j�D���ijA�E���y��Υ��L�?[P�?x��� �ʙ쾨����F��M?�F>C�>��>����
U����;Uk=���>a�G?Ս�>"�O?Dt?��[?J�d>�5�$���󼕿����>�=pMI?�D�?���?~|?:��>ý�=JD�U��"� ����M���G��w�F<�N>q��>6��>���>]��=. ����aG�N��<�*P>4�>�֣>Q��>��>ĉ=�tC?���>������g������R/���q?rp�?��?Z��=���{�R�l7����>�G�?PI�?�o5?��
����=��ȼV����4c�h�>ǒ�>}��>��=F�>$�t>��>~�>�D"��H�+ @��u�<�w?�<?99>�ǿ0u���t�#����ԏ<nN��Q W�n���'�U��ʜ=˳���B�=����_��5���"��Z��瞾�$z���>cA�=Q��=���=-��<�q�>��<��;=�T�<Q,=J�Z����;Z^�CU	���e8ڸݻ5<7�1=65л|�˾��}?=I?�+?��C?s�y>�I>q�3�s��>����<?�V>�cP����N�;����������ؾ�p׾2�c�̟��F>KLI�W�>r:3>}@�=iM�<��= /s=�ǎ=8kS�C=��=�8�=kP�=���=��>[^>�6w?X��������4Q�A[罩�:?�8�>{�=W�ƾ�@?W�>>�2�������b� .?���?�T�?.�?nti��d�>R��]㎽�q�=E����=2>���=]�2�X��>��J>���K�����v4�?��@��??�ዿʢϿUa/>��;>��>�T�_�.��R\�X$e��g[��#?%<��}ξ�#�>r�=�پ�N����=JT->%mJ=���90\�a�=���UN=Ns=��>�;E>1��=Vq��p9�=͘U=D��=��F>�����F�~�2�_�5=ta�=S`>G�#>�>�>_�?�?P�C?�j�>�:h�x|������G>���h?���=5��̣>	)T?�Y1?޷3?)��>F>�<�'�>G�>NK���q�	���雾7'�=��?���?Ev�>M�Һw���`�!�}�a�ƞ[�YX,?��_?��"?���>�!�D���(�m�L�r�^�6�S=2�<=E͂�î�zr���ؽu=fd\>	�>I�>��7>�<>�s>1�>��>��=~<��<h�<��<D�<��=��<�P=�v׼?y5:~���L=�ԃ�<��������&������w�=�3�>tB>���>���=�Q��T�/>2��MJ�=}�=N���TA�g�b��}�->-�=�0��eH>��]>5�k������E?2�b>��@>�h�?v�u?+�->aN���ؾ�����m�'�M�r��=��>E�8�4�<�`?a��N�!�ԾV��>-ۅ>ᑟ>F��>�.�Q�8���#=y�â.��9�>�E��Zg���$��~g�������bo���ۼ�;?������=]��?CrI?²�?v�>�L�����!J>��c�*3b����G?������
�?&u&? ��>���>�ؿӾm����>��7��#L������'�'y�9Z�̾C��>�ł��.׾&�?�i��+V����8�+���A
�>HD?6��?G������Jm,�T�����?�,c?��~>+<�>q��>E������`�F�W�<>�}c?���?�p�?eW=���=3��=U�?�QS>�l�?&%�?�r?.��g��><�;�}i�yd.����>�m=��������kB?i(?'T?��l7D����q��~�Z������%��E>x��>���>@C2>q��=Wͫ����=�hB>��Z>��=U�z>N4�>����f�w*?*�>H/>�r6?�$X>�My��~f�=$�=uf��Y��3]�W�Ľ����p=�n�Rb�<3�)�>�b���n�?�=PS�۳?��پ�-��n>�u>Eᙽ�]�>h�<>�)>���>���>onW>�>k>"Ӿt{>��+]!��(C�+uR��ѾԖz>������&�I�����I�V紾�i�&j���=��[�<�>�?Y��^�k���)�W����?a�>�-6?=䌾Q(��6�>ٲ�>�-�>\��ř��꽍�ۏᾌ��?���?�Qd>���>!$X?��?�h;�L+��Z��xv�i�=���a���`��|��*ρ�a�	�����_?��v?3�??�5<u>�~?��#����W'�>�{-�OC9�f�[=^�>�a��lX���Ҿ%¾�  �Y
N>�,p?���?�n?�Z�8i��r,>yg<?(�0?��u?s�2?��=?i���"?��(>Gp?�,	?�6?>�,?�9
?�,>C+>P��LK=Ԕ�G����ϽMs��H���<C=-�n= i�9�E�;+�6=�@�<����R��%�:����<ȓo=�Q�=��=4��>��j?�%�>H7>��"?�>H��2��@V���B?�{=N5�����l�M���>��z?ɱ?��s?�*�><[E�]�G���y>��>_�A>}�>��>�5T���'����=*�0�7Y;>_`>�� <��������d� �s�>&��>��z>Ƕ��(>�7����x� d>��R�����ƯQ�2�G�2���v�u��>�K?['?;�=��龵����f�)?ef<?�JM?E�?@ܓ=�{۾��9�ÎJ��)�㭟>-��<w��Ň�����}�:��T:��r>�����|�c>�R���۾�dn��hI�f6�p(a=W��K1M=����ؾ������=�>���ݣ!�SÖ������aI?X�h=�F���bW�^߾�o3>��>|~�>'�)��V��gA��䰾J�=���>4�6>Upd�O��LF�"%���>�>?�bx?�n�?p���0x��y�9@ʾ�S�j�!<�0 ?k�>�9�><�k>8�l=q�F��+;������U���>�"?�V��1R���E<�d!�?�7�ǿ�>���>��<cIJ?�c?"��>qmC?�Q?n�	?��?�aٽ���(?���?3�=Wϰ�p$���]�����K��>6h?i/:�68�>~5?���>�2?JPi?�}A?�\^>YS)��Y�p�\>R��>�Pa�`�ſ�U�>E'0?K>�F?��?�]9>|�+�H���O�콀����"0>�W\?b�[?tV'?�l2?�Y�>}(����\<�� >֢5?af?<im?s�>7�>|�R>cN�>����w�>6X?)�?6�?d;\?�a?�?*��<�}�Eժ���ۻ�	ͼ�)��`�=�ӧ=���7*�$��2�;��=�4s��V��$0q�G<k�1���,�?2�>�����>L'��:Ŗ=��B>�ɾ9¾a-*�G|���>���>��6>ix��9�z�u>�E�>:u��dK?��?3!�>@Gu���K��cz�rܠ�%4�>��T?�!�;�%��]���i ���%۽��s?9�W?�c>�f��ąV?�b?#g��\uN���Y��c��9f��q6\?�u9?GU�;�G�>��t?��l?֘�>n*��^�������c��Y��#F�=�W�>����bJf���>o�>?��>n'D=&.��13�;���ύʾ�Y?e�?Թ?���?�v|>|<I�I1ʿ3���>���^?A)�>�}��Z#?Z��Ͼ�,���؍�W%㾁�d��������>���r$�mZ���Խ=ڻ=�?V�r?�q?~�_?�� ���c�l�]����6V�����\���E���D��dC��$n��m�rT������9HC=�����I���?��?�m���2?6�ƾ���3м����>����w��>���T��<��=�yʾ�A������"?ᄽ>G�>"69?r/��>>�bp��7U�����-�Z>2+>n&�>��>{3<�7�K�0�_��	�i��3�ɴv>1�b?�L?��n?�+��0��΂�?J!��4��J���B>A(>3�>�NY�P.��d%���>�5�s�Z����x
��΃=�R1?���>~T�>��?bd?���U7��`"z���0����<�	�>�i?�b�>g&�>vFʽ� �`�>�(m?���>]�>�솾��'�y�๽h��>O�>�L?�Yx>�D*�Y�[�mɏ�������6��_�=M�h?������a�r�>/�O?���9=0x<�G�>��a�� ����4�&�oC>L)?��=19>�eľZ��|b{�8ۇ��-$?��?�,���?.��-�>��#?�>u�>�c�?���>�J���9����?�G^?�s@?�+?\��>f�%=�u��%ӯ����N�<ڝ�>N9U>�w�<
's=�-��in��H@��U�<[��=���s�����<9^s;���;���;#�.>�`ÿu2�U\徥����-p9�Q��cYc�xpټ@񲾬٫��������ZtD��������W�f�Q�/�F��?&(�?U���2N�ڠ��r��(���Vk>���>䨐�Ml�zϾ��ݾ�c2�R>���%��I��}���'?������ǿͰ��~:ܾ! ?�A ?B�y?��B�"��8��� >�L�<w&��<�뾟�����οV�����^?t��>���/��=��>���>��X>�Gq>���螾�3�<p�?@�-?Z��>P�r��ɿ���8��<���?"�@��A?�(&��F쾁�R=8�>�	?��6>4�%�����β���>��?��?.#\=x)W���&�p�a?SK�;��F�T�
�Xb�=,��=9�=���E[J>؎�>4��o�A�VCڽ�}%>���>
�X��&S��õ<��[>^;޽��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=7;��e����H#���"��<���<z��1�0�C^��/X�����5|�����=��=�q_>-o�>D\>p6{>ͫI?K_^?[R�>L�>����{x��1�Ӿ�L뼮�t����L����G���=��Vg��	�b�����ÅȾ%=���=7R�����M� �M�b�J�F�g�.?�t$>C�ʾ��M�#�,<<tʾxª��̈́������+̾��1��!n��͟?��A?�����V�����Q����W?B�0��v謾���=Ml���W=/$�>鱢=���3���S��+?�o%?O0���/���gw>l!����=��'?��?�E�<sة>��-?��������>�J>�Ǘ>��>��3>�㠾�����H?�Q?�-��و�E�>ÿξ�����<�V�=@:<��=�x�i>�Y8=K�5�I��$�� ��Xrf?�#�>h�Z�Z湾y�׾9�b�}�̼*v�?5Lm>/����Ӕ?d*C?|��H7j���L����dY$��h?��>�5�=-����D�������{?���?/τ�E�N��])��+�u�	�3v�>���?�^+?ƄA�����ݙ��_ؾ���>��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?n�;<��U��=�;?l\�>�O��>ƾ�z������3�q=�"�>���ev����R,�f�8?ݠ�?���>������m�=>nm����?�v�?Pξ۾=̇)�o�#���N>��[����$�=�|}$�J�����D��Ⱦ�t�`�>�D@�F��?�݆�d���_ ˿	�X� :���ʾLI?A1�>쁫��$�/a�n�U�δ9�~��[��,7�>��>T��$K�=�2��u����;�`�>>��>y'�}�b��O*��Z�1"�>��?�� ?\�M=�.��:�?��پ�!пf���Y��<u?5�?�$�?���><��؃�<��@@l<v�b?�B.?�BX?�Tc��s��߰�<��j?�\��JV`��4��GE� U>2!3?�E�>O�-�n�|=&>���>�_>�#/�;�Ŀ�ض�Q�����?��?vm�}��>g��?�q+?`l�Y7��qW����*���&��=A?�2>i���t�!�z1=��Ԓ���
?�}0?�y�/�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?t��>���?��=��>�>n/��'�v<ܕ!>�>b:��?�M?���>��=��>�UQ*�� C��IO����@��!�>$�c?s�L?��]>�Z��m�� �$��U��@
>��0�	�N�c�����#0>BLP>,�$>�-O��wھ��?Mp�7�ؿ�i��p'��54?/��>�?����t�����;_?Rz�>�6��+���%���B�`��?�G�?=�?��׾�R̼�>9�>�I�>N�Խ����Y�����7>/�B?a��D��r�o�{�>���?�@�ծ?fi��	?����E��V�}�k��f�:��q�=�87?��𾮃}>���>q`�=��v�ɶ���Os��V�>�;�?�R�?ۤ�>
�l?%�n�o0C�Q8=`�>.�j?�G?�eb��C�ZbB>��?�P�"��`k�v�e?��
@x~@ {^?�ࢿ�׿k���7�^,��c(=��C<�=+/��-Y�<羬<o��<��<L�q=�$�>E��>ᄂ>��>�
�>�(=>7P��e�)�>���-u��0 I�����k$̾<F ��0k�ۈ��fh��^�&�J�%���MVϼR*u��K ��t��A��=�U?�;R?��o?X� ?d�r��� >����'1=�($���='�>|Z2?�L?�>*?�ٔ=r����d��5���0���󇾡	�>�?J>@��>I��>>��r�/�G>n�=>��>���=�b(=���8�	=��M>�+�> ��>�.�>aL<>(�>�ϴ�r/���h�>w�F&̽��?������J��0���9������$e�=�_.?r>^��.>п�����1H?�����&���+���> �0?�cW?��>0
����T�4>�����j�&P>�4 �eul�g�)�� Q>xj?@�j>��v>�4�N[7��Q�ٰ�r�z>�M6?�.���9��u��1J�cX߾w�G>�*�>��P��������Ij�'Dh��}=�};?X�?��ƽ@�����q�7�����S>�}`>�=�%�=��J>y�u���̽ʭB��,=�z�=�=X>�W?�d(>�x�=���>~;��SB:��ݲ>��5>��->��?? �#?p�H�<,��S7r�S.��.`>���>١}>��>��D�Qh�=���>D.`>�p��䒽}�����*��	Q>�����Yk��7���=�3��Qp�=4Ұ=
l�J"F��=�~?���(䈿��e���lD?S+?b �=�F<��"�E ���H��G�?r�@m�?��	�ߢV�@�?�@�?��J��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�iS�?��?��/�Zʋ�=l��6>�^%?��Ӿ?h�>�x�Z�������u���#=W��>�8H?�V����O�d>��v
?�?�^�ک����ȿ-|v����>T�?���?`�m��A���@����>2��?�gY?coi>�g۾,`Z����>л@?�R?�>�9�c�'�w�?�޶?د�?\I>C��?c�s?h�>>x��W/��4��Ó���=��^;�k�>�c>����3hF�vٓ�i��R�j���~�a>4�$=��>�C��9��66�=Iۋ�:G����f���>A,q>�I>hQ�>�� ?9d�>��>	�=�l������3����K?�?���n�O��<yo�=��^�7?!04?��_���ϾP�>��\?���?�Z?�@�>A���:���㿿Uu��/�<��K>97�>7D�>����JK>��ԾDD��w�>Ϳ�>Ǩ���^ھ2H��"k��F�>�^!?~k�>�=?~l0?��>�>!������(�]k
?g�?�> ?+a�?�H?�̾_�K��飿y���o�;����=��?k�?/F>[ǆ�Kg��4 ��
��=!<.=���?��?�ˁ<j[	?��d?O�8?W�!?���}�n�Ο��~��Ѓ>c�!?��E�A�8;&�QA��r?e?���>j��8Eս�sڼ���c���=?5\?v�%?�2��h`��¾W��<rY�۵M��T<��B���>��>	���D �=�+>۰=��m��6�>Y<�=l9�>��=z�7����T=,?p�G�/܃�f�=��r�PxD��>KL>�����^?�j=���{�����x���	U�� �?���?@k�?�����h�p$=?��?�?V#�>�I��m~޾��+Sw��x��v���>���>��l���7������PF����Ž;��(��>��>�?C��>�W>���>����%����c���]�N��6�M�-�������Ns%��4�Ȅ����|�do�>V���*��>��?=e>�w�>��>o���u�>��_>f�>Ȃ�>/S>2�6>�O�=@�;�̽`_?8�m���N����J}���?a�?�.?ڐ��Gϔ�)��GU9?���?,�?�O>a~�\�K��G�>���>+"[��2�>[X.=��= P
>�撾~-��cY��L=��>W�e��EG�G�R�7��U��>��>u�
����E=Es��f,o=Q�?�)?��)��Q���o�u�W��S��D�TUh�^k���$���p��鏿{V���*���(�)=�*?,�?r�������1k��?���f>��>��>���>�bI>��	�}�1���]��B'������<�>rG{?u��>\uG?��X?A�H?j^^?Ǟ�>���>b�O�>'����H>��>$[-?)u>?��?�?@1?MF�=eS޽�����s�(?�<&?�?��>�;�>3���᜾�^,��O�V'Ѿ
�{�#}�>E�q>�_s������>� >���>�n\���ty���A>��?��>\��>dM��sc���]�gx�>��?���>�����%M���ܾ�?�$�?Y�D=5�1=�E�=Qj$>iK.��:ʽ�<:!���=�4a=����U݃=sm=�-�@��=�n�`5�=�>�� ?h$5?�D�>^�>��h�w�[��Y��=u�t>Q��>y��>�^#��I��S��EQf�E��=��?��? � >�=;A=~V���,����=©��o=P3?>�&?g�8?���?�FD?S�?i�=��)��H���JX̾+�$?�N?�*�>'A�3��4���&�E^�>ކ�>y�B�Z���X�5eW�;�����q��m��S3��篿��J��ѻ�a��r;��d�?�)�?庾#ܹ���V���K���(?�w6>�H�>$(�>��1���g���j���> ��>�d?�s�>2K?k�}?�TZ?��>>��1�.M���ݗ��u���0->�Y;?�
�?ۙ�?\�r?��>�,">3�<���龯��'9�f���s���<��_>�ɑ>�@�>���>3C�=!B��n��*n?���=��g>���>���>�^�>O�>��<�(C?�*?6ă�4(����s�վ�n?��?�%?��_=�վ.�Q�Ld��]�>c%�?�ݴ?՝ ?񏓽躦=��E<�JO�7���C�>�>,�>�[?=�2>мn>�h�>�>��X���.i1�� P��A?`
S?���>���[f�`���;Ѿ|(r<K�ٽ�oY���_�xt�yPE�{�
�T%�0�t�R�i�V!���X��zx�����S ����>��$>BO>�>�7=;����9>�s1>9��=0�'��#�<��=i�>��{< �X�u��2��*w=F:Ⱦ}E}?Z@H?<�)?'D?�|>bp>� ��.�>\��Nl?S�]>άI��
���K<�mU�����ڌ־�=Ӿ�.b�)����>�5��
>��3>���=�X<8�=��z=xk�=h唻��	=���=�X�=(��=^T�=�>\�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��>]��=�aK�p^1��L��sE�U�6�k#?��:�"Ͼ��o>J�=Ʌվ����v=��>�Pr=�y�B�L�0>�=l�U��xD= �z=3h>�<>��=�"��t�=1�I=���=o5j>��<���Hf���=uE�=r�d>GYN>���>�?&N/?��a?���>ܢy��b׾lž�yQ�>���=^̲>��=C�>>��>�9?lG?�NL?��>>s=��>Jy�>aj,���o���ᾛu��Br<��?�x�?N¸>&�<�D�g��?��/Ž��?)�3?�q	?6	�>�濞I��J��tzY��u��%2>�^(>�I̾J����H�|���Ǉ�����F�>g�?V��>�:�=�:�<��><��>�>>̀f=�f=�Q�=��@=R���5�>�a;�޼#l�Ʉ;P��<Đ\�}�^��*���tn:>��<;;Ͻ���=��>I�)>���>��/=�ç�ʍ!>O����K�G�=�䫾#JA���d�eJ����6�<� �Ũ2>YE>>�'�����4��>�Wr>�	7>2��?e�v?�>�=i��P׾�;���2G�\�%�c,�=0�> �%��9�x}\��M�B8˾c��>�<�>�&�>�'�>�K�<���"��G����-�#��>����`�н��^�����¶����k����#%?a�����cI�?yI4?�ώ?��?S/��D;����=I_��0->����܉�cWT�h"?1�?���>0��3K"�|����<�|>4����a�������u���.��/y?v���p�ɾ�C�������m�aC�c��t�>��?���?}���(��0�iU�*p��X�>A�G?�2�>�A
?�]
?��;X'��,����
>�%�?VW�?���?��g�l�K>��1�O�>U`?N�~?���?''�?�ū��|>'�E�@>$-��RV>�;?qI>*�����>���>��>��b�c�������۾'.���Җ=���;�>^x>Dl�>-;G>�:=#uǽ���pGc>j�d>pX�>��>�ś>��m����gdI?��>�Ë=�C?��g<[n=e��CA>�'��Wн�����}O��<�Q�>��2��Ƚx3��5�>�BĿ�?.�#=#���#?�������އo>�5�>3���0�>�wJ>uu>���>DMi>�=�E�>��>YGӾ:x>H���d!��*C�FR��Ѿ��z>����Q&�����r��8;I��k��>e�Aj��,��U9=����<�F�?m���Q�k��)�����ܒ?�Z�>�6?�֌����D�>5��>̍>�B��X����ƍ��i�/�?���?�;c>��>/�W?�?�1��3��uZ�&�u�[(A�e�B�`��፿����
����_?�x?4yA?�Q�<n:z>M��?��%�+ӏ�{)�>�/�';��?<={+�>�)����`�i�Ӿ��þ68��HF>��o?B%�?lY?xTV�sr\<�_`>�j+?Z�?�po?��+?��7?����"?�8>Mu�>��?f6?,�?=�>���=�>�G���I>cbq���v����#z�;i����ّ� n>��<ꮙ;L���3����=�Y����L<܅ļ�n8=uū�P7�=>�,X�>�І?UK?�z�=�VL?f✾�;�Uc��G�V?�ڇ>�N�ܿ�=�P���=��~�=�o?��?%�F?�w�>?�M������ C> �?N�g>�ܦ>r^(?lAL�F��C�e=F>p>8Z>�l >�)_;�Uξ6�&��&>���=T��>�,|>1�$�'>v���< z��d>�Q��ɺ� �S�J�G���1���v��F�>G�K?�?er�=b�dS��FJf��&)?�d<?fMM?��?rO�=��۾��9���J�A�? �>���<H��;���p!����:�]�:f�s>�%���m�kqA> B�h��YQg�3PD���վ��!>u�|?Q��� �&�;�HP��a�=f�>�`󾾍�ZE���Ԩ�>r<?�:m=�sk�ҶW�>|Ҿ��>�ȟ>���>4�׼i��^�L��h¾�n�<l^�>ם�=̄���Fݾm�F����	o�>J�C? �^?��?Rܩ���m�cI�88�gP����$�$)?�^>{��>R�W>�?�=���4D��U�(^U�ܭ�>�	?X[Q��9;��η=+�"�TdD�-��>R?��=��??��R?9ں>%-.?X�.?�L2?�%�>�_�vh2���?�N�?R�=k��<�|��N�]��R��{��>�p;?b���>a9P?	O	?��>���?´e?��z=�����d�B>J��>)?����`�=��%?���>�`-?��z? uA>B;���0��O ����=��>$�?�G`?�,?�'?`�?�1�����<�+	>+9?���?5y?��>t�?�A�=ݴh>N�<��'?ߣ�>��>��<?l�Z?l�?�9?�q�=w���J<P��=�"�c��<���ҏ�����<���~��ۦ�=�m<ӟ��lJ�_�]����������D=���>�xx>�d,3>�������	=>"���V���_4��f�=��>�b?�>~6��0�= �>Rǽ>%��MM%?Bp?X�?I�Y���`�rξ�nL��٪>�B?��=L<q�E����{r�|��=��k?��Z?�Z�y��<�b?�&^?����x=�>�¾�*b�|��P?_?L+F�˕�>��?$@q?j �>N:h���n�{�����a�d�g�!I�=п�>A���Id�֝>�k7?T��>j4_>�b�=��۾x����m�?�-�?�5�?0�?�7+>�m���߿�s���F���^?'��>�I����"?R����Ͼ5:��f ���+⾔*��,髾�$��1X��ʷ$������׽�y�=��?V!s?QBq?��_?ɵ ��d� ^�����qV���� �E�oE�3�C���n��d��O��Q���jG=$b7��6?��Q�?s�8?�(���4	?s��"�來k��ӫ�=�վ	�d��iI>�|=��t=m
�=�~Ⱦ{ƽ�������?��>ߝ�>�Bd?�!B��J��!Ǿ 7U�U�����=$H>�3�>�d�>�o���U�%*�P�%]��;=�Lv>�>c?^�K?�n?�K���0�R���4�!�N/�N茶��A>��
>���>n�W����&���>�G�r� �!���w�	�*π=Oy2?GZ�>O�>� �?�?7	��s��2�w��p1�l6�<�j�>Ei?�C�>��>�н&� ��@�>1 q?��>��Y>�1Z�^���ef����T��>��>r�?�(�>�C�d�e��a���i��v>9�@!�=hUp?�ą���n�Pf�>/`L?J�9��={ğ>,��H(����3s����=�\?�5>�0�>�+���$����a�T����(?eV?����n)��/�>>-?�� ?zŜ>�R�?x��>G̾
9��� ?x([?@�<?�s=?�Z�>�F�<��.�؟�Yq��9X=a�p>^�">�JX=���=W�,�,�T�K �#��;�m=}5���ޓ��a<��μ�\�<�e=9�>wп�hC�k�Ծ�*��,ݾ������| �x�����C=�����v���{��*�;��( =�����󛾑?x�\�8�&o�?���?LH���W��ҩ�T|��%�B`�>j�a��� =	$��%c��(���hyƾ�z�����4�)�{�Y��P�'?�����ǿ񰡿�:ܾ1! ?�A ?:�y?��8�"���8�� >NC�<�,����뾫����ο5�����^?���>��/��m��>䥂>�X>�Hq>����螾|1�<��?4�-?��>Ύr�.�ɿc����¤<���?/�@��C?��ZX��>���>���>U>T>��=�y>���(I�>Ē?6,�?�=FA�ic��;�W?���%�P�c��:���=K�7>e�r������6>���>ˢq��\��(��	�����>m�ͽ\0S�[o˾��Ѽȇo>�	�d�-�5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=�o��"���<V$����Mʔ=�	=�Am<�~�<*Ž��輨���K㚾��ֽ��
=�,->C>�OO>��l>��>��O?*f?泸>W!T>3 ��'��`�����s����$���R���I�k���⾂"¾�	�۸"�t�i��߮<�N��=�HR�?���,!��Gc��E�?�.?t#>��ɾ�&M��$<�̾�멾���gĤ��3̾\�0��'n��?%B?��hEV�LA�x�d���X?������ո�����=�6���=ޜ>���=~���U2�W�S�]M.?�t*?�k���¾�
_>3���N=�Y;?�&
?�}<�V�>0G?�B���#�n�`>
 �`�g>���>��>���,�&�:�%?"*N?B�ǽ�gR�}�a>��*����ӫ��棼E�������c�>�S#>�"�I,>#����O%=H�M?6<?� �w<��A9�AIH�������?h�,?��>.�?ӻ~?��:��3� �v���,��R9R?=I?��=,�1��~������AD?�^l?��>�=���f�$�]�Ⱦy		? �?�ň>�?=����|��H7�~*?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?r�;<��U��=�;?l\�> �O��>ƾ�z������3�q=�"�>���ev����R,�f�8?ݠ�?���>�������F>؟��}�?ₑ?�ʾ>1�<���x�����;g�<&�n;��4��"'=m�վ�3������T'��
��Q����>�@%�k�ue�>Τ<�3/翍ķ�ʆ�b����"�F�#?+ǣ>':�3���]�a(e�HpE�j�2�yf~��}�>zq/>�X���+��[2���$u���=��>rU���`>�돽N�Y�!�/�8lT>2΂>�m?ME>KF>Vy�O��?�����п�����!WZ?AfX?l�?�^�>����8i�<ۆ�@ >��S?J�8?~Bh?���N`j=� ��j?oR��Q`��4��AE�U>u"3?�I�>�-���|=`(>h��>\>�%/���Ŀ�ٶ�	���[��?��?�m����>F��?r+?`h��4���Y��C�*���<��7A?�1>�����!��$=������
?~0?e��+�Y�_?*�a�<�p���-���ƽ�ۡ>&�0��e\�oM�����Xe����@y����?J^�?f�?��� #�Z6%?�>a����8Ǿ��<���>�(�>*N>�H_���u>����:�i	>���?�~�?Mj?���������U>�}?�^�>$�?��=���>H��=氾�*��$>�}�=��?�}�?��M?��>�'�=��7�!Q/��+F��
R�Q����C���>��a?�xL?P'b>�d��R�0��;!�1Ͻ��1�(򼰼@���,��Bݽ�5>��=>��>�E���Ҿ��?Mp�9�ؿ j�� p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?[��D��t�o�z�>���?
�@�ծ?ji��	?���P��Sa~����7�l��=��7?�0�'�z>���>��=�nv�ݻ��V�s����>�B�?�{�?��>$�l?��o�Q�B���1=0M�>ʜk?�s?�Oo���b�B>��?������L��f?�
@u@a�^?+Y�ֿ�����;�˾���<�>yoN>�_9��Ϲ�(���V�'�4a�=v�=�">�j;�_�>d�Q>�r >;�C>���[�+����p���%�=��V��8�@�"�� Ҿ��1�����L酾M*�*��1��M%F�p�Q�1�����=�pT?+S?�o?'��>^�j�^�>������=�� �1x�=�C�>�52?<[L?P*?Qd�=E��z2e�����&��>a��%�>3�G>���>��>���>i�;�J>,�:>�"�>U� >#�1=w�L;��=�O>	�>�}�>m�>�N<> �>�δ�B.��1�h��w�&̽;�?����T�J�/���9��[����V�=0b.?Ja>:���=п����0H?����/#�g�+���>W�0?�bW?o�>+��6�T��(>a����j��Q>�) ��}l�M�)�<Q>�i?�$�>�g>P[-���^�e�Z�¾���>Y�??Z�'(���9u��Z��Aܾ�R�<�v�>��M�Y�������I���=aX?��>�}���8n�k҈�� ྙ�u>G��>(Oڽy1>�D�=���|�^�H��<	�S��=� >��?,')>0Jz=![�>�$��:�N��g�>�>M>�G#>�\=?�$?]z��х�=�����$�9�l>Ȉ�>S	y>L�>�nG��$�=��>z~d>����V��+:��D�$�R>�Ą��
f�+�x�3aj=������=x�=�&��4�D�\a=�~?���'䈿��e���lD?S+?a �=��F<��"�E ���H��G�?q�@m�?��	�ޢV�>�?�@�?��T��=}�>׫>�ξ�L��?��Ž4Ǣ�Ȕ	�6)#�gS�?��?��/�Yʋ�:l��6>�^%?��ӾXh�>&x�zZ�������u�m�#=Y��>�8H?`V��
�O�>�w
?�?�^�⩤���ȿ2|v����>U�?���?a�m�A���@����>1��?�gY?oi>�g۾M`Z�u��>��@?�R?<�>�9�R�'���?�޶?ί�?�I>O��?l�s?�j�>�2x��Y/�z6��o���}|=y2\;�d�>�X>����sgF��ד�Oh����j�C����a>$=��>�C佪4��r9�=I���f�ߥ�>M*q>U�I>�U�>�� ?.d�>���>e�=g��7ှ �����K?��?��E�m���<�ٛ=��^��j?X�3?0�`�THϾԨ>/�\?���?/[?��>����3���ֿ��e���5�<r"L>vv�>Kh�>��8�K>��Ծ7�D�wB�>���>V���81ھ�=���������>"q!?��>��=� ?$m$?3}j>L��>�oD�����F����>���>�'?k�?�?���m4�"��s�����Z�L�O>m0y?4�?���>�1��Ic��bk+���:����g��?��g?�M��?���?W~??��??�8`>ۚ�%B۾�Q����>�,"?K��{�A�_�#��D��|?U?��>�Ş����Fۼ����ѭ��?SS\?��"?���.a����sb�<�3J�=�;Z�<&$u��>�!>������=x�>~��=�3m���:�1'`<���=L��>���=a�;�����1=,?m�G�nۃ�X�=t�r�BxD�T�>JL>�����^?�k=���{�����x���U�� �?���?\k�?���'�h��$=?�?7	?d"�>�J�� ~޾��ZPw��}x�zw���>���>��l���E���י���F��8�Ž��½G��>9�!?�o'?.ܗ>"%�>�~ >�ĳ�G��~��+&�A�_��
�
�?�4o��0����x�P����E�~A����>��J��p�>CN?��=�7�>q��>l�޺���>��>���>X.�>�I�>}��>�C>� =�2 �XVR?aP��K�(����������??jrb?���>Ȏ��6�����B9?�\�?��?Lmz>ަh�Ј)�ۦ?)��>�z|�?�?��P=�	y�KІ<m�����L���I��S��>؟཰v9��	L�j��	?��?�aR��_Ѿ��ѽ�����q=^څ?a+?��*�v�P�A�n��Y�*�R�Cg�Q�k��砾}J"���n�j��֫�����>)���=�*?u
�?���5��	��Q$m���<��b>�;�>�>�{�>7�G>�
��71�_�\��&��\���|�>��y?��>W�U?�1?��?b�[?>�>la�>�� �>�<���>��>�5?s�C?�?�� ?<7A?��>��s={3߾��)�>m>'?�9?/�?� ?ƥ����ɾ��O>�6U=Ӳ���<[�d>}� �;X��:¨��j���[=nw?c�R�2�,'���g>��<?Y �>��>�wh��o�������>��?j6�>-]����a�0�g�>b
�?�-B�0�_='�9>���=�<�9ue��T�=A^Z����=ɷ7��x��菼��~= ��=�$��#X<a;>)�<y�r<�e?�#:?5��>~A>�OS�����Ē*>|>��>���>�j��%���������a�NVe>bR�?(м?PQ>ާ>��,>�X���[��� �%P���]�O� ?�R?� <?KL�?##i?�A?���6�!����bҍ� �Ͼ �?-�2?Uy�>���n{������[(�H��>��>ԍd������=�߽�A\����u&��o�����QP������`Խ$��?��?����7�
�6���:��s���7?�X�>��>�`�>M_���`��ᾜ�<�m�>�&?�G�>o(8?�ڄ?��P?K!>`��0��Ð���a;�2i>q�,?��W?���?�Vx?Ű�>nd9>@�E����n
���\���(�D'v��O=�D>�Ck>³�>ah�>�S�=h�l=���]�J��=�d�> x�>��>���>�W>Uɥ=�qG?c��>u7������������n^F���s?-8�?N�)?ȕ*=h���E�5��-�>��?�?��+?$.J�8��=9H������9�w��ϲ>���>��>[m�=Ma=OR$>j��>:�>H�|��f8��`��?)5G?<F�=75ʿ�������ܸ���|=j�\�h�}�<{��@���ս�޾
u��#���Ɓ�o*ؾ�)t�_������������>�7�=#2>m�#>�M,=:���*D�����rU,=k�=�f�=���=��<�S9;ڎ��}*>R��E��=��=3�˾�}?!<I?��+?��C?��y>-D>�3���>*���d@?]V>8�P�������;�����L����ؾmu׾~�c�˟�CI>�EI���>
93>�J�=cA�<V�={s=�=�fQ��=�*�=�H�=�^�=d��=��>�J>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�]d>c��=p1`�X��;"`�×���ic� �>?��H���־�w�>�!�=��� ��
]>�H�=�0=�Q���Y�R��=��ݽ���=1>GH�>�-H>3>����-�<��=��=� V>��<���D:��������>�(C=��+>���>
-?68?tD?J�>����O=b��Ⱦxץ;el�>P�?�h�B����?�C1?��)?�u?e�?&p>P��>Te�>"\��W�[�����ƾ���<>��?�t�?���>��5>�uĽ��7�W�v�J:"�J�>p�#?4�?��n>��P�Ͽ�_>�I�:�w��=��=��n�,qݾ��̽������о�Ǫ�ދҽc��=�.>_7�>�.�>mσ=�Nx>� �>�+d>/"=�YG=��=��3=��=iЌ<�
�=<:>�!�< �������a<<n�>��;�%,4<�N�=��=�=;��>hk>���>�=	���h/>ܼ��Y�L����=�b���(B�*d��H~�g/��]6��hB>��W>b���3����?oDZ>(�?>b��?ADu?��>�:��վ�L��W1e��GS�gø=�>q�<�is;�_[`���M��zҾy��>r�{>�2�>���>��Q��%��i���j.����>���&ѳ������q��m��l瑿��� v����>uE��8X��QI�?�I?�Ɛ?��?��H�O�꾭�>})�����= ���U�n?*���?��?Ν>c&��v�6�u<;�գ����>�i ��U�;c��#�����脱�Ɠ�>Ū��վF�j��-����k>�j;r�|��>F�9?���?�B���s��I;0��G-��PF����>im?�{�>�i�>�?�P;�%���&��{�=�?Ǘ�?��?H�����>�<ܽO!�>�d�>�d�?��?��?�\����>-O=�=��(�Q_�>B�><ش=IUO�|?wg�>2��>Ų����������*+e��	ż��9>�2�>��^>o�>bOn=?�u�v����B/>o�p>�r�=_&�=��>)�N>�����Q�)?�l�=؈>,�2?,�u>[�J=�졽��=��Y��fD���'������g���<G�~��?=k��E�>j�ƿ.6�?W�I>h2���?~<��E�+bY>�gO>A4н���>��I>�"�>��>�5�>&�>7t�>��&>�FӾ[>���d!��,C�_�R���Ѿ�}z>ќ���	&�П��w���BI�Nn��ng�vj�M.��3<=�uȽ<)H�?�����k�!�)�i���c�?�[�>�6?�ڌ�����>���>$ȍ>�J��^���Zȍ�
hᾛ�?6��?�;c>��>��W?J�?��1��3�-vZ�
�u�$(A��e��`�v፿ל����
�J����_?J�x?�xA?�B�<]9z>��?��%��ӏ�*�>�/�)';��F<=�+�>�*��.�`�3�Ӿ!�þ	6�qIF>��o?K%�?Y?�SV��w�L�,> A?�2?yh�?�S?�Ra?�m��##?B�K=l��>*��> o=?�$6?�	?g��=�C >u�d9�=�7������RP��($�C�_�=׺=�A�<����x�<��@=�8ȼW�a=��һ+�����==�;{�/@=iv�=��>Sl?P��>Z�:>b�?�m����0�-���m=?���?O�Z���d��N��Yx�>��s?���?`^h?�(�>�V�'6���K>��_>{b_>�g�>:t�>� P������Y>��9> I=	�>,6�=�Ƨ��x�-YG���=��}=+x�>3%{>�b��{	+>ޣ�p4{�cyc>�*L��ؼ��bT���F�t*1�b�s��)�>�<L?�d?2}�=.�꾺d��Y�e���'?A�<?\M?=?�U�=bھ#,:��qJ�����>K%�<��;��M��7;� �:ؿn>�㟾��!�v|2>W���2־�m�s�B�Iβ��>p>.i��d=�Y�_�ZF��B���� >��׾^�������[��-??�.>S~�Dy�1��ѓ����>#w�>�_�=֌��(K?�}Ҿ���LC�>A�*>N1>��ӾB�M�����>�IC?~�L?��?���3)g�h<n������8�� �e��A�>���;���>[�>�d=�B��B�M'^�UB9�}�>@��>��5��A�ۢ���5��z��C�>#�?¢ݼ��?�Q?�i�>��&?�C?�A?�\�>gH!<݌���4&?G��?U��=�ҽ�S�4�8��>F����>"D)?�C����>@?�z?x�&?�xQ?Ć?��>�� �6 @� u�>�Z�>]�W��G���`>�iJ?$��>�5Y?�ʃ?��=>`K5�#Q��A���	�=�>��2?]#?0�?��>IC�>|ߜ�Yk�=j��=&O?�?3�|?}�B�\�>�ꆽy>1A'��?�>ċ?�� ?�|r?4u?��D?I�	?뗮<v���?�:�����ɨ`�1p��@���b�J���T�*뼉�m�|��Y�����kZ|�Bɧ=�ˮ=�� �sMJ�J��>�w>V���N39>ǎϾzP��x�F>��j`��yK}��)��|�=�g>��>L�>M�+��p�=O?�>���>�2�o'?�4�>W/?����a�ͩϾ�R�X�>�B?Z�=�Eg�즕�{s��Ą=Bss?)�b?a~J����w�b?~^?)`�t!=�$�þ(�b�{����O?D�
?0�G����>��~?V�q?���>'Gf�:n�b��s3b���j����=[�>�M�&�d�t9�>l�7?�T�>��b>��=��۾B�w�ꀠ�c?T��?��?��?Ey*>-�n��-࿜Z��kH��"^?���>
a���	#?R��]�Ͼh+��8򎾝J⾟ ���ܫ��/��JV��A$��)��ؽ�8�=G�?�s?Z;q?o�_?� ���c�/^����j�V�������E�QE�5fC�9�n�t�R=��/���S�H=�X�o�F� �?*�!?3G����?�쪾����|����>������B'>���k�=��:>8�þ�����Ͼ�=?]�>�>�iQ?�n2��(��x,��xV�D^���=>Ac�>.>���>�&�=@�M�0ؽ����xK��|��Rׄ>�^?ɜ=?s�o?����.�	J��"}�{���������$>B|=��R>q"$�Jӽ�5"��P��|k�[e��������N_�^�?A\�>/݀>U��?��?����缾�[�R���k:�"R�>��w?]�>w۵>�m��@��*��>��z?�v�>\(>��T�����w��(��VM?��?)?I�>�o.���s�n��e���њ���>��x?�ۀ���{���d>c�F?��J<f^=�t�>葤�p�"�O��WP�s��=x�?�>M <>�;������c�"���-&?�.
?����-�)�>��#?���>�H�>��? �>�0ݾvJ��U?��_?�I?O�C?���>��=*�]�νν4�v�j=&�>NI>�/=�w�=��&���i�)d$���<#�=׿���9���?�<��m<}y�<=�h='$>��Ϳt�?����'��J�����B8��2�Mt_��M����U�Z�V����r��5d�=�̿���l�Q4��$�����?xv�?8k���m��y����������b��>����	>�C���=�ľqe����ӽI>&��tP��xq�@6n�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >^C�<-����뾭����ο@�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ǝr�1�ɿc���x¤<���?0�@�=B?H"%�����Y�=֟�>�7?1o3>[[��.\!��赾k��>��?��?H~�=�Q��M���\?*�=^�I�{9���-�=ا�="�g<|���H$[>h��>ɂ$�oI�V)����=u!w>M�3��{+�H�_�E�<�R>�4�J�A�-Մ?{\�vf���/��T��gU>��T?�*�>�9�=u�,?[7H�\}Ͽ�\��*a?�0�?���?$�(?ۿ��ؚ>u�ܾy�M?WD6?���>�d&��t�}��=�7�ǁ��O���&V����=A��>��>�,������O��P�����=� �Adſ��#���0~�;��L<Yφ�p��c�t��'ýHհ�v����E�۪<:ֶ=M=>�Ն>�m�>�G>'iZ?�ll?��>'x >�e)�M����Ͼs��r�� �ٽ8�X�,s��Q��[�誽�ʁ���n�Ѫ߾g6����=�S�� ����%��h� ?�h�-?�=>���^�B�ߚ?<U�Ҿu����V<y9�8�̾�d.��Dn��k�?�ME?���j�L����.ួ�����P?�%ܽ�s���6��OC�=37��=�2�>R��= �Ѿ��0��2S���,?x`0?�{����Ҿ�%i>��t�FL�:b+?Q�?�(���@>��?"=���U�ؤ>�C>�%�>;$?$J�>g�����T�Q�!?a1p?�������#݉>Z-�������m���W��q�$�=�ڳ>�\s>	�~���=kr�=Da�IGO?���>(:���(�oS�����2g�QW�?�� ?�@?4��?��@?�����{�F�U��g��_��=��_?�1M?4��=�28�~����:?%�\?̼>>g=���HG���㾊S�>ۤ�?��?F���qx��n�\+��}��>��v?�r^�_s�������V�s=�>�[�>���>u�9��k�>��>?�#��G��亿��Y4�Þ?}�@q��?��;<M ���=�;?�\�>��O��>ƾoz��e�����q=s!�>����{ev����gP,���8??��>�������[W>B��U��?JC�?ؽ����=�r)��Y��"���Fe>����i�#)�=���Ǆ9�4h˾87��V澤8�P�>�p@�Ē�6�?��u=���˳ǿ�mm�^����o�+;'?�~�=���e�m�v�>ߋ���=����!�2L�>��A>���� �=�Ւ�V[��k�A>�ܢ>�ȶ=_A�>���=ߜ�<�t\���"��[?�0?���>>�=׬��W��?)������|d����Wc?��u?�l�?ք�>I3P�`�=�}|��bX���U?�?�_?L�ǻ��=��߽`�j?�?��aM`���4��:E�R'U>�3?F�>8-��}=�#>
��>�_>< /���Ŀ�Զ�~���g��?��?k�F��>s~�?oz+?ge��4���N����*�:la��A?1>v����!��=�$�����
?F�0?g@�-�Y�_?&�a�L�p���-���ƽ�ۡ>��0��e\��M�����Xe���Ay����?I^�?i�?ܵ�� #�Z6%?�>g����8Ǿ_�<�>�(�>�)N>�G_�t�u>����:��h	>���?�~�?Lj?���� ��� V> �}?'�>��?��=�p�>܎�=c���67�g�#>���=܋@�A�?�M?�>���=�a8��
/��cF��?R�����C����>��a?�nL?�Ib>�?����0��!���ͽ�E1����n�?���*���޽ �4>O)>>yg>��D���Ҿ��?,p�,�ؿj���o'��54? ��>�?����t�/���;_?Cz�>7�,���%��^B�Z��?�G�?3�?��׾�Q̼#>3�>�I�>��Խu���������7>��B?���D��;�o���>���?	�@�ծ?ei�A	?]�K)��0P~��N�qU7����=��7?ՠﾬ|>a��>�ά=DMv�����bs�"m�>,�?�?�?��>�Vl?>co���B��<=-��>#k?�f?�[�J3�8�=>	I?O���Ў�qQ��pf?�
@k@{�^?ݶ���5ܿҫ��V׾BwܾC2��l}=IK�>:�s��=gA��u=�F�E[=�=�>���=�=�U>w]>1�x>D�c:(�_�������(,�_��rt���`��gQS����:����Ѱ��2��2'�R�`�J���?f���<h�'>v�H?t�(?H�r?�6+?�s����2
���0� V�����=��>�=?WOM?U�,?EZ�=/��)IO�/M�Py��B_�
[�>��>��>ǟ�>�>Pg�+��=o��=>��>0J�>��=>�>�w��lz>�l?2��>���>�<>�j>�ʴ�R(����h���v�z�˽[�?z���ܱJ�Q'��熍������=	Q.?ZC>D���/п���$H?Aɔ�>��	,�x>��0?4eW?��>�ڰ��U��>�1	�2�j�N>e3 ��l�V�)�o�P>A?q��>|.c>��5�Q�;��]����⬚>��T?��Ⱦ�a���k�2Fo��@�	^-=m��>���<C*��$��K��i�O�=��P?���>���־*�K������Mt>��>А�;0�>-<T>'��=��"����_dB�e߱���=W<?Ж%>S@a=�R�>G��>�Q��K�>�2W>XS>��;?�&?�m!����I9��,��n>g�>��>�q�=��E�2v�=7�>I�S>�G��gb�1�%�A���S>�*v���m������_=�������=~ψ=4� �B&G��=?=�~?�|���ሿ#��D��erD?�2?`�=`�G<�"�$���R�� �?J�@�k�?�	�S�V���?�?�?� ��>��=Qh�>Zʫ>�!ξ��L��?�ƽJˢ�4�	��/#��P�?��?��/��ċ�&
l��'>]%?e�Ӿ�h�>@u�@Z�������u��#=���>�8H?T��ݴO��>�w
?�?�_������ȿO{v����>H�?T��?M�m�*A���@�-��>Ӣ�?�gY?qoi>�h۾JfZ�ǈ�>�@?wR?d�>�8���'�/�?�޶?m��?J>�f�?� s?�a�>k�iS/��]�������y=q^�:��>[�="A���uE�f%���G��^k�C��S�_>��$=X��>g:�h��}��="<���M��]�T���>/�m>��J>R��>@`�>7��>|��>1�=������U`���K?���?����&n��w�<:k�=�^�N(?�C4?k]�^�Ͼ�Ψ>��\?s��?B[?�\�>���<���俿|�����<��K>�*�>�I�>$8���MK>X�Ծ22D�gk�>`ח>�e���5ھ2"��^���G�>�g!?[��>��=� ?��#?܏j>�ѱ>�BE�@+���E����>V��>!u?��~?�?�͹��r3����}㡿|[�T>N>|	y?)E?i��>����x����B�sH�����/��?�_g?���Y?l)�?Sx??ՇA?#�e>G���ؾi���ẁ>��"?���FB��#�Z	��Y?L9?�S�>U?սRD��㼭|���D�?�{X?�M"?�t�9OX�xľ��=Ņ��g�;�N��P�0�&>>��>6���x��=^4>�F=��|��1Q�ܱ�)t�=�*�>2��=�xT�����=,?��G�=ヾ��=�r�vxD�e�>Y]L>����^?V=�u�{����9v���U�b �?��?~k�?�#��^�h�"=?��?^?�$�>�F�� �޾��ྂYw�C�x�v���>1��>E�l�v�V���?����E���ƽ�����q�>Ϸ?�8?���>�-|>Yux>�˞���vѾ;�
�
vG�+�PO��N8�x#�\�Ѿ�t��P���žOn��߸�>�|׽��>�	?td>uo�> ?�>7=�n~>��=���>ô�>���>yT�>�s$>N!=��ý�DQ?�N¾4�(�ef侂����@?9c?��>����k���j�@�?�?�<�?\	t>��g��(���?v'�>�wu��T?ǳ-=u0�����pʯ�ކ�|��v^��~�>���6�
BM�h!w���?T?#�ּ�GϾ���r����i�=.q�?�3?	�#�ٖK��x��wb�۲S��V���n��`̾���VoW�r��R����ڈ��{.��խ<��'?M�?@��Q|��|���r�'D�o��>"�>;'w>�Y�>��>���D](���R���(�A���/��>W�x?���> �:?��.?�K?�/I?JPX>۴�>���J�>��W��-+>L@�>� F?Ċ&?�l?�t?,�-?�D�>�2�<��澇FԾi�?wf?�"�><�?Q�?mՁ�D�3�Hh<�p�;:���98=��7=��归w����>G�x<�0�=B�?G���5�(��΅s>��???�>�>�>~8�����e
��]��>��?x3�>l'㾾�d�c��{�>���?�?���=`>��=iǱ�6ك�=����%=L*�����n�<w�=�~P=��<�N�<U�6=��%=K�0=6v?�F?��>��K��5:��u�.m>����<�Y�>�f�>�WH>1Ш�U3��요�&�q���s>ᨓ?q�?�̋>��=�E>⛾G����޾T<z�[��<��>,?)Te?�?*�7?��?�Zɽk��㓑�^񈿵q��u�3?=J1?�d�>?���Ï��,�����5�[��>p�>�CW��x���.�%ws�0�J��=�8S�H��N��ɺ���O���>%�Z������?���?��ؽ<���"�Xܵ��Ƣ��0?.R�>�n.?��>����p�bv&�ǂ+��c�>�L?Z��>��L?3-h?��`?��>@=��Y��t2���䯽�9�=��=?���?���?��z?ǂ�>ͩN>c V�'�Z����z�� �u���f�=�Э=�ʔ>w?H�s>�E%<�=�*9���=G>��5>�)�>̾�> �?F�`>��=,�D?m��>"-ɾ?>	�\ꮾ�ٝ�� ��.d?J�?�]7?�R=b���Q�7������>J;�?R��?��+?/�6��> ��}¾#L��I��>���>/>�,�=g��=~<>5��>�~�>�3"����]=�t8.�l&?]C?��
>�Zǿ�(u�H�q�������<ͤ��v�^�����#Y�l�=�����)���ą]��E��凙��Z��	
��3vk�v��>Ẑ=���=���=�S�<ʌ��E�<�=X=d��<ǧ�<�N��(�<�+��-�<��8�);��!<�/^==I���]˾��}?�0I?ژ+?��C?h�y>��>ύ2����>4��n0?3�U>w�Q��d��d�:������5����ؾ�t׾2�c������`>1�I��>U�2>� �=8�<�;�=��r=%T�=J!1�~�=�x�=ظ�=���=(6�=1�>l>�6w?X�������4Q��Z罤�:?�8�>i{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?Ati��d�>M���㎽�q�=N����=2>s��=v�2�T��>��J>���K��A����4�?��@��??�ዿТϿ4a/>���>��<��m��������U�_�`|m?�k]�o�\� ?\�ڼT�[��퀾LU$=�e�<HB��!;��r��N�=��սO>A�r�p>�>.k�=e���0=��=�|9���=F5��,��(O��c�k=������g>_�>q('?"� ?{==?���>Ӆ��������*e>�\�:,�>�_`>�cl>��>�}?�9M?2{a?�j�>�A>́�>+�?]Q�/~��Xk�	���ﰾJ�O?�@�?�k?�w;�����C���F��n$���>v�?c+?�?C#�9'鿢�"�ӕE��p�",�=�	>��B�ٚ_�c٩=� .�`/��PP=g&4> �R>�«��u>��
>�G�>	��>�/a>Qw�=���=�}�<X��:�"��;�d�z=��f=@#����= V3<}ʵ����=��=:3�<4�h<�c��b��=���>%9>o��>b��=`���D/>����?�L����=9A��,*B��0d��D~�j/�O6�#�B>�DX>?����2����?�Y>3l?>Ȅ�?�Au?Y�>��M�վBP���@e��VS���='�>F=�U{;�Y`�i�M�ʁҾ&��>ɢ>I�>1�~>Q�?��D'�!�9P7�	@:��X�>k|����P=��>�Uw��<Ϫ��Q��kSr��(��A?�b����F=�߅? 7?�%�?��?V�l��Θ���O>{�?�P=�� �l(��E�b?�?��>V�����̾]C��6H�>J�G�vP��&���0��#�It��N�>�e��r1Ͼ=^3��D��*D����B� ir��S�> �N?#��?�;_��a���N�j6��>����?K�f?���>֦?��?���0�Z��ht�=�Lo?:��?_��?n�	>$��=����,b?��>*�?�}�?�M�?�1����>$"߽����j�ޘ>r�x>v=D5�=�?]9�>jO?8�����,���e���Z/����=Ҡ�>�7�>��v>�>Δ=�)�=��>�*_>%K\>��*>p��;���=¡=������T<?��=A+>�V2?NJ>��R=㽟��+�=���(�6��߽i������2~=�ĭ�.����۽���>��¿��?DcN>�2���?2��*ދ�n�>1aj>"��C�>2�w>'��>�>���>�Ӭ=o�>]5!>�"Ӿ2t>����L!��EC�wR���Ѿ��y>�����&�{���^��xtI�z������$
j�X1���S=�7�<�1�?����p�k���)������?�?�>46?�ٌ�D���K�>���>U��>�x��]���
Ǎ�Q]�$�?I��?4Cc>R�>��W?��?�v1�e3�~zZ��u��%A��e�v�`�a⍿d���C�
� ���ƽ_? �x?MrA? �<,5z>���?��%��я��1�>�/��;�f�<=;/�>�4���`���Ӿ$�þ�B�{vF>��o?�%�??X?�WV�'����E
>G�U?�{!?��v?��`?"�W?H~!�e�?`b�<��>?l�>f*?�?y?(k�<��X>�V���MQ=R�Vsn��,ͽ����{%�
��</�w��E����=L2<��>������u��=�PL>�nٽ�G�$y	>��S>B��>]�\?�R?�>��3?&B��vN �������7?ר=�,ƾ���?;:�g�þ}6�=?k?Iz�?�H}?
��>��[�:����>z��>��5>"�>�?�>r�G�]��}�>�||>ID�=\��=��������[X��U�S���=���>%&|>�N����'>�w��<z��d>0�Q�tܺ�T�8�G���1��\v��e�>��K?�?���=�E龹o���=f��#)?>]<?3HM?��?�1�=��۾��9�r�J�l?���> "�<D�����k!���:�b��:I�s>�8���8Cb>���uz޾A�n�J�E�羡]M=�l�-�V=N�_!־]�R�=��	>:����� �����٪�o?J?�Yl=4n��vYU�Zq���>Ǉ�>�ۮ>4�9��v��@�x���@��=q��>I�:>о���bG�m<�_��>�)<?j�m?�}�?�A����h��QG���g�;fR����?'ض>=(?S�>pv#>夾����g�&�+�$��>�
	?]P��[N�H/y������/�K�r>z�?��,=�8?5�B?��?�4_?�"?1�?m�>삽�\���'?�7�?��U=n�i�a�&���0�ҾH��ֱ>i-?9Ӕ���@>�i?ڵ?#�?`�M?	�?Y�$>�r��\�����>�w�>n�U�7n��kY�=��B?+6�>�Y_?h�?q��>nA�����C�2\�=�5�:�~2?�%?�B�>$5�>���>�O��oӝ=@��>fj?��{?��e?��=5��>�w�=�^�>��>�>Є�>�N?�O?�yl?��E?���>��<C���i�޽Iݙ�ﲐ�^����l<���=�6l�"�:���缉+=�ר;;FO�-)3������⋽��+��xv<& �>�n>{*s��=yqȾ�5޾��4>i�X=�W������n%~��/�<�k�>;q�>��j>�iN�t��=�?�G�>��?�*?;/$?*�?{��=�A��?}��P��>�>p�9?�I�=l�f�� ���r���&>[�o?dz?z�㤹���b?n�]?f�[=�r�þ��b�X����O?��
?H�G���>3�~?f�q?0��>�e�1:n�7���Cb���j��Ƕ=`o�>�W���d�zC�>��7?�M�>��b>��=_s۾�w��p���?6�?��?��?	&*>��n��3�ȡ��N��f�]?�(�>� ��s#?����b�Ͼ�I��L���%��[���`��Y���|���A$���2�׽���=q?�s?�Qq?��_?S� ��d��E^����jKV����0��E���D�JZC�-�n��N�����-��=�C=a\�,YI���?�?]`�1�?��X���Ѿ�Z�W�>!�����U'��i��Y>p>�1����.�sm��f�?gի>"/�>��m?X�Q���F�vE���O�bt�yջv��>ι�>X&?2��=�#�P���ݾʾ�k��^�v>�c?
[K?��n?Y���H�0����$�!�ٺ0�>�����B>��>�P�>^'W�V"�me&��>�1�r�R��c���H
���z=2?�Ń>�Ȟ>��??`�	��O���gu��0� �<�u�>ki?_l�>]�>�(ս�,!�g��>p�l?��>��>u����`!�Ƒ{���ɽ�.�>�ǭ>\\�>��o>Z�,�s\��N���~���9����=ѐh?̲��a���>B�Q?���:�$N<6��>vx���!����H^'�*\>i?8��=��;>��ž�A�*�{�e��d)?"d?�撾�\*��}>��!?=��>F"�>�3�?�қ>b�þ�W�Pa?�B^?��I?J[A?�v�>Nc=����Bǽ%�'�&�*=�.�>Y>�o=�?�=�v��Q\����I=��=��ϼ���D�;]|����E<6��<`1>��ֿ; P���t�,þR���Q���q��pK��k��O��pҷ��J���ޖ��`�:$Z���]�{k���;��r��?���?��l�+C��Ӈ�#������>ha��A��=�ݾyș�C�'�m#�������.G3���A�P�{��'?M�����ǿ(�����ܾ �?�' ?��y?q���w"�%�8�%� >�q�<齞����+�����οi����^?Ӹ�>n(�Z���	�>�W�>XX>��q> ����/����<��?j�-?VV�>~�q��ɿٔ��=��<ռ�?��@|iA?�&�E��R�(=9��>�7?��<>gP#�+������=��>���?K��?�1D=-�W��$���e?쨩<��E�y��� �=��=X�$=����C>_�>�%�<FJ��S�	�6>�m�>\�4�����+_�ߨ,<j&Y>�Wνg[��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�󉤻{���&V�}��=[��>c�>,������O��I��U��=����ȿ`'��&$�==��1=:ڼ�&ѽF?���7����~�s�׼�#m�;�!�=�E>�wm><C&>:A@>��V?��k?O~�>��>�����݅Ҿ����3d��Y������J�����Vm���Z����y�y.ܾYa,��B$>4�N����t�޾�Wi�qk�j�?9�>y�W���V�g�澖�V=6R�˔���l2�Mk�� ����[Į?(�s?�Q��_��L*���a&���C?P��=��ܾ����m;xg�>��3>��>�8<4�~�>[@��j/��M>?j?ƥ�?&��<��#�'�9>�"?%-?~��=R�D>���>����T�`g>��>">�>f�=><0>� ������?��H?P<�ۻ�q�>*��fƃ���L=�>�� �$p�}|F>�+�=�Ҿ�͚��E�=[���UkU?��>�`7��$1��־u�۽��=�χ?� 
?�I�>�>0?�UC?��=(��w�V�]��
�>��n?UY?a� >�m��!���#Pq�v�?>A?]%�>�)��
���<���Ծ'-?-�X?�3?�H���p��%v��Q��I�A?��v?nr^�;s�����N�V�<�>�[�>���>:�9�kl�>5�>?�#�eG��ú��CY4��?o�@u��?$�;<�#�z��=	<?�[�>��O�#=ƾ|v��������q=�"�>닧��dv����+Q,���8?���?ē�>I���A���>�G�����?���?IPȾ k=���w@g��(�.>=��>��9�O��M���������*]!���̾���c�x>��@���D�?a�"��Xڿ�Qտ� ����־���?��>һ=|����A���k��51���M���5��P�>#Đ>u��W|���}��s<�u�Z�^o
?�z>,��>���-����=��ܽЧ<@u�>��>$">���K?���o��;���l4��=??���?�z�?�I�>��>��ʾ;]-=��n�s?�y?ț4?��"��۟��d>�g?YU����b���=�@[��G�=5!*?��	?ua"�t�0=�U�<*J�>C�S>W��6ÿ����9Ͼ�2�?��?�����>�8�?�=?B �%���P��3����� 1?O��>����8��Ϋ�� ��Ά�>:�?E"���]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?���>��?�b
>�>���=ॾ�ض=��=L��=������>`vI?h��>"@�=�W��p3�!�L�NRP�&�����G��4A>��S?me:?%4�>y��<!���k(��P�N-	����<�����C�~��`>�>B߄=����5B߾��?Jp�9�ؿj��.p'��54?,��>�?��}�t�����;_?Sz�>�6� ,���%���B�a��?�G�?>�?��׾dR̼�>6�>�I�>*�Խ����`�����7>/�B?I��D��q�o�y�>���?	�@�ծ?ei��	?��ON���^~�܁��7����=�7?=-���z>���>@��=umv�8���0�s�Ĵ�>�B�?N{�?���>��l??�o���B���1=K�>5�k?[t?L�m� �m�B>��?�������K�� f?�
@�s@��^?�좿��߿�����о��׾Ɛ�=��)>�hd>)�½)��<�yp=�n=�ε��=�"�>�]�>���>��*>h6�=R�=
���� �����<d����D�����
�}؊��� �~
X�ݞ徭���-f;;�/�����¸��Y9�KQ���P]���>��9?��@?d�k?�@?(��=A��>.e
���!�M�ν�;>�ܕ>' ?��>?��8?��J��%��6l���s��P�����>�>2B>��
?�I?(�o>��"�!x>�y�=<'�>�p>�	����=��f=�8">6H�>���>�B�>�C<>��>Fϴ��1��k�h��
w�r̽1�?���R�J��1���9��Ӧ���h�=Gb.?|>���?пf����2H?'���y)��+���>}�0?�cW?!�>!��t�T�4:>6����j�4`>�+ �l���)��%Q>wl?��f>a%u>[�3�bZ8���P�_s��	s|>S26?Pʶ�)9���u��H�^ݾ�L>S��>�A��a�C���x ��ri�
<{=�r:?�?�B��$㰾�}u�q:���@R>LA\>N�=�i�=�TM>��c���ƽ�H��9.=	��=pi^>ڇ?7�N>T��=�p�>54��H���
n�>��>1Lh>��6??s)���h��ˊ��>��&`>Z�>Xhi>+�>4e����<#� ?�MY> �/���&<Vw����%���$>�҈�����u�����Ǿ?�gz<>�E^<�,�14��>��~?���(䈿��#e���lD?S+?p �=%�F<��"�E ���H��G�?r�@m�?��	�ޢV�B�?�@�?��E��=}�>׫>�ξ�L��?��Ž9Ǣ�ɔ	�()#�iS�?��?��/�Zʋ�>l�}6>�^%?��Ӿ���>����c���)���v�K3!=_f�>�sH?C����6M�#�?��s
?�?"e�#�����ȿuv�{�>(��?Lޔ?��m�������?����>�e�?E�Y?�Mj>�۾TC[�f��>��@?��Q?ԛ�>g,�	)���?Wʶ?ną?OI>���?��s?/n�>�+x��Y/�=6������&J=-dY;�g�>�\>����AdF�Y֓�tg��,�j�����a>ژ$=��>�K�|6��>�=�����J��I�f��>
&q>�I>�U�>�� ?�`�>֥�>��=;h��g߀����y�K?���?���2n��Q�<䠜=s�^��&?rI4?h[�O�Ͼ�ը>˺\?]?�[?�c�>W��O>��5迿M~��t��<*�K>4�>�H�>#��rFK>��Ծ�4D�^p�>З>4����?ھ�,���K��1B�>�e!?u��>�Ѯ=ș ?��#?��j>*(�>�`E��9���E���>���>�G?��~?��?-Թ�-Z3�=��q桿��[��=N>t�x?/V?Wʕ>�����)�E��GI�V���
��?jtg?�R�t?�1�?_�??��A?6*f>&��Zؾ]�����>n�#?�޽R�:�<��(�/�?��?��>)＄�Ži_������ʣ�>bDN?6�"??W ��c�����L=4�Q��4��W�7;	�?��>}�G>/._�k��=kVL>~��=ܐd���4��o��Z=៑>'d�=��7���� ,?�5A�ʑ�����=˥r�ǕD�{�>�iN>�{��z�^?�;>�/�{��ି�I��q�T�I��?T��?�~�?烵��h��|<?.�?��?��>哭�n|ݾx�߾Jw�kw�E���m>e&�>z�e�o��G<���s��p;��N�Ž6����V�>j3�>m?)�>;;0>i�>2׎�._Ѿ����N��>���.����L)�T�����!�5��x�־�ʔ� |�>���G��>�/!?h>�^D>٭�>r�<N��>L�S>ԷB>S��>]n�>�*>��=��e�(��~'R?;�{-(�<C�~ ���P>?Z6c?a-�>�Oq��݄����yz?t��?я�?]4l>��j��7)�l�?�U�>y"���	?�"V=oO;���<�3��L&�� ����A����>�����!:�VMK�(�b��7
?��?��׼
�ξ��佭���\�n=UJ�?P�(?��)���Q���o���W��S��y�H7h�Ct��Q�$���p��\��#��١(���)=8�*?"�?*�����  ��*k�7 ?��_f>�	�>�$�>�ξ>P[I>%�	�Ĵ1��^��J'�����Y�>'R{?��>��=?s9?A[?ƴP?��>���>Иھ�_�>ʢ0�>Ѻ>�	?�?a�3?o�?��$?P#(?�_>N�.��&��:�����>t��>��"?!t�>n?�忽��]X$�k�=Qv��7�ʽ��=�f=�k=�+�:=�\�=�S?m����4�/�~8�>�=?��>:ټ>׾��
���ɕ=Z	�>���>�J�>4S��9r�a=��H�>�}?�P��<��>!��=�2��ar��,��=bԥ�S�y=��O���4�������=+�Y=1L���:!ɼs�;t�=�� ?2%?<�y>b�s>����P��0��:�=��e>��]>)��=��Ӿ�l���d��W�g�e�j>Ȧ�?{�?'I=�h�=�=���X���ֺ����R=c+	?��?�L?���?��B?%�?�>!���㔿�򃿶,���?��,?ϳ�>K��)۾�l��.>�I�?�k?�Y�̵��2�_���)�A�Z�=>7����+��n�"�k�~���]r���-�?ȸ�?�˜�!U2�J/�~�����Ѿz<?F��>�/�>���>B���z]���4%�=��>d�??G�>�#P?���?;XZ?Z�j>Z��(���WĞ�8 ϽƆi� 7?�xQ?�|?[X�?�S�>0[�>t����U��c��YX�r�V��J��vd=���>��>z��>�W>�T+>y��f�ӽ�l,���=�x0>�^/>�S�>v%?jO�>wrE;��G?wx�>�־,���ؽ��2���y����t?���?@�(?3�������1����r��>\��?P�?�;$?�,1�2B	>q���"���f�$��>Q�>�,�>�F>��:d6>s��>D��>�,H�JI�c3�����r?�d8?�=?�ͿS%��!����)���5=���g�F�b���K��=�f�3��߭��Ql�� {�Ͻ���Ⱦ�
��6�c����>&�=�K >���=������nm<V�=��=�<4��`��G�U�;J�K�ҽ1.a=�=�(�;o�n�ھʾ��|?��H?׮+?SGD?�|>1�>��9�?ԕ>qށ�ea?n�V>d1T�7���Y�8�$S���p���Iپ��׾�xd�88��9y>nH���>��4>���=n�<i��=!�m=��=�/L��p=���=ǹ=�D�=��=�p>,�>�6w?U�������4Q��Z罡�:?�8�>�{�=��ƾu@?��>>�2������xb��-?���?�T�?@�?Eti��d�>^��5㎽�q�=d���>>2>���=��2�H��>��J>����J������4�?��@��??�ዿТϿ,a/>�f8>`v>�{R�!1�k\��b�h�Y�ww!?��:�B;̾�V�>込=�6߾D�ƾ�-=ڊ7>�c=�/� �[���=�|���:=A�l=^T�>��B>I��=.S���۵=�DL=w�=�O>@���c�>�,�*��r1=���=2�b>�{$>���>��?�b$?�\?cv�>$���߀�����Q�=X�����>[֩>�fp=/F�>��0?g�8?��?ız>.�>��>(��>- 6��u�!i���?x�8!���H?lq�?|��>�V�������¾�4����k��>^�-?{�>���>'��o��<�=�N��݃;�4�>^��>;;�]� �=c��=zfy�}z��Fa>>�>ȱh>·=�Н=T�7>5=�>5�>�E�=�i�<O�n=r��<O���}�="�Z=;T8<hА��YW����=�%��z{��v����m:�&)��f=lj>Z��>?-$>���>Az=Z����X>�[��[�B���=Is����:�n�^�2x�/t$�� L��M2>ضS>-�b�����Lw�>"am>߼)>��?�b{? X->"�#���ھ����̿@�n�8�}�=~>���8�f8c�}(P��о��>�֍>e�a>�^>tK9��PN���=}V���[G�״�>����n9����!;�f7�u板�祿�Y��>EH?�u��2ل=�?�?Q�Q?���?�.�>�n��*��o�P=�HԽ�i>�b�]~s�Zg?���7?/R?@+�>�-��,7��F̾,������>�nI���O�i����0��{����ܝ�>T����о�3��e������B��'r�>�>͔O?��?��a��L���IO�d�������_?�xg?$�>BB?+?���}Y�=�����=��n?���?;�?w>1��=�Aདྷ��>?�?�a�?�ؒ?LKu?�a�{�>t
0���>"����#��K>�=>-�>=x��>=��>��>�k���������8�C�J�ع�;Ű�=�ĝ>��\>7#U>hy>E�*�!K�<9�%>^�>�>�	>�p�>���>�h��W?	�P(6?4� =��7>�\7?o�>�4=>R��*�>��<!j`�ᴾ8�&�d6�<���=��;:��=K�����>(=ǿ��?��W>��Q!Q?��ξ*l,���=n��>���"�><��=�O>���>���>����������= 4Ҿj�>�Y��!���C��rR�־Ѿ��}>OK����#�:�	�j��[�G�ҵ������i�療���;��{�<0�?�� �/�j�ti)�wG���?Ǡ�>1x6?��w����>�v�>�b�>ec���S������I9����?���?��d>���>Z�[?�n?N�#���,��^�'y�m�?��ih��X��f��m@z������ ��S�c?ʃt?9{7?2q=(ys>؝~?p'�����3�>K�(�xm9�%�<�#�>�q��Cm��iھt���ӂ�l>[�o?�~�?�:?3�X����Fi�=H�&?��<?��?�(D?�]=?\�\�c��>I5=tA?6;?VB ?�;?,A?'o�=�Ƽ�r�N�n� ���⏾f4/��ǽG�h�!�j<^�.=�ށ=8��S���Ř�={_g����ܪ���v�@��W����7>S�>�B�>�X]?I�
?�?�>Dl5?,��j*N�����l?�'*������׎�s��AN�=eO�?�9�?�#;?�C�>�W�B����B<�>
�>>��Y>���>vBv�4o5�~=�<�E>?�>l��Ҽ�����ܧ��2]�A3�=��9=���>�x|>���z�'>3n��	z��d>k�Q�������S���G�:�1�bv��6�>.�K?)�?��=�v龪���s3f�>)?�<<?,M?;?�Ք=�۾��9��J�Ʒ���>�r�<k������5����:�H1�:$Ss>R���Π��qb>���V]޾��n�
	J�����L={��?V=����վz&�b��=7
>V���� ����Ҫ�,J?��j=�y��u�U�Q�����>*��>y�>�+:���v���@�䝬�w��=���>�:>���D��7uG��1�|�>�O=?
�_?��?'A�h�^���;��V�%�ľhp��I�(?T��>}��>�ߋ>Uj>��x�����g�݊>�AW�>#�>��r�N�"�ƾڪ��\�s>�?��>���>�3??I�?�5H?�
?���>2�f>�	�8F��ڊ&?y?3��=���������)��$ �:�>�5?�x��B�>L '?��(?��?VB??�>�y��6�	��>��H>ӎn�����(�=��I?	��>��f?�jp?��<�M�Z�T���=�;@�C<=�T??��>E�?+��>,����-�=���>�c?N&�?3�o?�C�=E�?B�1>���>ܖ=i��>���>�?iPO?y�s?)�J?̕�>q��<1E��VD��G�s���O���;3I<z=�]���s�z0�)�<Ӳ�;�ⷼ�́�0y�c�D��t��F��;�M�>F�z>+j�����=2r¾��о��={�$>��p���7�t`�Ӵ�=�?=ض�>)i>x�b�`=���>W@�>,F8��I?�?K�?�dS>��4�n1��5׏�%�>�_?}�>*H��N@����n���@>�K`?"p?2I�&��I�b?x�]?�g�=�*�þx�b���r�O?u�
?+�G���>a�~?8�q?(��>E�e��9n�����Cb��j�Sζ=�q�>_W�2�d��?�>˛7?O�>��b>$�=s۾��w�xq��I?��?��?��?�**>G�n��3�&�L7��d�T?�6�>�����* ?�*��Ծ݆��t��оF��nা덒�����������#YԽ�2�=��?U1�?��s?Cr\?{U ���k���i��\����L���꾷���I��MG��FG�Sj�b��Y�޾�p���B={�G��Q���?��5?�┾�?���DǾl举X�>��ξ�%t����<Q`#��[�>
�=5zھa"J��:��^?gT�>�� ?�%V?�s��'���H��&_��<��n�=�ֈ>s��>�?aE7>C����=�@��U�澾* �J�v>�Rc?�fK?��n?����0��,��
�!���2��j���D>��>|O�>I�V��I�&��>���r�~��^f���	�)�=\2?V؀>��>��?��?�m	�`z����w�z1�v`�<��>c�h?��>JX�>s]ҽ/!�9��>�l?Z��>��>혌��Y!���{�$�ʽ�(�>�ݭ>���>��o>{�,�K"\��j������A9�K{�=��h?m�����`��>�R?/,�:4�G<�|�>��v�M�!���򾴽'���>�y?��=O�;>�}ž�$�;�{��9���T)?IL?�꒾j�*�?�}>�"?
��>�)�>(�?��>{þgg���?Դ^?\5J?�AA?��>��=W!���Ƚ��&��+=�U�>��Z>�zn=9�=����x\�H�F�C=+_�=��̼ ���
<%��6�K<}��<4>�jӿ�D8��BξG��{�����&0��&|-���k��h�<;oh�!ܾ��{�,����N��	>��[x�ܼh�Ѹ�?U#@��:��FY�(T���M���d+�2�>�'����=�.��劂��^���u �����B�J:�0�7�\\���'?����ںǿg����9ܾi ?�B ?<�y?��S�"�:�8��� >GT�<6p��9��斚��ο����E�^?���>t�NV��|��>��>Q�X>i_q>����㞾w�<��?�-?Ң�>��r�ܓɿ�����<���?�@}�A?�'��{�i�R=�&�>lR	?��B>�/�>l��p����>w%�?��?K�6=��V�����c?�cP;>E�{�ƻ�3�=ש�=̴=��4�M>�Ŕ>���H�A���ؽ�1>�"�>"���ͷ_��j�<g8]>Fnӽ�Ώ�5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=�����ο�>�;�D�K��=6�4>X�=/c�)`D��Z��X����[���V_��kU�:
=Q�>-��>W�2>�G?m�T?k��>7J�=��&�Rա�$�־ֈf=�C^�`<�����~XU�DFe�@E�����.�(�σ9�ɏ��r��<�8�R��=kL�῏�����Gf�0FI�n� ?��/>C�����@��7��%>ƾ�3���w���Hg�������%�W�p�s�?�<F?�C����R�Fh�F{����ǽC�\?k§�H��� ξ�n�=7�=Z�<෠>�d=���X6�NY�"�;?_�?�澥���/Wk�2��U-@�Q�U?�?��'�3�D>�{<?hߔ�Cl��V�.���v>Q0V>�?�B�=�Y��,�-�"wB?�:k?�HC=~�Ͼ���>�E��u���>E,�>�k��� � �9>:�*>����ͽ��н��rW?뚏>��*��H�%���h%�1=E[y??4͚>��f?�9D?��<T���;T�_`	�}t{=��V?��h?�
>�؋�Ǘξ�䥾��4?-Xd?^�P>�]�Տ�?�.��� �6?��j?��?]ȼ0�x��Ւ����?7?V�v?:j^�m��*����V��'�>�O�>N��>��9��>��>?K#��K��<����Q4�gÞ?��@<��?m�:<k��{o�=�;?�f�>��O�Z&ƾ���|���q=x&�>`���7fv����$v,��8?;��?~��>\���ʢ�>z����?4�?J�� _>�c��Bh����&��=���<�՗<aq�=�E���r������%��dо��Խ�9X>]@������>����n�׿y�ؿ��z���O���U2?�[U>�@L���ʼ�����rV����MA����>(��>����wp�/��#d_�k(3���>�%�>s��>{J����G O��0�$��=M�R>+?��V>�c%�d�?��Ҿ�)ɿӇ��f�4�؍8?�Ku?Ś�?1�R?L������mze>J��$�-?��?�?6�U��=�)�=��j?����_�u�2�5�E��=Z>�f4?=��>��*��Ef=��>��>��>n�.��.ĿƉ��`���j@�?_[�?O�׳�>���?$[-?���ؙ����%�+���;�@?M�6>�����B#��[:�Ԃ��.�
?�i/?@q��l�]�_?+�a�M�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>e����8Ǿ��<���>�(�>*N>lH_���u>����:�
i	>���?�~�?Qj?���� ����U>	�}?<��>g�p?��=�?b=�Yo���O>�Zm=��~>ido�A��>��C?cG�>�BS=3.7�o�7�bl6��oM�L��m:�9�u>Hh?;�7?�7�>�k���_R���6��,=�;�a���=�I*�M� �;���>�>�=�D�=(��J�
���?�i�ƖؿCk��#�'��/4?���>?���,�t��i�q>_?p�>N2�-���"��4����?�C�?��?�׾��˼?>1�>E�>�ս�ǟ�!�����7>>�B?P
�G����o�
�>E �?��@Ӯ?��h��	?��O���_~� ��Q7���=��7?�+�m�z>��>���=�qv�����s����>XA�?J{�?x��>��l?�o���B���1=�S�>�k?u?.1p����1�B>׵?������M��f?��
@eu@��^?�뢿�lѿ�����b̾&Y׾�Z>�>�U>�.Ͻ�=��j=#=��绿�>��>;�.>�MA>��5>�H->��A>E��I�$��c���P���=�+������M�}R���{��#	��Ŧ�=kƾ��
�n��(`½�,�ċ��p�J�)<H>�=?�<@?�ib?g?��=�L�>��EKʽm���>���>%�+?-ZZ?��?ϔ�@�þ�AX��֌�!���7�x����>�N�=@|??-�>��6>w@{���U���o>�s�>��"�z��=��=>#=�?�=�qh>���>1<�>!F<>��>�δ�w1���h�t	w�w̽� �?�����J��1���6��~����[�=�a.?�|>����>п	���I2H?Y����)���+���>��0?2dW?ʞ>E��!�T�6>����j�uY>�- ��l�Í)�#%Q>�l?��f>�u>�3��U8���P��g���|>�#6?�Ӷ��)9���u���H�Yݾ�9M>�þ>��G��i�$���l�	�i�L�{=�y:?_{?��Ұ��u��N����Q>VN\>��=�_�=[WM>m�b�7�ƽ�8H��8.=��=8�^>Z�?�s.>J�=�t�>�:��'1W����>%�H>�3>8??v�!?L-L��fǽ+<��H�$�V/|>b��>pc�>��=kX�T	�=L>�>@ d>�à�h]D�����D1E��Y>� ���R��b����k=����O�>y)�=�ٽ��D��=�<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�m�>�e��Y������u�>�#=*��>�8H?�E��XP�H >��y
?�?<g�]���+�ȿ�uv�\��>��?��?#�m�h@���@��|�>���?-fY?Հi>c`۾iZ�册>��@?�R?q�>�;�C�'���?;ܶ?C��?�?I>u�?Djs?���>1m�zV/��񳿦u��`-v=z��:)��>/->(���d�E��g��2��0Cj�(��ZZa>$=���>��>���@d�=LȊ��ϧ��e�a�>@r>#/I>^��>l� ?��>���>L`=�����ܥ��r�K?���?����n���<��=�^��	?Y?4?��X�	�Ͼ��>��\?���?��Z?x�>����:���鿿|�����<��K>&�> ^�>Ј�$K>��Ծ<�D�gz�>�ߗ>���oھ����_ߞ���>oS!?:��>ނ�=�� ?#?�zj>!�>�eE��8��w�E�w��>β�>�C?>�~?��?�ι��X3�����䡿,�[�HIN>�x?}V?���>ˍ������E�<I��������?�pg?"���?�2�?~??ϣA?�f>Pi��ؾa������>�"?X)��/A���%���[�?�s?�z�>r��Ki⽂x缦���(��Zm?�}[?��%? ����a�Cx��-��<��@��e����T;4<��B >1�>M:��8Q�=|1>�Ч=�k���1���;�4�=F�>�=�y6�ꅈ���&?�Dr���w�&Ĥ=ىh�vC���>��f>h۴�l�_?�8�P�~�JW��Y��L�>�Ѳ�?"��?�a�?���Y\d�Z1?j�?*�?���>�y����ӾO ߾Ay��v����̮>���>{���ξ�N����xh���L��c��a`�>"�>�?�\?��K>�!�>3��4'����'��2�\�(�#"6���+�9��*���$��������Xo{�g��>������>��
?�g>�}x>�5�>E0عo3�>̡R>4Ӏ>jܥ>��R>�2>�k�=e�;��hTS?�÷��}&��ھ8����A?+�h?Kg�>�%�秃��
�$�? �?��?�FN>I)i��Q)��$?z�>�Ђ���?��}=��=���<0r���l�4$⽫������>چ���h7��LS�&�T�{/
?�?���z�վts�՜���o=�F�?��(?�)���Q���o���W��	S��w���g�����~�$�v�p�7쏿{V�����(� @*=�*?�(�?�~�#�&���4k��-?��Bf>c�>M?�>Fپ>�"I>3�	���1��]��='�+����^�>�E{?��>�5I?�$:?glR?�&P?�|>Q�>b����C�>St�nr�>W��>Q�.?F�.?��3?�h?u�&?��^>��ʽϣ���Ծ�x?�9?G�?�?�� ?�w�X��mY�����m�K�%�/h=ߴ��pս�Q��>�<}�">S04?o]��P�,�}%�g��<\�D?�?2�>-a�	�Ͼ)��Y?��T?���������h�����H>��?9;��~���j�=pa?>n}��u��=x}>-3F�l@>Ju>\�Ƚ���%�<��> �I�g�#�tF6=u�>�Rp�>�?A��>�@�>�;���� �-��؏�=!Y>'S>�>SKپ�~��$��	�g��_y>+y�?�z�?�f=��=.n�=Eu���K�����`뽾'�<%�?�F#?�ST?Z��?��=?i#?u�>�$�_L��r^��$����?��,?~�>�&��˾fᨿ��5�n ?�R?{`^�i)�}�(������N轗�>0�ɪz�cc��\Z?���㻢���������?	�?7��7����3�����Q�D?8�>纞>���>�I)��b��G��	9>A �>�.O?�>��;?���?Y�h?�y>���,V���g��� ���p��(@?G�+?7:X?��?���>�>���CF���ֽ���P=���C ѽ���>%/5=+�>�j>��/>*,�� z���^ս�_�����p�>d��>�K�>���>��>�mD?A�>.d׾�6���Ǿ0ٔ�(�ֽY"�?h��?�j ?��e��P�?�P���߾�<�>2'�?��?��>?kJ����=�I������
��h��>d�>���>X�>˵f<�O�=��>F�>�/���9�d�.�0�=�V�>$�9?;�*>z@ӿ/���n�޾L�׾R(g>������J���<U�h��z!������N�{3��`�6��(ξP��äƾ�쮾���#�>Uv=�s�=&��=1�=���hg:6��<`�d=�>H������c�<��=��<|#�={�F=Wht��;�/�þf�{?�G?�~,?��F?m&e>b�>��c�p׆>E���D�?	�V>.�h����)�)����h��8DܾIؾ��^�	�����>n$��ש�=�1>=5�=]<��>%��=�fw=��P<Q�J=y�=eܟ=��=D��=X�=U�=�6w?X�������4Q��Z罥�:?�8�>h{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>N���㎽�q�=L����=2>s��=w�2�T��>��J>���K��A����4�?��@��??�ዿТϿ6a/>K�8>5h>�^R�$1���[��Hb��X�	R!?��:��C;߅>'v�=ءݾ�mǾ��1=Q�6>az^=b��x3[�Mj�=X�}�N�4=�=c=Z_�>8�E>���=���@�=�M=2�=�O>�lI�2C�*_2��#2=���=^a>�	&>��>��?}]8?k�d?�`�>�>��q��e@�T)>ĈE�2ȿ>�2�=ܷ%>f<�>Q�(?ݏ[?��J?��{>�Q<>2�>AV�>��/��\�����a>f�z?uJn?ͅ�>"Ԍ=�ӽ��%�pH�_�r�m?� -?9l?;�|>W(�(���}D���'�_b=EC	=��#> i����Ľ�	���B<,J��)T�=�̝>	Vt>�>3IO>#�=4��>tx�>r�=�G����=݁�=]��=�9�����=f����w<a��Y��;y6>=>/߼�C<��=sR-����Dy>�=��= ��>M>�d�>(�=�J����.>5��A�L�Px�=�;���EB�8dd�H&~���.�f5�cUC>"?Y>���3���?�UZ>��?>�u�?�Ou?|� >tF�JVվ����d�[:T��{�=1�>O(<��R;��_�)�M��0Ҿ1�>1"�>5Ƞ>��g>�9,�&�@���h=�ھ�3����>n�����O�Q�n�?p���L��}�h�C <B?K~��	�=b?��I?�M�?��>!����ھ�P)>Mv�c=�w��yu�	���*�?��&?/��>U�뾄*D��Ѿ�!�����>P5]���E��[��DA3�ū,����!��>擾�Dﾢ�2�j�����|�8�H}P�L�>WE?�߯?;���<|���H��#��������>Y�c?�>x�
?B��>NL�C�޾�C��\��=Kh?H*�?%��?��=�6�=�)���2�>�;	?x��?�m�?�-s?	�?�̚�>u�Q;��!>�/�����=��>�Ҟ=6��=�[?]
?��
?�M����	�(��'�񾅰]�� =0��=qq�>uH�>��r>)w�=�i=}�=�+[>xO�>��>��c>�/�>K��>*֞�m���7)?!�>/�>\'6?`b�>7�->K���>�伽=@T�����m�[�ju�=�h+;�t=�=�=�[Լ� �>�Fȿ���?Xt�>�$�"�E?�@���� �9�=�X>��@���?��>��Z>GQ�>$�>ʣ�pP�=��>ϨѾI�>a���.!���B���Q�{]о��z> ��$*)�	��n���,E������EPi������=�a��<�	�?u��E�k��*��]����?���>�
6?�V��|���e�>�I�>Ya�>����qj��"���Iy���?¤�?�Mb>�h�>��W?�J?x�0�7�3�Q�Z�Žu�A�@�lXd��"`�P�������j
�����$�_?��x?,A?�.�<�v{>À?��%�L���@��>6r/�3;��Y>=�?�>☰�M}a��Ӿ�\þ~=��G>tUo?�1�?��?��W�ɌS���->��9?�=2? fu?k.?��9?6���?��)>5�?�{?OS2?��/?e�?�(>W��=�F0��=_�� <���ѽhwֽ���g�<=q=�z�:�Y<�:;=��<Jh�^�����5;��\��< �!={��=u�=s�>y�I?AX�>5��>��E??⧾���r&�����>0������h��nt�ݙ˾���>��f?���?;<I?3�>�I��퀾*A�=���>�6>q�>t��>^
����(��=P�5>2O�=���=�̽��K��F�-����o!�=x��=��>$*|>�:����&>K����{�Ac>`"O��2����Q�6�G�v2��ry����> �K?�$?˴�=ݓ��!����f���(?5\<?u"M?��?~{�=��ھ�9�vJ�J���>Hǈ<���l���-���::��ߢ;��s>����P��Cga>����޾Mrn�d�I�s���RN=�O�0�W=n��վ�~��I�=v
>/g��3� ����ﰪ�G-J?[�l=5���c�U�f˺���>=k�>���>��:��0s��P@��P��"��=2��>5)<>�>��G��G�J�R6�>�]F?�s?���?�莾�R���KW�F ��m��j�)�t�??��~>�h?eſ>�?D>�&���羞�M���F��T�>-R?�R��@8�ǖu�7����B�w�>>DJ?�6��>�W{?nL?k�8?=?���>y�7>i��<�Gn�wb+?d��?d�>J��<�o�O1K���:��"�>��?fLྀ�O>$�6?;sC?ӎ?��I?vk?�1>;�ž��S\�>$��>�&h����A2>��g?rT?�KJ?gT?a�f=�cU���齡�C<�6=���r?�N?P�?ɹ>��>F���;'sY>�Ed?��?�t?��>��"?o2U>	�?�,:�h�<[�>�a�>�N8?2�u?#�J?I?	�=8���V��\ｌ�n��>�#�<�΃=���I��_���+���t̼q���[��=���&��<ǃ˼�=���>�>h{���O>�ľ�nZ�k�n> �����gݕ�Nw^���=�2�>�>�>!n�>QO\��	�=^ �>GR�>�����$?�P?�s?A&I=�-`�Qh��K��^�>"�M?�{�=qTj�WD����o�I�w=�Fh?+�P?B_a��3�O�b?�]?�g�=�3�þ�b�����O?��
?��G���>��~?��q?'��>�e�K:n�����Cb�f�j��ж=<r�>X�	�d��?�>s�7?-O�>��b>%�=Zt۾��w��q��?X�?��?���?~**>S�n�34�hK���a���]?���>8��L#?�*���Ͼ���؎��⾟ȫ��嫾To��>�����#�D��ؽ��=!�?C�r?�Sq?�_?h� �5�c�F^�n��{&V�G
���\�E�Y8E��oC���n�������☾i�J=�=�&x@�wp�?�o.?��|�\,? \���aӾ�H;��r>�U߾�>��QrL=&���f�=�W�=���.^ �X���?�ϖ>Z{?��j?�`��53���P��t]�8$����=�^�>��X>��?[��=�&�r�-���ﾲnܾ����}�v>'[c?v�K?� o?�� ��n1��:��`X!�X�;��ʨ��F><J>�Ή>j�U�n��s>&��W=�dDr�&��/��E�	���v=��2?e��>���>�!�?�?����ܬ��w�א1���<���>�Eh?`.�>�ԅ>��ս�!�Ҳ�>��l?���>k��>�P���}!��{���ʽi�>�u�>RA�>��n>i,�n�[�D>���t���8�j��= �h?9d����`�Y��>0R?oة:k?<[w�>��u�Oq!����k�'�k�>͓?�\�=�0;>�ižj8�գ{�#���ͫ'?iv	?�H���f$�(܊>��#?�-�>E��>q��?S��>q̿��^<�?��[?�%J?�E? ^�>��ѻg���Dν�K7�n�<�z~>��T>��s=���=;����Y�0���X=j��=D���Zf���LQ:��ɼ�u<��<U2>Eۿ�L�oݾ��M��F	�Q.��@D��4냾�\�����o��z�q�q��/� �Q�P�״i�����*i�r8�?� �?�;���
�����5�����R��>�s���U�G量�����(߾D ��/O���i�ue�)�'?;�����ǿ찡��9ܾ�  ?mA ?Ҧy?����"��8�v� >�4�<�>�����l��� �ο�����^?���>�	�)��i��>"��>ҟX>�Eq><���瞾�0�<��?a�-?���>̍r���ɿD���l��<w��?��@h�A?m�"���辭-H=���>p	?�PE>{�/��`��緾\4�>�ß?�F�?��\=��U�E�/�
�c?��{<�A��ϔ�/c�=�A�=�4�<�X���h>�q�>��+��{D��-Ƚg�*><r�>���*�f�a�`m�;�oR>��ƽ�Q��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=x6����{���&V�}��=[��>c�>,������O��I��U��=Y����Ϳ�8]��@�>d�=S�f=zT>.���R�:�A=����b��ס	�,7�<�i����->B���

��Ml>��.?UZ>?�"�>a�(=r�H�^����ݾ!F�=��2��o ��ͽ��<��~��}�.�����"����u�.���@��1%=��R�y:������i�B�7�?+?/i�=�H���<���̽~)��r����(�`S<��ھ����UL�S`�?C?+^}���?��!��%��� ��Y?�	ҽ�Ӿѱ����9>��>칅=�D�>/�[>�{���]'��@d��A0?��?1+��������)>/2��/�=��*?_u?�O\<	ĩ>3$%?�S+��彦\>�J2>4��>�a�>ks>0Ǯ���ܽ)~?��S?�2��q��>�ý���y���h=eb>�5��0��ȴY>	�<ݍ��H�D��̏���<�XS?��>�� ������[�Dt=3��=�bq?C� ?M�h>͆Y?�"C?0��<�X�
O�.���}>��Y?q�l?7�>]D���޾�H��-�"?�Sy?�ъ>rޙ���=�������?"�W?�?���Et�J)��������&?P�v??V^�li�������V��7�>�L�>��>��9�Y~�>�u>?f�"�N������ag4�6��?�@��?C�><Q��Ȏ=V@?J-�>�sO��ƾ ���M�����p=�
�>�O���av�:��ɥ+��p8?���?�_�>v�������.>e<�����?�w�?�̾���=��!��Mn�b��B�<��`=@d�H�<`j���~�7������ھ)a��&�>��@iݽ��>�����R:ѿH��0����x���	E?F�>������xpZ�v�U�;W���U��a��^��>욅>Qj8�X����ي��yd���J?�̩�	m�>������=� $y�ֹ>?��y>|��=��⾪�?:�ΆV���4���9���T?�%�?5ݏ?�@?&?>|�b�m�L�x��'?�Q`? <?�K�=����[�߾j?�_��iU`�َ4�]GE��U>S#3?�C�>�-�_�|=�>^��>%e>�#/�p�ĿHٶ�������?���?8o�6��>?��?6s+?�i��7���[��?�*�Z(��<A?�2>g���;�!��/=��ђ�ּ
?d~0?�y��-�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?Ե�� #�g6%?�>d����8Ǿ��<���>�(�>*N>cH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?� �>��?��>?~�>���=
���3�=�*�=�N�=��E�K�>�I?C�>6ј=Z�����6�PnA�q�?��
�+A<�_ �>e�f?-D?�>��,��9)��J��{н�F����Q<�=�������<7>I�I>!>ߌ8��"����?�o���ؿEh���P'�64?���>:�?^��4�t�5��
5_?<g�>�6��+���#���3����?�E�?L�?��׾S̼	>�ޭ>�=�>9'ս�矽k|����7>��B?�'��B����o��>���?s�@Ԯ?A�h�g	?���P���`~����7����=�7?�0�,�z>{��>C�=nv�߻����s�c��>�A�?�z�?���>}�l?�o���B���1=<J�>��k?�r?�|m�0�h�B>n�?������*L��f?��
@Yu@z�^?��տ�ꟿڔ����n�3>&I;>N^�>����۽�y=t��;ΜȽ��)>o�<>��>���>���>��>�ܼ=�8���$�$r�������5U�!��])���g�F/�!s���{3���{� @&�͑�D'D<T�þ����:��U.>��S?W�K?߾i?~��>7H�x_o>Q���.¼sz
��� <���>��(?9?8/?|��;qF��*�N�|�d[���(���{�>Nz/>���>���>���>�)�<�6N>q!v>��>6> T������<柀>���>���>���>�Y;>:�>%ϴ��9����h���v��̽��?:G����J�h��A���k�����=�q.?�l>����@пDޭ�#(H?����8���+���> �0?:W?�7>c���)�Q���>����j�:� >W�����l��)�t�P>�Y?��e>_it>��3�ɉ8���P�Y_��/|>46?`����E8��xu���H��Eݾ�FM>��>&F�d�������~��4i�f|=dt:?-�?g���ϰ�6�u������"R>�\>��=�t�=�L>�<f�\Ƚ�>H���,=}s�=��^> *?�[F>.T�=�>xׁ���h��/�>r�1>�>��3?,�*?K�)���	�}�l��AQP>�>�>4�w>W�>Q�@��}�=[��>[�t>ø�Ĕ��
_�IL,��i>�!� �N�[_�kM�=t��D�=lE�=W�	�ɃF����<�~?���(䈿��e���lD?S+?] �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��J��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�j�>�j��X��x����u���#=���>�6H?U����O�z>��y
?/?C[򾜨����ȿ{xv����>��?d��?W�m�%A��@��}�>]��?ViY?�_i>$h۾XWZ�3��>ֺ@?�R?��>�9�f�'�#�?�ݶ?���?��I>�8�?�_s?�V�>��m��P0�lY���㋿�Vf=_�:��>��=����E��䒿���D�h����e�b>M%=�E�>��佲˸�Mr�=\�������h�#۸>Yu>� F>]
�>�X?К�>�>M={q������`��&�K?���?�U���l��N�<��=C�Y�o�?:�3?�m�$�оh�>�\?i�?�'[?,0�>���0���#���f��HZ�<(�N>��>-4�>�5���VL>�HԾ�bC�|��>3f�>�(���۾�����Ǆ��|�>:� ?��>�N�=� ?�#?��j>�(�>
aE��9����E�4��>ߡ�>�G?�~?�?tҹ��Y3�U���桿��[�`<N>o�x?�U?!ʕ>H���ʃ��O�E��.I��ɛ�?�sg?�P�!?2�?��?? �A?�'f>c���ؾv���s�>t�!?-��A��%��Q��?,]?I��>뎑�ءֽ�BѼ�(�����Ʈ?K�[?B�&?���[�a��Y¾��<��D�m���o��;�I��>z�>��؁�="�>`�=(gl���6�MUm<2��=�ӑ>���=�6��G����:?�P�="[����b�_���]OL�(��={��>2����g?��ľY�n��p�����������Г?���?Bv�?-6z���V��Y?4��?�'?z|?�y������3F)�/[���z8�6E���[޻5z�>2��>%z�����'���p��Ll�e����>%1�>{�?;3 ?�>G>�Ȳ>7#��(�}�쾋��_S\��k��o5���+����,�Y!����$�þ�X|��ۗ>�
���>�C
?$�f>J!x>�=�>b���7�>u�Q>>�=�>�P>G&<>�	>�2�;�BƽjcT?�C{��s��f���;ľ�GL?>�g?�B�>9���Z���j��*?�1�?>͌?jw�>P!���[��K?�(�>����R?��=WS=���=����
�3��hv<ל�>���z.H���L�0`Y��q?�G?���%s۾�dv�����un=_=�?��(?��)�u�Q���o���W�S�]<��h�)���{�$�Q�p���e���.����(�&�+=��*?f�?�~�Yn�z-��J&k�,?��df>���>��>��>i,I>k�	�?�1�4�]�(@'�ᣃ��[�>UD{?�b�>��??h�=?r�U?	R?�t>Q��>�h���$�>�'8=hQ~>eY�>e�-?�j?�h=?�?�>�?K��=���B���		��ӿ>�V�>x�.?��?Qlq>>\X���Ҽ�O��Jy<�E�l�̼&�>ޅ����!>ݧ/=@��K��=(%?���ғ��о�%4>K�V?ٟ?�1�>o
��p�Ҿ�����#?UF"?��C>�?�43��������?u�t?����0��S=�K>�������=�2>o�,��Rg=CQF���=�F/�)��=�3<��=���[j�����;�lC:�u�>��?�a�>��>�	��� ����ັ=�HZ>�MS>�f>�پǀ�������g�xpy>.{�?u�?��h=�C�=b�=�Q���O��c�� ��<��?E#?�HT?!��?�=?%<#?��>,��8���K��Wآ�p�?f�/?R�>��������t���R:�GX�>�;?�Ie��]���;-�D�Ѿ+;�k`>��&��k�v��� �>�%����T��Fɽ�N�? ��?7�=��'���Ѿ����M���U,?��>\�>mB?�\��VS���"�J��=�9�>�0B?�U�>�/_?���?�n?�=AG�2�ɿ��ą��Z5Ӿ�6?��?i_�?p>�?K��>.W�>��<O���͜��䦍��ǽz���8ؼ�6,>��>�P�>��2>L��p�m�Ww��qͽ�*}��7D>���>�w�>�{�>���>�7�>�sL?�x�>�ݾ����8!�^���
��?��?Q85?��G�8dK�޹6�5��>��?���?��N?�ã��=>�j�@-�6l��1�>S�>Dݓ>}��=�l>�f)>M��>�s�>���������K�wZ<��??�?��=�3��h+s���
��62�)��=�F�;2�,�/�B>�=�J ?���î����s�����_\���j�"=�r>���>���>OT�>,��=���=�,Ǽ_aν������<�:��>�������
�.Jq�h)�XM��P�A>x��=*/���}?�I?�.?_A?��_>$�0>�z�����>�[]�	n?DQQ>��(�.<������د�ר��i�Ͼ
bҾDd�'���r�>[��.�#>�>>�k�=�O�<��=�A�=rܘ=+x���+=���=b<�=���=���=���=�R>�6w?<������� 5Q�,n罱�:?6�>䑭=�{ƾ�@?��>>.2�� ���Lb� +?K��?�T�?��?�xi��c�>����Ԏ�hv�=&����;2>s��=��2�}��>��J>��� K��P���M5�?�@Q�??D⋿��Ͽ�^/>�7>�L>(�R��1�x�[�F�a���Y�!?��:���˾�h�>m��=T߾rZƾ4|0=z�6>]�`=�t��
\��̙=ц{��D:=�k=�؉>W�C>3y�=���<�=�AK===�=FgO>g���*:�8�/��c0=��=c>�V&>1��>#]?i <?��S?�.�>�t���Z˾���	m�=���K�>�x�=8t
=Xo�>�|"?�:?�??|��>[�=�hX>�6>X�@�^�A���z���\�1c�>?؅?�$?���=����U<��1m���$��>6ME?��>̴>U����Fc&���.��w���Ĳ6`+=�_r��OU��B�����A��88�=Kx�>M��>��>/+y>`�9>׵N>��>_�>��<�.�=pc��tǵ<�h����=ᑼB��<�ļ���)� �b�+�Ƭ���;��;9@Z<_��;��=���>�>�O�>���=̗���->������L�[��=9����1B��qd��\}���.��k5�7*A>�W>"؈��1��H�?7_\>EKA>���?�u?Vt >��8׾z7���6c��bR�$��=n�	>�;���;�Nt`���M��PҾ��>�6�>�)�>-�l>�[+���>�l|m=��7���>�Č�$b������n��Ԥ�#��a�h�1��*�A?䁈�V�=�f}?�vH?0��?�X�>�#����ؾR�3>PS���:=�d�Zo�sa����?�%'?�)�>m��r�B�v�Ծ�Ƽ�8>=��}�?��3���p'��P���K۾���>^�+��+�.�+������y���A�.��_q�>��K?�ް?J��=��N�+o̾fW%���ؾ�J�>sR�?���=�f}>��>�Y����m��K���7�>T�?�@�?�J�?}����C>����>O>2�>�b�?7�?I_?6��<.y�>�O=27�>���=�S�����= ��x��=i� ?�	>��>SoN�����L9��`ܾ$^�&m�<�
>��?j&�>Ô>�p>��ϼS]��{�<)��=��<�v>Z%	?l��>���,����*?_ژ=�m}>�h5?І>$�>4�,�bJ�=P��1V����1t���O�O��=��>m�>�ؼ=o�>��̿���?[��>Bf ���&?A�)�ɽ�<�=M�>>o|�՞�>���>�Ƅ>�)�>7=>%S=>:�">5��;{ԾR�>�8�!��|B��Q��+Ѿ�Nx>�z��1="��n�ؑ��C�I�����^�i��{���V=�L��<N�?�A��Q�j�!�)��M��uJ?��>^\5?�������v�>��>���>�=��lC������������?B��?�!c>k=�>�W?R�?��1���3��nZ�h�u��9A���d�E�`��썿������
�0ÿ�/�_?��x?
kA?9�<��z>���?��%�L����Ί>Y=/�");�F5@=�>r&��d=a��uӾ�Cþ|��T�F>��o?�0�?c?w�V�j�2��?->��9?o2?��s?��.?��<?��#�8�?�U3>.n?w�
?r62?)?��?o�/>�K�=�ö�=�����9��$�н��̽z�i�VM=�'O=�b<2�;N�=×�<4���st���<���~��<hMc=�=���=R��>.o\?��>�؈>8"5?�"��q2�a���v*?m�2=��g�$��ȧ�����:>�2g?U��?#'Y?,fj>��@�9J�b�>K�>��!>N�]>�E�>�8ԽgT8��L�=�>L	>�g�=�ሽi�x�d��r��y�<��>���>���>���;�2>,ݩ�y��;>u�0��
���$-@�qi(�9���N� ?7�7?�!?��ם�ǒ[�?�r�*!?�<C?p�C?�ؒ?<)>�����A��}B���R�1a�>��=�vʾO㜿�����'��1Q=�z>O�y�=Ϡ�� c>S��U�޾3Zn�G#J����8K=�%HY=���e�վ��~��l�=�	>������ ��񖿕����JJ?�o=^X��
V�^>��]�>��>�Ԯ>�:5��lq���@�tp��y�=���>�;>!���5fG�m���>%@?y]?<��?��"�WIh� 0C��L�����z��km?���>r��>l� >��8>xV5����-sx��N���>C�?�H�9JT�	"ʾ��� �0�4#�>6 ?�l=�J�>xpL?�$?�09?��>K�>䊨>c�8���J+?VX�?�<�=�.�{�`�+�K��3�C�>!�.?죾7F�=�f.?��&?�n?�1?5�>�>�{ྶ�fl�>$�>��s� ���9�=�jI?o?�HV?&�k?��j>�oO��L4�0�,>��=���=^�{>�F ?3�/?��D=��>�,羑@��5�>��x?��?��{?-C�>c��>��]>�m?񳍽��8>�`�>�?�A?��J?z�1?�4�>^��<���Sa�2ǋ�ZO��u+��Fm=0]T>��i��3���䋽/��<X��<�,�f۽q�/�0T=���=�/�>�Y�>S΀�)T�=�s����"�=��>>�t ��k���(�U�;g(T>���>a4�>*;��?>�g�>fq�>D�L�&z	?H,?��#?Ϡ>�X�:F��?��?�$>?+a?KM>�+������R�B�Va�~?vR?�n����9�b?s�]?�U�=�$�þ�b�_k���O?*�
?��G���>#�~?��q? ��>T f��:n����Bb��k���=�j�>�O���d�jD�>��7?VB�>�b>W��=Mt۾�w��r��,?H�?Y��?x��?�*>�n��/���� H�� ^?�f�>�L����"?5���xϾ5J��厾��v ���2���p���k��e�$�%����ֽ咽=l�?s?�Nq?��_?�� �=�c��,^���"ZV��Z�r�E���D���C�ҙn�-[�<$���ј�W�H=o�H�rM;��Ļ?^�*?������?�=���A��xp���P�>��˾J���uC-=f#�h�=>'7>Z�i��'�ds���A!?���>XB�>�pS?�l�67���?���a�����D�=W��>��Y>*��>��(x��ic���q˾en����ϼ�!x>��b?�uK?'�n?B���2�/��E��Pu"���I��O���A>�i>��>�M�%���A%��>��r�����f���.
��v=#�1?���>��>�l�?�?�	�bˮ�L�n�21�_�8<�h�>b;h?���> M�>� ݽ�Z ���>��l?j��>L�>y����Y!�y�{�թʽ�&�>-ݭ>m��>��o>��,��"\�j��q����9��s�=9�h?������`�w�>�R?:.�:.�G<�}�>��v�׻!�`����'��>�{?̛�=��;>�~ž�%���{�j7���Q,?�?h,��	�,���j>��?���>5 �>1\�?ү�>;7ؾ�5=UQ?��V?��G?�1?���>��_=�ȳ�vW��2��O~<�ڏ>u�E>��=��=�='�9`a��X.�H�<�w�=[�:�Ź��	b<XM���1(���= h?>�~ǿ���vmԾ���������ʨ��L���e��޾�'���þ�h����ڽU�ɽ�Ҍ�5#"����%�~��o�?p��?k{�%(��ө������շ1��O>y�.>!k|>ټP�zv���=��7���>�u����N$��l]��\��s'?�ܑ��ǿ���*&ܾ� ?M< ?|�y?(�9�"�W�8��p >��<O���+��⚚�3�ο\r��<�^?G��>O���&��5��>R��>P�X>�q>����,�<0�?��-?Η�>��r���ɿx���F�<���?��@�@?�?*��C���"Z=��>0|?BJT>�3���tf����>V��?D�?�Xr=��S�P�����\?gη:��A��	�����=|ؚ=�Û<��
��bB>�=�>��#��mE��_Խ#F>|�>�>*����1�W�o$�<F�P>��Ž?���5Մ?,{\��f���/��T��	U>��T? +�>R:�=��,?X7H�a}Ͽ�\��*a?�0�?���?%�(?8ۿ��ؚ>��ܾ��M?_D6?���>�d&��t�߅�=Y6�뉤�{���&V�v��=[��>d�>Ƃ,������O��I��Z��=�r�[�Ŀ�H&�� ���=�$Ͻ�9���[�����f?��)��\�Dվ~c��]ʓ��߽�� >Co�>Xo�>�D?eqD?;.�>�Q>ыѽ����ݶ���ü�=߽���a{|�i��=(˰�����|�b�&��'�\i �`ؖ��5�E&>�F�V{����n�?aO��;?��y>ۛ��:;��E��Ჾ]���{�����kꪾ���T�`�v/�?��P?��t� �Y�#�1����Q�x��G?�������C Ծ���=��=o�����>�
a>g{���A&��zD��n=?��&?�׾�\���Wy<x9�{��=[?Q�?b��18�=]�C?��0=�3�Zp�>��̻�N�>?��>v!�=+]����A���/?��x?�Dҽ��V��>�~������M���I�@>ŵM����;�d�><����N���%WJ����<��X?`ҟ>��'��n ��쏾�Y*����=�Zp?��	?���>�ES?��I?y��=M\�F�'��=V�R?L]?��>�3�����	���:+?Qig?k�s>�p����`�)��:	��R?�n?��?g�����#h��s���r�4?��v?�q^�[s��k��]�V��;�>JY�>���>��9��j�>�>?�#��G��⺿�X4��?f�@`��?��;<�'����=�<?m^�>��O��@ƾMu������~q=� �>7���/fv���YO,��8?Š�?X��>��������
>[���U�?uo�?�Ҿ"��=�,.��n�k9���y>� j=	C���� ;o�����tt@�ZPӾ��þ�</�G>>
@�L���?���6�Iݿ\ÿR����⾻����-'?�ʩ>9�W���HV�sBb�8�(OW��-��N�>Ӂ�>�77�(F�kΔ��wW����T�>-��>��?�T�H����	 �`�b��f�>cW? O�>,:�=����o�?Սʾ^+¿ ���x&6��De?�\�?�(�?_�7?��麹.��t=�?ݽFZ�>L�?V�H?#�$>aA�=ݝ��N�j?wv��M^`�X�4��'E�JU>�+3?C]�>�-�9�}=Az>){�>�_>5/�ĆĿ"϶����U�?܂�?u꾰��>�|�?c+?`��1��]<����*��%C�r2A?;2>�k���!��$=�ْ�!�
?/c0?����@�[�_?)�a�K�p���-�x�ƽ�ۡ>��0��e\�/N�����Xe����@y����?L^�?h�?͵�� #�f6%?�>b����8Ǿ��<���>�(�>�)N>?H_���u>����:�i	>���?�~�?Lj?���������U>
�}?	��>*�x?	)4>2�?�L�:v��W��>JpU��e�=�����9>�st?�;?���>�N]�K��]���H��,�M�:�9�H>��v?��5?RJh>��ɽj�c��%�cn���QA��S>�Q��)��H9>��=.!U>ɔ�<�e�5"�k;?E���ؿ|9���K%�f�3?C;�>	(?%u���w��1���]?P�>�h��������[��ǫ?3��?�%	?��Ծi^���n>Y&�>"~�>��ҽt6��*~���8>B?���|	����n�j��>��?WS@�˭?"�h�S 	?� �L���\~��u�M�6����=��7?2C񾉨z>^��>��=�wv�Ÿ���s���>�9�?�x�?��>j�l?@do���B�"2= J�>$�k?km?Il{����8�B>��?M��@�U@��4f?��
@�p@�^?���,޿������ľK�ξӣ�=%޸=��%>�1ʽM϶�寣<y�<@��Tyd=t�7>D�6>��c>�U>{jy>k��>�c���2�Đ���f����=��\#����^f����`J�O��Ⱦsz;-W�N^5��u����������	I�>�?��8?5�|?{D	?�6V>Ye�>�7#�d���������>K�>N�C?���?z��>)\�� �E�A��Rҡ���龏5��y�<��=?z+�>�3=l��=�m>L	E>�5�>
6�d ��K@u�S�>R�>�.@>	JM>A�>XE<>+�>�δ��1����h�w��̽� �?����J��1���7��褷��g�="b.?Wz>m���>п����2H?���*�~�+���>��0?dW?D�>�����T��6>���ңj�+^>* �j�l�m�)��&Q>il?d�f>�u>��3�[8���P��t��f||>+6?�㶾�Q9���u�!�H��Uݾ�JM>P¾>(�D��m�3����
��yi�|�{=�x:?T�?�9��3氾��u��?��gTR>�=\>(�=7f�=PIM>�mc�O�ƽY
H�V�-=�y�=[�^>z�?��>!=�L�>����P�/�gK�>xU>B>lX@?�0+?��'����ewt��;�7�n>��>�w>��>s�R�+V�=��>�V>);���t��[��?aK���\>����T�m�&�G=W���,��=3�j=*�f�H�D�Y<�~?���(䈿��e���lD?S+?\ �=&�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��H��=}�>
׫>�ξ�L��?��Ž6Ǣ�ɔ	�-)#�jS�?��?��/�Zʋ�<l�}6>�^%?��Ӿ�V�>���-Y��p��V�u�X�#=4��>L8H?W��U�O��>��r
?�?�c�ު��l�ȿKyv����>��?+��?��m��>���@���>���?�aY?�pi>Um۾vaZ���>��@?RR?��>e>�9�'���?�޶?2��?z!I>�x�?Ǔs?X��>$Ru��7/�H��ʒ��m|=l8/;�x�>J>����F�$����2����j�����Qa>T�$=��>�佉0����=ͬ���M��Od���>]5q>-LJ>Z�>�� ?���>�j�>�=�[���$��d��6�K?w��?Ψ���m��~�<�D�=S]�E�?~�3?��`���Ͼ�L�>��\?�Ѐ?��Z?Q��>���1�� 꿿)����.�<�IL>e�>�H�>����ĽJ>�վ-E��U�>�.�><禼�ھ됁��q��OG�>�%!?10�>�%�=l� ?S�#? �j>�(�>�_E�:����E����>΢�>�F?j�~?�?Pҹ��X3�P��塿|�[�z3N>��x?�V?�͕>���������F�	\I������?ug?�U�?�1�?��??��A?z#f>6��� ؾ����+�>�?�d@�pH�k��_��?�?��>d%�������"=��
����~?��H?b{?�� ��$W�;��"v�<�9]�mW�;!<������>�@>�D2����=+�>�5N=c܃��U>�"�;.�I=�o>��=��7�A� ?�=�=݅8���x��t�2�Z��Z>/�>6nܽ�ir?b� ��s�����Is����X�Fg�?ט�?���?��l3��6=�>�[�?�.?�0?�!ǽ��^����8��F�׾|��<���>���=ns���u��h��셿�X޽�P`�W��>���><C�>��?�ZW>L_�>ے���~0�Cu ����ͧ[�8)�~7���A�vd1�q���
'���<2ќ��ݙ>��C�Tu�>�+?O_>��:>�x�>qS�<,�>�~">&Ke>r�>��>�z�>OE>��8��X�R?�㺾 '����W�@?P~e?[h�>�~U�$N�����ɴ!?�Y�?"'�?S�v>�oi���+��o?���>z(��*?c�j=��<2��<�ڶ�������"����>,w˽C�7�hWK��G]�,#?!l?���`о�ٽ����ce=��?d�(?�x)�«Q�^)o��W��R��^�Qg�[����%�H{p��ۏ�h�����x�'�� 5=�j*?��?5;���,����j��?��g> �>ͨ�>Aٽ>5iJ>�M	���1��F^�^�'�i���x�>~P{?t��>�K?�K?ߤY?.-G?�E>��>"�F�>�A����(>��>,*?H�1?Y3?�,?�u3?�I>#������h����>$w?d�?ù?(� ?��4��b����:9��=v��Α�,��=r�J=5������>�佲,=ú?&掾��X����H�>�R?��'?��?��O�}=9���n>M�>��>5��>i���K�D)߾8�>�BT?O3�v�=��U>�l�=�#
���o�Y�>�w����=B@a�%K�P��L[�;"x;��H�g�+�j�ɼ����|V�u�>=�?T��>3C�>A��/� �����h�=Y>
S>�>hEپ�}���$���g��]y>�w�?�z�?2�f=Y�=
��=�|���T���������:��<��?�I#?�WT?m��?4�=?Kj#? �>'+�PM���^�������?JU,?��>���V�ɾ�����3�V5?��?L`�ڧ���)�o���F�˽�>q�.��O~��⯿ �C�Ҝ~�k��5К����?Eӝ?J�>�c�6�,�d��������C?^B�>]ڤ>� �>�(���g�7��:f8>���>��P?� �>q#P?u9�?L�w?�mq>�i�ͫ�\D���S ����k*?A�S?#8k?�n?m�>�(�>ٝ�=X�E���}"���֤=氞�W{�D�>�6�=�$�>4�:>��=��i�̵ �cs��U,�=D�O>��h>!N�>®�>T��>Hc
=GuJ?Ɂ? ��9qJ��\�LT}�Pۂ�0�?�r�?E *?%�\�껇�A�"����?�3�?���?�VX?�8P��r>>;����A���Q�>l�>���=x��>>�{<��&�ql?�	�>7����Ծ��&��#�#�>ۓ"?tBX>��Կ�Ď�J��c���n����������S�����gS��q���Ł������Ͼi:�b �P#׾�bǽX�>�Y�>;c>t�>��=Ē����;}�4=a� >遽^���x^߽)��d07���
>�<�P��z�=JJ�=(r���˾y�}?�:I?p�+?��C?�y>l9>˭3�#��>m���M@?V>��P������~;�����3!����ؾ�v׾:�c�ǟ�(D>�gI�&�>�/3>gB�=>r�<@(�=(s=MƎ=�cQ�a=��=T�=Zf�=���=B�>�\>�6w?U���	����4Q��Z罟�:?�8�>z{�=��ƾu@?��>>�2������wb��-?���?�T�?=�?Fti��d�>T��d㎽�q�=���>2>h��=��2�L��>��J>���K��C����4�?��@��??�ዿϢϿ4a/><�8>�0>-�R�IE1�qX���^�H�U���!?E�:���ʾ��>�߹=�z޾��žlF"=@4>&�]=���-�[��f�=�rv���==�j=�P�>�yD>X�=����!$�=�-E=�I�=�'M>�r̻��?���+� (=���=e`>MH%>X��>f?��7?��e?��>����\��|�ܾ�]n>z�<���>�=:�?>��>�$-?�H?�4D?���>`,�=-�>Tk�>�&�q�۾ $���5�x��?�?�>-���k�+�P�
���:��X���E	?i(?��
?��>78�2��h&���-��ğ��-���.=Np�(]�F���Q���뽖*�=��>^��>L��>I)v>ԧ7>uQ>5�>�>�<�<�ր=������<�`��Ў=>u�����<�K�0���A��Ai0�cB���X$�<$<� �<xy�;8�=���>�
>�u�>���=F1��S�0>����H���={٣�!�D���c�m0{�|++�g�'�T>��V>I���	<��K��>ںd>�aI>���?�x?fB>%�M�׾n᛿`i���E�|b�=\�>�5���:��_��O�оU��>��>Eޢ>�Sl>>,��&?�_x=��\05�M��>5���X�^���q��)���埿u�h��|��2pD?(D�����=O>~?��I?.׏?.M�>T-���ؾY/>������=U6�lq�i둽+�?�)'?Pg�>63���D��ھ�yҽ��>�%[��;E�������*��1�;�-����>F]���ؾ�d8��ㄿ�Z��_�J� ak����>� M?-�?�"�v�w���H�6�t����>�X?G=�>q�?D�?m㰽��ھ8bq��=&>k�y?���?�!�?g��=��>����#>ur�>�Ϝ?J��?/p?��>�>"��=r�>h�廣��;�R�=�Dy>,dt>%M�><��>4�>�%ý��r�+��Y�\���<��'>��?b�N>�<>P@�=���� �Ǽ��l=y�>(؟>T�>�
?A�?���-���6?o>�(�>�A4?��9>��>P��:�}>.*��uc[�0sQ�>l�QI	<)
>�>���tZ���w�>�ο���?�R�>7	��AN?���.���7�=�
4>DN��7�?`��>���=C<�>n)�>@l���n>�[>c.����T=l��G����9�?�M�w{�����>������N� ���!W��pw���Ǿ�l�Wt�
T|�i��h��=�?Xߏ�G \�x�+��&~�4	�>�ԍ>�t3?�ǜ�J���c�=Ċ�>��>�y���m��H ��.�о�Q�?d>�?�!c>�؟>8�X?�9?�0�R.3��Z�\�u���@���d�ǽ_�8S��〿�	�Ig��/�_?� y?;"@?i��<]y>��?#�%��*��Ad�>�M/���:�}4=>~�>�ǲ��\`��aҾ�¾�����E>3�n?�?>?�S��Bm��c'>��:?֞1?�Ft?��1?%f;?���e�$?L3>�8?�l?�J5?=�.?��
?iE2>���=��je(=�4��yي��ѽ$�ʽ�N��3=X2{=�bP�C{	<��=�
�<:GټXc;����<�3:=�B�==P�=ܶ�>\�d?��?�>�4?A�L�EH�Π۾]?z,�#&��u]a�$t�\BϾґ.>�o?��?/�O?���>,7E�M[��o�=Ew�>�j#>�a>�>�C	�1�|�I�=>��=�i>��g=U>;��E5������D�����<7Q*>���>�>5Xn�ٷ+>C��ֲ����X>�nL�J���O�O�E��1�k�v����>)�K???*��=���zu��UVg��j&?GO;?M?�<�?	s�=@�Ҿd?9�rJ�D��L�>�_A<Q��Ɛ��Q���J8��D=��'d>@�������d>_���}޾�n��I���羏�U=���ROV=u����־�}��	�=�*>c����? �8���yv��]�I?}/h=����-�T������>�y�>(l�>ͅ9�ke��iA��4���e�=w��>\�;>�o�쾶�G�R&��܆>>+>?�"�?ی?펽�ax�knS�Q"�0�þr�$=o!?4��>��?Wc>Gܺ>;���f��[w���:�k-�>�(?ۑ��*^�n�vD�KI<�~_�>�t+?�*�4��>v!Q?$�(?X#Z?��?]��>s>=��:�Ȿ�i+?KI�?��=�]^��3o��42��U�y �>�"D?��پ��[>��8?/T?�??&q7?��>��$>��ԾoY��ة>���>1���lA�����>RwP?I��>��m?���?h?s=�O<������=L.���_�UE�>���>��?K�o>���>;�꾇`��9R�= e?H̄?�*�?R�>���>�KT>'��>4bN���}>=��>��?ϹM?uu?4i?FZ1?�<^��v�f�^h�Ry�=�F��L�=;!Q=W��=��&>�V�=z�=�c�=5�M����!v��%���	���ӽ1n�>&w>�Д��(4>_�ž'}���B>�墼3���Y鋾ō3���=H|>2�? �>p%���=���>i��>�����&?>~?�H?���;�Ka���վ�N��'�>�>A?��=Sm�H���|5t���z=�rk?��\?(NX�������b?�]?<e�r=�Q�þk�b�v��U�O?Y�
?�G��߳>g�~?��q?���>��e�T:n�����@b���j�?ȶ=rn�>=U���d�{F�>K�7?RL�>��b>��=@o۾q�w��f��7?9�?���?���?*>��n�;1�T��==��>�]?`^�>����"?GB��ѝϾb���7�����$	������dP�������$������׽8��=F�?�+s?[q?��_?y� �vd��N^� ���*V�������E�E���C�ԛn���W5���y��W?F=��_���;�5�?zC7?�򕾯�?�������%�꾌�>�q޾�S=3��=�pZ�z$7>��Y>2@��D6��־�r#?8��> ��>yk?˯g�,P3���J�bނ��8��{>3hD>�η>d��>���t�Q[�=e��8��R]u��=�>o'b?��C? Bt?{�����"�syp���&�� лz ��G�x=��">��k>�"P�����4�BiF���z��9���������=	�7?���>��e>rb�?�|?#������Q�����/e=�D�>2^?�q�>_||>������>Y�l?���>��>/ꉾ͠�>Fy�8ؽV��>���>��>�m>I�0���Z�0?�������9�E�=
e?5���H�^�2R�>�Q?��8<כ�;Ԫ�>"z����!�f��uI/�ҏ>q?UT�=��;>�ƾ��j|�����1�+?��?i����+�I6{>�� ?^�>%��>;Ǉ?F͂>�Ⱦ��<�?}XX?%@?l�7?��>�%e=�O��vﯽ�*1��ق<7 �>f�X>�8�=��=��-�b�C��j�&=���=������&!<��ݼ!�ԼV=�f->J{ٿ~�R�o)�VH���Ǿ۳�Z�����]�vNB���q�>�p��Tv�I;��9�A-�J�{Ϩ��>ܾ�P]�<��?.,�?�ɘ��`��ׅ���ޚ��@N����>y�"=�f^<�>�yć�\�J��侐똾Z���3$;�J����Q�U�'?L���ٽǿ䰡�;:ܾ9! ?�A ?�y?B�3�"���8�^� >zK�<t2��ԝ뾚�����ο������^?���>��j0�����>ӥ�>��X>bHq>����螾31�<o�?�-?���>��r��ɿT���*��<���?�@WA?s(����I�Q=���>~	?Q�?>cl0���3����>a�?	�?��M=�W���
�Je?p_<��F�Pٻ���=�{�=�T=���GK>/��>�,�D�A�+۽�i4>��>�K#�
��E^�Vƾ<9\>D?ԽS��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=���z�ʿ%�7�J�-��;�=؜�=R��<������n辽m0}��"_�X�ｑ4�=^�#=4���BLA>��]>"u>s�O?CHf?�'�>v>�����:�� f;�υ=�Ti�$օ����W	'�o&��-˾I辜��r��2���!0�^d$>c�O����Ȓ6��넿�Wn�%j9?�$�>����b�r^��@�.���h\*�5�L>XS��$V@�SbF���?��]??L���S��C�������^Yd?/�뽓!���Ծ8ź�o�=SQ=d}>��7>�����T����A�
VF?��&?�5ؾ��R��Nf=�ϡ=�I�<J�
?�}?�����>�"?i�/��Ԅ���>�
I=hը=r��>�\�=u�����#��7<?Z�e?M�E�OXn�^ا>R�Ǿ�����>�\>�k��KC��1d_>MH�=�\�O=+�6�⽻����Q?�}>��/�'2!��7�ߢ=(��=��s?� ?�ʋ>N]?�+5?��=�
��$S����||c=6�W?��n?G�>�#�B;ƾo���	+?��\?4O>1i��侷V'�����D�>� P?�
�>��~��f��1��p�� 91?��i?�e�C����
�e	��m�>f?��?�SL�ϗ�>K�*?g<������k��^�8���?�?@���?rw>=1�G�=��?7q�>�S��ī���������3�=��>=���=J��p�������O?�I�?���>Sao���龬`�=25��k�?�S�?�*ξ��L�����t�wy��!>��g<*�;�{{�����W!�i?��;���̾��ڽ/��>K@_rV�?@�>�t� �꿧oͿ~'�����������$?lS�>H���h�{�_���f�`�:�nLW�������>9�b>��S�����QW��0R������?!9�=g!�>%�v�f��X����P��(#>�1?�%�>k\���Ϲ�?�?�m޾��#w��2�#�p[?ȕ?�
�?'�?#�@>)+̾fG��} ��y*4?-;h?�A0?���=	�H�)7����j?Wg��T`�<�4�/E�BAU>�'3?�N�>��-�}=�9>�r�>PU>�-/�K�Ŀ	ض�x������?I��?�_�*��>�|�?�k+?!b�*0��ak��B�*�s�H�;%A?�1>M���E�!��/=�В��
?�a0?Ua�8�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?n1�>�?���=���>~~�=�ː��<�%>��&>_ഽ�-�>��=?h+�>˨�="�F�0��)K���G�j��il=���~>Əc?��J?¿y>3����ļ�-!��W���*��7{�V�N��ܪ���Ƚ��:>�D$>
9>�`��V澟�?�p���ؿ�i��Gl'�	64?���>P�?���i�t�3���9_?Uy�>�7��+��X%��(;����?�G�?��?��׾RH̼�>#�>uJ�>�Խ��c���A�7>��B?���C��b�o��>e��?��@]ծ?!i��	?($��N���^~��x���6�F�=@�7? 9�|�z>E��>�˪=Tjv�ﻪ��s����>�D�?!{�?���>)�l?�~o���B�>a1=h<�>n�k?/r?� f���4�B>Z�?G���􎿑F�Tf?�
@ir@d�^?�碿0#ٿ����˾��޾���=~����=�7���G>�V]>0(���d7�~R�=�w�>/�>s�Z>�L=���=n8%>�o��"�!���sV���o8��������P��8�` �b񾄽ľ�Ͼ��d�+_����n�g�ӟ��K߽�Ud>��L?��I?���?��?׿P�t�M>�r����\�N[��^y�>v�?�<?~;?��%���羰�q�ڄ��Z��nҢ��`�>�~+>���>���>���>�F>x��=��\>GR�>��=ԫ*�a�Nx���>n��>P�?��>KN<>^�>'ϴ��1���h�^%w�.e̽��?cg��ʮJ�[3��[B��/���]>�=kX.?��>�
��r:п��J3H?����4 ��+���>��0?v_W?��>���I�S�+>J��X�j�E�>5 �=�l��)�
Q>c?�t>`�~>ز0�(�4���O��V����t>�p2?"y����0���z�E� N�Y�U>w^�>ޜ���@����_�{j��pe=v;?h?��]�Rϳ��Kl��V��|�9>�s^>���<�`�=;K>�_��J޽��J��*0=@��=K�A>���>�M>Щ�=wt�>�3���c1����>��I>��+>G5?J2!?�l�/�/�A�<�i�c�8>.��>֊>Z�]=��j��c�=��>�@I>��T=�
�L���!W���>�m�;>����.�<�����M>��<d���N��w�;�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�h�>lu�wZ����� �u���#=u��>�8H?�S����O�v>�#w
?�?4^򾳩��Z�ȿ�{v���>��?m��?)�m��A��@�g��>��?�gY?�oi>pg۾_Z����>R�@?1R?d�>�9���'�h�?�޶?���?�J>pw�?:4s?-��>�s���.���������
��=�(�:�>{O>I&��F�7z��0����j�%"��!_>�w!={��>���=溾���=����z$���Ci�_�>�dp>�G>ʞ�>>� ?�:�>���>T=�"���큾s▾�L?���?k��4Gm����<�Ξ=�u]��g?�_4?�,u��[Ѿjè> \?)y�?�Z?#��>_(�4B��}ʿ��u��� �<�K>���>8
�>R�����J>�Ծ��E�N'�>p�>c!���5پ������3�> � ?x+�>ˬ=� ?Ԝ#?��j>(�>aE��9��S�E����>}��>�H?��~?��?�ӹ�OZ3�����桿t�[��;N>��x?V?0ʕ>t���у���cE��=I�l���W��?�tg?S��?2�?��??��A?�(f>��rؾ*�����>�`"?��	�Q@��0$�}����?@?��>t肽�=ܽ���H�����%(?o8[?��#?�t��`��jľ���<���oJ��t<�Z���>
�>�͓��~�=�>��=\g��O7�[W<ă�=��>�?�=�b>�����\;,?�vG�nփ��ߘ=p�r��yD�:�>�SL> ���^?�w=�&�{����Lr���"U� �?0��?~i�?!0���h�!=?��?[	?B+�>D��n޾��ྉ]w��|x��o�F�>��>m�0�M��� ����C����Ž�t���0�>܊�>&�?�d�>m:]>=`�>>��cu�w�;5���fQ�^�*��y�i���������-���c�;�>[��}�>[��I�>��>�փ>U;>��>�2�<@�->�#�>D�^>S�B>��>,��=}Q�=�z��
2��<S?w����l(���J���ܞB?�b?���>�L9�)���Xj�a�?�u�?���?�.q>S�g�s�+���?���>[|���?��P=5;��+<N���m�����,�az�>��Ƚ�?:���M�\d�~_
?K�?>���[�˾��ڽ���y�n=oA�?��(?��)���Q�"�o��W���R�2���g��i����$�җp�!鏿�M���%��x�(��X*=��*?/-�?Fy�fq�9c��Kk��C?�Byf>�7�>�=�>��>'�H>f�	�̭1���]��'������(�>�O{?㮍>dI?�;?�fP?�L?���>�Ʃ>�ί����>s�;� �>��>7�8?�-?�/?E?� +?�c>�l������Wؾ��?R?�c?�?g�?Jj��!��ێ����c���y�6	��`�{=ъ�<?ؽ*t�C�V=��T>�4?�2$�̚>�m��s�>�I?��	?R��>+�3� ����&�<��L>���>�c����
�SՇ��9	�@;?#��?��a<�L)==	;>�[>N����&~=��=*J����û7�u��Қ�o���5<r�;=��?�X)��wl=
A�=tt�>-�?���>�B�>�>��9� ���Qj�=#Y>�S>�>�Fپ�}���$����g�\\y>�w�?�z�?��f=�=t��=z|��DV�����������<�?ZI#?eWT?ӕ�?��=?vj#?x�>�*�#M��+^�������?s,?VA�>��0�Ҿ\�����@����>�#?z[N�+�����=�b=��%<)��׌>hH���`�C����7��Ƚ�d��&̽L��?�?���=��.��ӽ������"ܾ2�??;��>e>��>Z?
��gk�g���A>}��>��2?0�>["[?��?�|W?ΝA=Q8L��O��������پK�񽩚;?1 �?��?�`?�@?��>T{�TȪ�Z����׼0�"���ɾoZ=}>��>���>�f@>�UE�>V���e�=����ܪ��+�>.��>"5�=��>�s�>�ě>YrC?b��>�I��Y%.����4����M�<%�?D��?��;?�ꎾ�8��#F�<}��YT>�z�?�?�D�>�Z��<�#>���Y�׽˞�]��>�C�>mv�>�-����?�>�s}>5{�>�6;-����E�{����?=�+?����п2�����K`���*�=��4�x �8Dý�,�p��=U�;��Vs���̾����������žK����0�E"�>�"�=���=��\=�nü���<B�)=91=���<޾�����z~j=�?��:�<6�]��d�<�8>�[=-L˾�t}?�*I?��+?z�C?��y>q�>��3�⫖>v_��P!??�U>`�S�Z����D;�gҨ��P��}�ؾSc׾�d�cܟ��>�[I���>#�2>D�=Iч<��=qt=,��=m�N�f=W��=�}�=ډ�=2.�=��>�k>�-w?���諝��5Q����?�:?pO�>b��=Q�ƾ7
@?��>>i+������f��!?���?�R�?��?��h�SW�>����Ȏ�,c�=�����&2>��=�2��Ĺ>��J>u�N@������5�?��@��??�㋿�Ͽ�N/>z�5>ZP>�QQ�L61�J-]�|�c� S���!?W;�Q�Ⱦ'r�>:5�=͚�z]ľ˸(=a05>��x=q����[��g�=]�}��2@=��g= ��>JWF>��=���,��=�QZ=�r�=NQ>�S��_�I���έ-=���=�|c>��'>	,�>�?`.?�f?�z�>�Mo��n̾��۾�/Q>��=���>n�=��.>���>��C?��;?��=?�F�>�(�=l>�>?��>�%���i�յ�����<_�?�=�?w�>U�I�c�P�h���T5�׎��#T?��"?��>�V�>z^��9濚;?��4�8�<�@w=���=k?�_������=z��;9�b��k���Ғ>�^�>/�G>"��=�~<OpW>�p�>6�=A����9�=gV�=ND>x��=Eû�GB<S5���!�=��<z1��Bm��$�{96�h�<�I�=�3�<Q��=
�>U�F>�>�32<X�о��0>�BP�S��E>XӰ��%L��_�S�9���G��,�Ae�>��W>�+�H���m��>J��>g,>>uE�?" r?M��>��Ͻ�� ���`�o�\��d=
E;��;ÿ;�&-N�2�E�}�;��>Bߎ>4L�>&�j>�},���?�oco=��޾�5�Ks�>Jڏ���8��t�n/l������l���9e���N�1A?;r���x�=7�~?��I?q��?�-�>�R�� ؾ�^%><P��ĝ5=i�H�m��蘽s�?��%?�C�>��C}B��FϾy೽���>TSI���O�����!5��`Y������v�>�➾��־�.�C��3[����9�1Gx����>*SM?��?m
=� ���3,N�	���缽K=�>ӝg?�Ơ>5�?/�?�5Ͻ����nx��0�=#|r?���?Ȓ�??p>�*>q���
|v>A��>��?M~�?!v?���<��a>�콠Z>��T���������� �w5����?�p2?�_4?S��6�����h������.��=��=��>��=@:B>% �=�	����">��=9�>��>���>`�>M�?,���)�0?�&�=U�F>�t?�I�>�+>��{��wf>��"<e��8e��iP��l��H=\	C>ӝ>t������>bɿ�	P�?��>�����6?�F$��PZ��m>�[E>[օ�}�'?פ�>��}=LA�>,{�>�����1>�g�=�CӾZ�>����d!�:*C��R�#�Ѿ{z>�����&�5��n���;I��l���g��
j��-��X:=�"ǽ<8G�?������k���)�k���q�?�]�>�6?،����}�>I��>ō>�L�������Ǎ��hᾍ�?��?�;c>��>:�W?�?��1��3��uZ��u�Y(A� e�F�`��፿�����
�����_?�x?,yA?+S�<	:z>F��?��%�hӏ��)�>�/�';��?<=e+�>
*��Y�`�t�Ӿt�þ�7��HF>�o?:%�?kY?TV�כm�$'>{�:?��1?�It?��1?f�;?p��k�$?�U3>�M?"r?�I5?��.?9�
?f2>Q��=lǨ�V(=�'���ꊾ�ѽm�ʽ�}���3=�l{=eL��t�<�=��<���l�ټ�g;�١����<�9=R�=C3�=���>N]?z�>o�>�6?�����6�D��t�-?�N=B‾.���or��^ﾬ� >�j?��?�/Z?�a>��C�33C�yi>+ŉ>zg'>u�]>5'�>�a�s�A�_��=�>@>Ħ=8]���|��r	�搾���<�� >F�>w�>i=S���>¿�憠���9>���F���载��U���4��Č���?��?�� ?؁(>� ׾��+�}Ji��-?&�L?��P?\f�?�@�=e����9�kZ����v�>,�A��h�/C���	��<�0� �<�z>Ӕ������e�>��!���˾����K�Ōʾ0U,�Ȟ5���>k����@��얾��<�`l=\I �F���k������̸[?�l�<�Ԩ�mA~�a�L���(>Ӎ%�ӓ�>܃ѽ���=�!��4���A�����>R}\>�t2�����9��o	���z>d�U?�1[?��M?G����}��
Y�<rǾ����j���?��>�q?�>Q�>�RȾ��.�s��p+���>�A?7�#��B��փ�"���XD��zH>�>�>�I�=�&?]9?w�> ?�??w�>>z>v�q�������?c|�?Ǟ|=tUW��ҽ�4A�'�_�G��>��>}�P�w��>�?<X"?�*#?AZK?m	?4�>��̾L�*���>��>�k��թ��t�>kK)?�`q>�>?���?�B=xX$��!��~�(�����>6�J?�|J?>x1?���>#��>�å�5R=���>�a?��?�=�?�Q=>dL<?\�=ԑ�>���>���>Y-?�ST?NQ?[�A?�0?�<��� �S��ɂ�Om<�;�=QT�=��6=�3�`!b�H6���7�8QV�j�=,ۇ��(��?¼�'R�C!&�6b?'�q>�S��b�>�4�����o�N>�5�o㯾=��������\>a�0>�~?�]v=*����<�IT>�ɜ>��,�߶?��,?�kJ?O�ڽp\��W����w��n�>��F?B��>2C������=s��T�> "�?e[?��۽6��K�b?��]?4h��=���þd�b�ǉ�1�O?��
?��G���>��~?w�q?���>:�e�:n�%���Cb�$�j��ж=yr�>;X�&�d�z?�>K�7?wN�>��b>�$�=ru۾��w��q��d?x�?�?���?�**>��n�14�����`>��޽]?2?�>ƴ��p�"?�0ݻ��ϾgE���_��pY⾅*������z����妾1�%�Ps���yٽ��=N?�Os?Fq?u�_?�� ��c��G^����Y~V�������F��OE�jC��qn�xB�Of��4U����B=u݃���S��u�?��>�[����>	����8���־',�>#ر�y�i���1>�e�tք�"X>�� )W�����?5�?��<>�#G?��c�n=��l*���8�N���#�=y1�>�x�=0s$?��>�t8���!������3���hv>nFc?T�K?-�n?�����0�\q����!�D~1�A���uB>M�>�܈>��W�g]�b3&��,>���r���\���R�	�8�=��2?w��>�6�>n8�?l�?rG	�C@���w�R1���<��>�Ei?���>u�>�;Ͻ�� ���>)�l?��><�>���}Y!�u�{�ɜʽ!�>`ح>��>��o>F�,��\��h��u���e9���=}�h?u�����`���>�R?2�:�G<�|�>)�v�}�!�/���'��>�~?��=Ʃ;>;�ž�'�M�{��;��C")?�8?�Ӓ���*�p#>�"?�R�>	a�>=.�?���>y�¾ԯ��?§^?�4J?�hA?���>5� =?���;cȽX'�"�*=�Ά>��Z>��k=���=����\�ͷ�rB=hL�=@�׼�6��'`<����c<� =�4>�ѿr>>����� ��+�r2��Ն�"z6������X ��vվ�T��	@��`���%��N��7�������v%�j��?�.�?�ͤ�"�~�����bs��B较�>)튾v��=C�[��~�D�ξ� ¾����������tT�s���}�'?z���˽ǿ6���%3ܾ�! ?�? ?��y?��*�"�h�8��� >��<~
�����������ο���b�^?X��>�	�(��� �>���>L�X>RHq>���Zힾ��<�?օ-?n��>��r�۔ɿ����-m�<z��?��@��V?���<R���=*�?��?�0>
������,����>�E�?��?<�=��w�)D��|1?بN��O�-�M��(�=�l�=]Z>����Y>��>߲��������B�b>9�>&
=3����=w�H�_��D�=��W��܉<5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�򉤻{���&V�}��=[��>c�>,������O��I��U��=���S¿om.��I��c#�q'����=jؽ��t��9ؽ��Ⱦ��X�1�b=�8ƹ�*���.�=�©>��>��>yEO?�Mg?�-�>��#>s�ܽ��c�Z����ོ�I���N0��͋��H�P����䨾��羈��<P
�8�&
ľ��<��v�=4R���ן!�BFc��jE�9�-?�">إɾ�5M����;ʾP��k�������ɾ7E1�l�m�%ϟ?��A?ǅ��uU����������vLV?�;�0���D�����=����p\=��>��=D�ᾪ2� T��&?��&?�)��!؋��m[><�����˸)?0��>ȑ�!��>�5&?_�F�&@�Uɗ>�>���>��><{/>f[��8���]?�XX??kA��������>$�þ�?��۴ּ�ei=��<�=�I�>^��=;ӥ�A����z�\����w?��>��H�U{� 2o��3�gAֻ��j?�B	?�+�=�a?U�g?��.>j[�N�^��4��c�=��`?w�?��>���/cҾ"�۽�b?ދ?��>���3?��ZR�l���r6?�8y?��.?���8������!��?��v?s^�xs�����M�V�d=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?M�;<��Q��=�;?l\�>��O��>ƾ�z������1�q=�"�>���~ev����R,�e�8?ݠ�?���>�������j�=�쉾���?��h?0c��������8��:���D>6
>��sh>���� M1��[��"���b��<݇�>��@ݕz���>\yW�[^�d�ƿ�ꇿU��� ߾N$?���>���~�4��=8��uw�@��dL���̾��>}A\>�'��㠾��i�{U��3�o�?��=u(�>�.5�����H_���̀�z�>���>�~�>qG
=]�ؾg|�?Q��:�ӿ_q��*��|�W?�Q�?�Y�?;K;?tk)<7G۾VE:��� <Ug?��<?�?d?��9=�k�6�Ľ��j?�Z���S`�R�4�ABE��&U>� 3?�7�>6�-��p|=�>��>.|>�/�-�ĿQض�:���*��?q��?�s�z��>��?�v+?�k��5���T��<�*��J �!@A?� 2>ϔ����!��-=�dʒ��
?�0?|t�*�z�_?ܘa�p�p���-���ƽ}١>��0�c\��d��N��Xe�����@y����?*^�??�?<��� #�F6%?K�>A����6Ǿ'%�<g}�>J&�>['N>dW_�ܬu>����:�m	>���?~�?�k?֕�������G>�}?|H�>��?�=�~�>
��=�°� -���">���=�s@�m�?�M?�^�>���=�Z9�/�_F�BDR�,&�N�C��>��a?��L?�	b>�>����1�-!��dͽ451���� �@���,��v߽��5>d�=>�>��D�<�Ҿ��?Mp�9�ؿ j��#p'��54?0��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�>;�>�I�>>�Խ����[�����7>0�B?Z��D��u�o�x�>���?
�@�ծ?ji�T	?���P��a~���17�d��=��7?�.�4�z>���>`�=wnv�ʻ��j�s��>^B�?�{�?��>y�l?b�o�"�B�l�1=�K�>�k?�t?�/o���԰B>t�?=��e����L�2f?��
@Au@��^?��w"п�ї��l��@�ƾ.S�=R��=�e>�ҏ��q�=�%�<�Js�>�����=��>��b>@�>��?>�zB>`�6>4���d�"�T>��aŖ�	�A�VM����CVQ�#���B��2��21��0ξ�H��[)����~���p�B8�ۚ�|��=ϕT?]�Q?4Us? ?�`c�gj>2���=b�"�)^�=�#�>w.?�.K?��)?kj�=Mқ���c�������T��[��>�kL>N$�>�9�>���>��/��R>?�9>���>R��=f("=R�
��@h=MvR>�>�>���>���>�C<>��>�δ��/��'�h��w��5̽���?�����J��0��oH��`����k�=0^.?	]>#��D?п�����1H?����7&�`�+���>S�0?�YW?�>"��F�T�z/>¹�]�j�r>K6 ��{l�3�)�#Q>h?F�u>��e>�5�H<6�lq]�"����x(=-��>7�ž�EŽus��`i�����3�>A�f>�m���+��T�����\A��@��D�R?�.�>,<���_�XՊ�u;`��>��i>����y�>��<M�P<?��Ao�F��<��9>N~>W?0,.>��=�ð>���:F���>6\->ܼ->�/=?U�'?���ү�𹀾3n)����>�x�>��{> ��=�KP����=�U�>��g>�5"�H��q>�\^?�ved>�Ã���S��\��1�h=�r��f>���=���I2�1 .=�~?���(䈿��e���lD?R+?W �=�F<��"�E ���H��G�?r�@m�?��	��V�?�?�@�?��J��=}�>
׫>�ξ�L��?��Ž7Ǣ�ɔ	�+)#�iS�?��?��/�Zʋ�=l�~6>�^%?��Ӿ*h�>�x��Z�������u���#=d��>�8H?�V����O��>��v
?�?�^�ݩ����ȿ|v����>D�?���?]�m��A���@����>9��?�gY?Voi>�g۾�`Z����>Ȼ@?�R?�>�9�ӏ'���?�޶?ǯ�?II>���?��s?�h�>v1x��Z/�x6��.����P=d�[;ud�>�S>����dF��֓�3h����j����Q�a>��$=��>OJ��5��9A�=�򋽈K����f����>�$q>�I><X�>�� ?�a�>ʦ�>�z=�g����������Y�K?���?���2n�V�<果=x�^��&?I4?�s[���Ͼ�ը>��\?d?�[?d�>��>��迿�}���<�K>d3�>�H�>�$��gEK>��Ծ;3D�ao�>�ϗ>L����?ھ-��@<���B�>�e!?ד�>�Ԯ=j� ?�#?��j>'�>L`E��9����E�ͳ�>1��>)I?��~?�?�ѹ�$Y3���E桿d�[��:N>y�x?LV?�Ε>����؃��D&E�[PI�������?<tg?�`彤?C2�?�??��A?�*f>����ؾި��E�>!�!?� ���A�J&�z5�[n?8?���>C�����ս�B׼���0���b�?�\?.&?���$4a�cþ���<o%�9K�^��;+3D�h�>�;>�������=^�>�y�=�,m�y�6�E�k<`��=s�>H��=3�6������5,?:�C��ă��Ø=(�r��tD�A�>�dL>�����^?�U=���{����)m����T����?���?�j�?!���c�h�]=?�?n?���>3@��gg޾���iw���x�6��`8>��>��g�r���������O���vƽ�i$����>� �>H�?*��>�A>���>=����$�g�۾2����Q������F���(����� �����8���)ξk���鿧>�v��#��>s?��x>?�>�z�>�
<�ќ>p�;>�>P��>'�<>6yl>&s�=U<
=�2�`�l?}���L;�cǃ�����EeL?Nm>?�Q>	]^������w�UMX?�:�?N��?RŽ�u���I����>kY�>�	��u�>KHm>�u'>��X��\3�����ٽ��>k0=(E:���F�3�����?���>�f=ҙξ~�=2�����o=�A�?��(?q�)���Q�:�o�`�W��S�%y�Ah�������$��p��菿ba������(�)=�*?;�?q�� �����M!k�[&?��3f>Z��>=�>1�>(6I>��	�M�1�U�]�A'��΃��M�>3{?C_�>�P=?.2?�vp?�=?��>#�>[¾�?;Ɇ�H0�>h��>�Z?�O?��/?�u&?�f1?Z
�>���;�h���-о�O?�,�>�.?�#!?�?.�1�FQ �_�o�<�սb��hB�:�>�0��E�����d�=��j>_ ?#����9�q�����s>��7?�J�>7*�>�����Y��<�<���>m?�U�>BU�.r�?x�dk�>Ȁ?�a��=j�,>�s�=瓼oع�:�=�ڼ�k~=��e��M"�t��;�)�=�n�=�;ȹ����~>��P?�c��<�t�>y�?ѓ�>+C�>`?��F� ����vg�=�Y>�S>g>�Eپ~��p$����g��]y>�w�?�z�?��f=��=Ԕ�=|��T������������<��?�I#?WWT?ڕ�?��=?Gj#?�>r*��M���^�����<�?cn%?xc�>@+���˾�e�����ܦ�>e��>o%V����<�u����|��
E>W�+������ɪ� *E�mY	�4_�����"N�?u�?K:w�|j�����#ʓ������\=?�=�>��?��>�
C�q�I�~V��]>���><�>?�n�>X�P?��y?��Y?��X>Z�8��|���e��h+���>pg>?#
�?��?�hz?q��>݅>R'���⾞E��^�C��h���l�\=��P>�8�>���>/�>���=ILǽB㞽a�<��Y�=r�_>]��>��>�q�>�m>` |<��N?U��>�Ӿ2��瞾⦾�!�c�?���?<?Q�:li�lI8�����ѿ>��?ߨ?h�8?��v�Q(>fA����Ծ�K���>\��>�4�>�.�<�s�=��=�j�>��>}�Ͻ6���?B�����?�o??�$�=�xÿ+k{�F���c���iG�݂����
�P�������=�jþa���0���m��\Ӿ�������荙�rL����>�V=$�>q�)>��L=�@�=�>���=�&_=Q��ZA�f���I��`=�U<��D��_D�<~A��V�ʼ�i˾�j}?C%I?��+?��C?nlz>h�> I2���>�Ё��c?�U>�P�����;�J����9��{�ؾ ׾fd�Qǟ��)>�L��{>��2>�;�=��<�[�=�As=��=�[��l=���=�z�=`��=���=��>f>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>bC8>�>H0S��v1���a�vd��k`�ra?��;�Mʾ�.�>
��=���3Jþ-�!=�R,>�rP=�P!�6)]�CP�=1x��G�I=\=6�>��B>�&�=������=%�A=�"�=]P>j�n�N��ӌ=�4q2=��=4d>�#>�|�>	O?j�!?��q?L��>́���R߾b*޾	�|>*�y��?���=�Xt=���>�kJ?��>?�84?'��>iډ< �>۫�>`.�Ř[���R��~�-=aJ�?;�?�}�>�`̼�6`������G����;�(?6�>?�}@?e��>������+��R���S������i=P��%�<B����|�ؽJ�=0K=�~�>G�> �+>lPx>.;{>S��>u=>��=
�=�;���н�ܽ�n���J�=ƿ=:��;�6>ɉ� �;3 �� #<-y=0�=���=l��>�>\��>W[�=v ��9*/>�����L�/ڿ=qb��aB��4d�tQ~�w�.�^6�D�B>�1X>�̄��1���?Z>�l?>��?G-u? >�����վ�J���$e��/S�J?�=��>X�<�?_;�0W`���M��dҾ�>j@b>8�>e�>1wA������F��:�?_C��R�=`Ӵ�,���O7��*��9�L�S1̽��>NM���'<5�?�.?nS�?C�v>j8E>�)��| >��X��&�=�������V7����?73e?�%�>I�����Ś˾;��>l�I��O�ؕ�@�0��t���h��x��>�l���7о��2��T��^����KB�L�q��8�>I"O?��?��b�Wz��[bO�1���ׅ�c�?J�g?:W�>�N?v�?"���G�C�����= �n?,��?�K�?�,
>[*�=#�߽o��>O}?C�?�ƒ?a�~?1a���b?%OD=o	�>���կ=/��=`Y>�E>���>�?!�?�Ͻ1'�A㾅F��Of���Q�	�=�>_N=>��F>.=��<�ZV=��S>���>]��>�ey>|�>5��>忾b�0�\�w?��s��҃>B?�Y`>$�>��ν1�>K�<�

}��H]��T��m6f��>�Q�����=�t����>џĿ<�s?��$��I����?�k��m�>�"C>���>�R'<�,>6F{>�k�>�,�=���>$��=P��>���>FӾ�~>����d!�-C��R�N�Ѿzz>���&�������BI��n��Fg��j�.���<=�բ�<�G�?3���.�k���)�t���g�?�X�>y6?�ٌ�L���>���>�ƍ>cH����Ǎ�xg��?K��?�=c>�)�>L�W?F�?�v1�F#3��xZ���u��$A��e�Ѯ`��ݍ� �����
�k俽��_?�x?�wA?)��<5-z>���?��%��Ώ�,�>/�##;�!<=n5�>V(����`� �Ӿ��þ$E�?VF>�o?L'�?�\?�1V��F�Hɜ=��?4S?�8�?�g?Kq?��=,�v?�r�>|�J?M��>���>�?��?pC�>�30�.T���>/�
�T;���d	��쭾~�n�lC���;E<�5�=-��=*X>�A=�p���׳:�,����;0���� �Pɕ=��+>Fo�>-�?���>�A�<TT?$���VS��5i�.��>�n�sI�<����`�����K�>��`?i��?���?W�>��>�h���X�>��>��=��]>���>!�t<��`��F<Lސ�k>5�����<6�ν�)%�����*��_>?��>T-|>�����'>J���_)z���d>�R�sͺ���S���G���1�p�v�v[�>N�K?��?s��=hb�Y��!Hf�4-)?�b<?JMM?�?6#�=O�۾��9���J�W6�y�>[��<����¢�? ��1�:�F^�:��s>M1��i�P�-�>�>�w�_��`��gD�`�*�`�=�@#�46��jT���z�R-��� �<�1�=r%���A��B��K꫿7T?�[�=�+򾪶���5a��)�<�=�<?�_���h����2���PtW�
P,?è>������þ�zN���nے>��P?�H?��k?j����^�@�$��E����b�8>��#?@?�,-?�
->KV�>3���#���_]�r7���>�i�>���=�(�T��]��=��#�>�B�>>D=Mf?l�&?�J�>�tv?r~�>-��>.V�>��E��+���k2?9��?��_�������=��f�,�V��w$?���>TT~�;��>�$?�!?$�<?�)?�&�>$0�=���N6C����>�4�>?*r�.����>�K?�="�W?���?��<U�>��_�.ү�6�&�{����/?�?�T7?���>H׻>����*>A��>�5?�:1?��^?�d>;?�l>Gn�>�#���L=8�k>�p�>��`?�(w?p�6?��,? � �3]ɽ"K��l��D��2�{���<�� ֨���8�R(�:��=���=�w>�y��<�/��e�> ߂>a���YtQ>����Kq��kb>��>�;7��͏�#8�b�=E��>�
?��>cJ$����=�>"5�>�S��W?��?�U?q����_�)˾ �9����>0;?/�=Xzg�'���n�p���d=��k?�a?��8�&&���b?/%^?����<�
��� `���� 3O?�
?xH��_�>�!?��q?^[�>�e�qn�X)���}b�x=i����=�j�>��� �c�O��>&�7?���>g�a>g��=��پ7�w��\����?�Ռ?Qү?	Ί?,�+>�n�	����;<���]?\p�>�[����"?�1��8�Ͼ�[���&���� 8��~���i������~�$������׽���=n?�s?�4q?��_?� ���c�e2^�`��IRV�\��:���E�*�D� �C���n�Wi�%T�����hbE=�|�
�#�=�?c?|Ğ�P.?cӃ�*���d���J�>r�a&B�١B>����' U>�~Wľ������| ?�x?j��>z5?fl��w0������.T�I�쾰��<��	?��h>u) ?w7��_-�yZ����ž�Z_��dT���v>�{c?qdK?��n? ���0�#5����!��74�����/B>�>��>�|U�Ϫ�8&��>�;s�����P����	���=��2?�>�1�>%�?��?�9	�����ͤx���0�M�<;��>�h?���>���>�vѽ�� �9�>g�m?SX�>$��>2�p���%�+�v�����U�>�µ>�#??��>�7�1�W�fr����0�ˌ�=>�e?)}��X��1>��P?ad2<&�<�>&̷�L�#�W�����D��<>F?�X�=F�=>��վ�t��8��;/���0)?��?�b��|e*�BU~>�"?�z�>/U�>E*�?�@�>�þ�v�y�?m�^?��I?AEA?�l�>h�=H��!Ƚ��&���+=O�>��Z>�em=��=�H��V\����'�E=�Q�=��м9�����<H��I�N<`��<s$4>��˿CU5��̾�d������;�Y�7������>�g�@�Ҿ�ߏ��݇���޽��G��e���������?�#�?|N����j�	�7����A|q>��D��&>�ޖ�'��V���߾�!��R.�Հ��<l�9�����'?a����ǿq����۾�$ ?2 ?�y?��2�"�ʆ8�X!!>���< [��E��v���n�ο㬚���^?���>w� ����>��>��X>W�q>�*��\'��V �<	�?��-?W��>Br��ɿA���鯢<���?8�@�oA?�T���Ծf3�=wa�>,�?��L>2�L�����澾���>�v�?I=�?�~�=�Q���F���Z?�8��';��G����=$�=餂=Z3]�+3>�\�>2�'��/2�s��~hA>
��>��4�`��Vf��=�r>L*�����5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=��������̘)��aQ�Т�6�Ӿ���<L���&=)ve�#O&��	(����7ү���>�f%?Vj?��>R�>�E5?{\U?�V�>�:>�+�Q��Bh��Z�x9��������ؽ>���w�Ӿ������V\������Г�{�;�b�=ѐS�h��&� ���b��H��$.?�!>}�ʾ�rK�Ӳ9;zdʾ�+������μ�YOϾ�?3�Ʒn�h��?�hA?�#��.W��K�+���3Ƚ��Y?����[��ǭ����=h���aH=�٠>�@�=~�M�3�BMR�@�0?�?%���&Ȑ�*�3>�#���W=g�)?8��>Z L<�ѩ>��%?d�'��ս�2Z>�.>���>"��>R
>!�� '�_6?U?������_�>	���:z���c=I�><�4��2ܼ�4^>�g�<�`���6�v��1�<��g?h�?L�=��PR��.�>$x%��b� ^l?�?�!t=�G&?��S?b:�>�����Xa���e����??��)?ű�=����7}��0�^��'?��?:�>*�ξ���<�/��	о�"(?�:?5?JN�=��z�Hܜ��(�l�X?��v?s^�ws�����I�V�g=�>�[�>���>��9��k�>�>?�#��G������zY4�$Þ?��@���?��;< �H��=�;?i\�>��O��>ƾ{�������q=�"�>	���ev����R,�g�8?ݠ�?���>��������>k�m�ѭ�?�.�?i�ž�r�=����^�������=yɘ=9O�G�T=�3��3��ٸ��!�e#�����d�>��@=?V����>p9��&��x.ÿ�������@��4?U��>����u�aPQ��V���2�)=����Q�>�>������)�{�@g;���̼��>@��H�>�DQ�r���՟��!<��>i��>�>����
l��خ�?"��Iο���5����W?�o�?���?:�?>��;�Ex�/Ux���r�bH?et?�X?/G$�}d`��)7�$�j?�_��rU`��4�hHE��U>�"3?�B�>N�-�L�|=�>���>'g>�#/�u�Ŀ�ٶ�@���T��?��?�o�
��>o��?ts+?�i�8���[����*�L�+��<A?�2>���D�!�;0=�IҒ�ü
?X~0?{�g.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?nB�>;4�?�D�=qm�>��=>0�����5=��=X��=�b�����>�qH?L��>��->-$��-0�`�D��Z����d�@�ܣT>Yjn?8IX?�=�e��ܼ�G��9������.�r�b�����}�0><�d>+�a>l�-�����?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Ua~����7�j��=��7?�0�$�z>���>��=�nv�ݻ��V�s����>�B�?�{�?��> �l?��o�N�B�}�1=7M�>ʜk?�s?{Ro���i�B>��?#������L��f?�
@~u@^�^?)"cٿ��u1ʾ�v�������<�7>���a��=��~���
=,Rl�=9V�>�
�>,�>nm>�|>�>|υ��Y*��̡����
�X�}c9�����S�{������e����N�>=��0=UQW�ǃ�MF�����>�U?�Q?8Uq?[��>��/�	�->� ���<�&���[=e�>;�6?�R?�$'?%/�=�N���e�J}�m�� ��(�>yy]>�g�>Mn�>J�>��]>�`!>�W�>���=�ƈ=�$�;�A�<�Z>KҴ>���>��>6>��9>Z
�������NU�J��6���l�?��㾖�Y�$oy�$M��I��{/>h?�Ζ�+9����׿F����??�~�����K��N3>VO-?�Q?I,�=ŉھ��ٽ�`%>ÅN=������=�Tľ���;(��}Pl>���>�k>V�s>�W4�P7�OO�Oh���ar>l`5?r%��I�;�8ls�5�F�!q�L�K>��>�و�������W���i���f=��<?f)?�8ý�{��,p�R^���-U>^�b>kH=`��=bwR>��}��nȽ5F�p4=�*�=��]>$?q)>��=��>�)��VD�i�>dL>>�j=>2�;?��$?/;���肽>�~��11�u�w>���>
��>e�>�_I�Aژ=���>�!a>�Ҽ�������DC��ZL>Q0���j�Ĥ��Pu= ����>�u�=���%SG��]!=c�~?�X��7���z����dD?61?UǏ=WI<��"�k��D�?[�@�S�?�v	�x~V���?U.�?����~�=���>���>WϾ�
M�0�?�Rƽhf��'�	�f�"��?�?��?�E/�������k���>�}%?L)Ӿ[h�>Nx��Z�������u�÷#=H��>�8H?�V��:�O�c>�w
?�?�^�ݩ����ȿ9|v����>T�?���?f�m��A���@����>:��?�gY?Poi>�g۾0`Z����>ѻ@?�R?�>�9���'�{�?�޶?د�?�I>"��?V�s?�k�>ePw��`/�m.��������~=�^f;�l�>3�>�����^F��ʓ�3a����j������a>O�$=]�>�G�'���'�=3ۋ�5��(Yg����>�p>0�I>"�>�� ?�u�>��>	+=�䋽���xᖾ�L?蓏?���l��l=&��=wHT��o?>�0?B8�"Uо�>�\?G*�?��Y?��>���󂛿LW���ִ�I+3<k1V>��>ڵ�>\�����O>tӾ��:�;�>�2�>p���پ�U~�`<@�<�>/�#?� �>GM�=,v ?P�#?�Th>կ�>[E�	!���7F���>���>(?��~?�]?����}3���8�����[��"L>D1x?��?3��>S����h����9� ?O��՗�Ă?��f?�O�+�?��?��>?BB?]�h>�V�/�׾A���ʀ>�!?�<�afA�x1&�j���?�?�c�>�$���9Խ]߼���8���$�?Q\?�&?Ա�'a��þ�d�<�e*��VH�5<�\P�xP>�>�ʇ���=��>�ձ=��m� �5�E�`<
�=���>.[�=Y�6�Tz���6,?
D�Ń��
�= �r���D��>?L>���@�^?�=�<�{����+q����T�n��?��?f�?������h�u=?��?�?M1�>�8���Z޾ġ�vdw�لx��|��Q>���>z�l�(��=���X���fO���ƽ���_��>ǅ�>ZN�>�j�>�ą>�~�>�䉾��(������*�/H����Y�@����G'�-l¾*��w��E�Ⱦ�2���?�>uBp����>�r?*�M>��>�O?��R>��s>糋>Ւ>��>,(r>�>��]-+��c^?�� ���/��쾐|4=��S?��Q?��>݋A�y�ȅ��g@?��?��?�?>d�y��DM�?�>/�?J�z����>Ĉ>�d>�����[���>���`�^��> ���"G��x6�-Ƚ~�?�u?"�=�bﾎD��ޛ��g�=�fM?�a2?�(3�˪/�D�b��)b�c�M���Y=^�ѽ:�׾�E���u��h����݀�N���s�*����q�C?#��?{#�s�N����ލg�~r���<>!]�>�E�>-�>*5	>v�Q8��<9��bB��������>��H?�à>4�A?��Y?>�?�=?���>
�
?|��I0 ?�0L����>���>�R?T/?��?��?��:?�V�>qY/>Υ�@�¾��>�>�>��I?D�*?Q�?=���,�l=9NY=B�$�4���d�Y�C����$>�9��V����ݽdE�>!I?L��<9��+���h�>)9?Ԏ�>u�>򓾼I����<gx�>?�
?�x�>���?ht�����g�>b��?G���Ƣ<O->���=��㼘2<�]�=� �?O=��A; �K�r���4�=m��=(~�;�@��_�;dVj�*{�<�n�>��?I��>�_�>9��6� ����>v�=�CY>�S>�7>h"پw��� ��n�g��Gy>�s�?[y�?��g=�=�m�=儠��E��������Z��<�?�J#?�PT?U��?��=?�h#?<�>�.�O��7]�������?I0?O�d>�s"�e����c���� ���L>�:�>D�~��7�3���?���(Η��%=EOt���s�ꫣ���M�ʱʾ�5�O)罹��?%��?�\^��ؾ\��@�#R���v?|�=+@�=�[
?�	7�
7��#�v��=�$?M�L?r̸>�[?� h?*�<?�s>�@�����'����&��`L>�Z;?uf�?˄�?�tb?���>zd	>4洽��پ+_�;��ýj�P�2�μs�>���=�0�>�>Xb�C<6�?N۽�/��C>���>{}�>P�B>��>Kp>!�<��G?<�>�H����ٿ���߃�R>��u?���?d�+?C$=i���E�
%���0�>�g�??��?�9*?đS����=v ּ�޶��q��*�>bȹ>�5�>��=�G=�8>w��>Ş�>�G��[�jn8��M���?F?�a�=-�ſ�)r�ìp�)W���H'<F����e���W�PЫ=�;����������_�P�ꤐ�)N��V~����z�df�>y֊=��=�^�=�c�<��¼<̼<��F=��<=C='n��5<]-2��
�81��6��:ꊀ<wP=����D�˾�}?Q;I?ɖ+?�C?��y>H>��3�^��>΃���??�V>(�P�>���͍;�Ҫ������ؾ�p׾��c�;ʟ�C>P�I��>�43>~/�=�l�<��=�7s=�̎=�S�u=�+�=
K�=Ib�=7��=t�>=N>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>\�]>�8>id��.�QwP�9�i�~6��:*?x�L�l뾚��>m��=����:��&g��k�>����s���q�l��=Y�ӽ�A�=L�*=��y>�r>�>�<��7�=���=���=wh>�Q=�o����U�=���=�G{>��=��>o�?�,;?�K[?D>�3p���������n>󭑼���>.n*>��>`��>�?��6?ubI?���>��>�ԇ>��>�v���P��	;� ھ�L�=�Ys?�q?�h�>�OT= ����7�!M0�k�=�
�?�{V?+) ?z?�'���濴^5��TV��g���N�C�<�&X��J$;Wq�.�+�m�F��n>��>?��>�ji>HI >�:1>;޾>x��=�nQ�r�=_=�9/����I��=��=�#>�ֽt=����K��G󝽥���h=�t=��=(��=��>�->*4�>���=- ��4k+>����GM��~�=c=���;�ԓc�3|���*��X0�J|G>�T>�)s�<P����?U>3D>W��?��s?�.&>?�)ؾ\����q�f�7����=�>��7���=��b��#S��ݾ:�>T�p>7�>S`8>(�-�C���P�h���G!N��?�2��
��၄��Zu� u��쵦�fy���=� ?ϼ���?�=�9�?*�6?SH�?���>(x=vY����~>�e^�]�a��8��e�G��ξ�A�>?g�?�L�>�������H̾���:޷>�@I�6�O���C�0�	��&ͷ����>����L�о`$3��g������čB�Mr���>õO?��?F9b��W���TO�����(��Nq?�|g?��>�J?�@?�&��z��r��#w�=��n?���?%=�?>�U><�����?��C?��Q?�U�?��?�:=
�M?��Խ���>>=��4>�Z��� }�V<�:|z ?A;3?);>?I�ƽ����Y���[۾�E��dd6�W��cx9>�+>-�n>��=�~��I�>��W=�>��>�F>�>��=�LM�M �e,B?�
>�>|>�E?{�*>};>8���.π>>ܶ��ܽw�-� �꽓Y2=�˺��V
�������
���>�K���f�?IU�>�U(��?���>6>(��>'�<��"�[��>4��>F>���>5"�> x_>7�K>�Jn>CӾc~>���R\!�,.C�+vR�`�Ѿ+Wz>楜�2�%�������4I�>���ar�Ij��.���==��ڻ<�G�?�t��W�k��)�����ޏ?j>�>0
6?Ԍ�~���>���>m֍>�Q��q���Zȍ��rᾴ�?���?�;c>��>��W?ǚ?%�1�Q3�QuZ��u��'A�7e��`�፿������
����:�_?��x?yA?V]�<+9z>ࢀ?k�%�gԏ��)�>!/�';�<8<=Y*�>b*����`��Ӿ�þ�4��GF>h�o?O%�?1Y?{PV��R@��5�=��:?�1?:Ii?�6?�m<?,�U�3?�F>U.�>$�>[�#?\&?f��>xgp>T�)>���i>N=k��쉾���Hcj��Z���>�m=>��=�'�t0�=ͮ
>y�X=��ἥ�<�<F�*D���u;�&�=�۬=4ڜ>oxe?$Z?��->��)?C����0�*DϾ�C�>6�J>m&N�����������¾e�1>��p?&�?'�c?��>�%���B��g�=�F�>���>	u�=���>��s�Ѵa�bo�=CE�=b�>�9r��Tؽ�QZ�����[��_<�!��=���>�X|>7W���'(>dv����y���d> .R������ T�:�G�W�1��u����>	�K?O�?��=as龝��rCf�G)?�y<?dTM?On?�E�=��۾j�9��J�y���"�>9	�<���6�������:�T:�:�t>�֒���wI>T���.���	������𾩦��E��n/�r����T�9���
$�> ����O�1ֱ�������\?�C�=�Ḿ�~��� ��2`�>H��=���>Li����b�"�x��cJ>|{ ?u>v�<s2Ծ��#��"��>>6|B?ʢU?#7{?G���І�ŀZ��ܾ���J.>a�?�v�>�]?�W�C s=�&���%�J�o6���>�?n�U�e6R�j难��۾��U�#�>g ?y����V?#�?;�>�|a?��3?�}�>�a>sK�=q޼�C�-?�K�?巼�ƌ���Y���G�;�m���?��	?��g�{]�>?�?��? #�>�|Z?���>���=�l���7-���>+M�>ݟc�RJ���Ƭ>WQT?��F>��B?&��?3��=�;��ƫ�~(ʽ��>f��<oM?i�?�?�j�=Y��>�A.�#ß��#>�["?R�?��?�]�>Ql/?�"�>L$�>w�̽ݭ�>�'7>�5�>[L�?L��?��W?3	?��<S*=��<£������d��>�����*=��="[H��&��Y>,���|!H<���<�_�kO���vѻФx<��?��>Z�|�仾>����|6�צa>��X����U���V%�L�:>�\=R�?���><*��|�����>�<�>���+?�/?` (?������U��?K��o��?�?��=4�x��2`�0a�K�=<&v?��b?�J���� �b?��]?bf�=���þ��b�\�龌�O?��
?8�G����>#�~?��q?���>��e��6n�����9b���j���=Hw�>�`���d�LF�>|�7?�;�>w�b>�i�=Hv۾��w��x��v?��?���?��?<-*>�n��3࿝����J���H^?O�>������"?�� �@[Ͼ�#��$A��Z������	���P������9�$����`�ս	�=��?L�r?q?��_?�� �E�c��^�<��T�V�O������E���D���C���n�5C��������~H=q����+��?��-?�F(=	e�>�?��,2Ⱦwﾛ;�>�B���;/�>�Z���a�=�^���n�+$��n�2�
	?��>�խ>��S?N5��P�~�B���.������>�h><��>��?��.�©��^����Հ��U����ή�q>��c?o!K?�zm?����[/����ҷ �d@��0���(D>-->I�>>_��b��%��V=��
r�6��Ĵ��49
����=�"4?媁>�|�>�×?� ?'"	�����~���/��e�<ư>V�f?6��>#_�>u佤S����>��l?��>��>>d��A!���{�˽A�>o��>#��>u6p>#�,�\��l������19�RR�=�h?x}���a�A߅>3R?Wa�:�/H<���>�@w���!���򾑝'�6�>Hc?�Ԫ=<�;>��žk"��{�z
��f�(?;�?!u��9�*�\�>�!?�e�>�ϧ>�Z�?�֙>�����7:l_?�\?mH?�A?� �>�}A=p��5+ĽZ%��#=�!�>*�\>Lj~=���=���@X�[��V�-=��=�ɼ̬���KO:�Jż�I%<m�=U�2>�߿4/D�6�;�M����"�+��`�r�(1j���}������0Ҿ[����=�Y��4}b�t���ω��n���?%��?!����������J�b�G�޾g��>M�[5=�7z��λ��)ž����,�C��Ć�Ѝ�[����(?+,���?ǿr�t�Ҿ1�!?�?��u?�����"��8�v�.>ƺ<[J�7(�륚���ͿRh��ʊ]?�(�>`[���%��>'J�>��Y>�v>�T��&`��iQ<{0?�c-?��>��i���ǿ�`����w<��?��@�N?�"����Mx�}[?��?o�u=�o��1#�]�ž7��>��?��p?�>��h�>V��EB?��	/�@A�T�;Z
�=�$>�)½�]>tM�>>n�P���A��O"]>�B�>�e;���H��TC�&�5��y>	x �Q��=Մ?X{\��f���/��T���V>��T?�+�>d<�=��,?7H�7}Ͽԯ\��*a?�0�?��?h�(?�ڿ�?ٚ>c�ܾ��M?>D6?0��>�d&���t����=�2�3j������&V����=Ы�>�>�,�����O��I����=C��ƿ�_�R�'����Z�����r�5���ͽ6���G��w�x�$��G�=�C>��t>$��>0��>�pg>U3^?u?�h�>f�>ر/������ؾ�2;��P�wWڽ���󢉾CZľv;��i:��k��`%�x�%�����=����=R�!y��G� �Z�b��F�n�.?�7$>˾�xM�u<�wʾI媾�ǈ��Y��̾j�1��n�Ο?Q�A?�셿3�V����)?�����[}W?�����֗�����= г��{=ټ�>҂�=9;㾏3���S��O.?�7?Xg��+ۉ�w�=>0�d3=(?���>���®>��'?e�6��Mý��a>n~>O�>?��>SO%>� �����Ѽ?rcU?�S��Ex��-ܟ>�����Xo��=�a
>�<F�)�H�x:>�c�<�����[ʼm.o��=!f?x��>�5��,;��6���=?+3��ga?*8�>C)d>ǳ3?�P?l�=/达��a�f#���=J[C?�*?�>�g ��оT��b�H?��?��>�����k+��a ��Z5?�q4?W�-?�MP��4��Z}�����+�<?�fu? �^��R���?�:IR��p�>To�>J��>O�7���>��>?:�&�2��便�3��a�?�[@��?p�<���d �=�� ?���>�<O�
^ľ*����{���o=�X�>�ѥ���t�L"���(�}�8?=��?��>Ͼ��%��n=B&��?�Xm?�|�c췽n��j"_��Q��'R>ֲ=f!�<��0<�D����]�������Lc���3����>jP@`ۜ���>�����o�_ο%����������O�I?��>9��=GF��IQ���g�1k$��QI��Ǿ77�>6>i������B{���;��������>o���ψ>R�Q��ȵ��ܞ��t<<�>���>��>�<��xQ����?����=ο�����d�gMX? �?�N�?Tl?tD.<H+u�yl{��='��KG?'\s?�FZ?�'�(�[�y�?��k?e`��3`�>e3���C��V>�C2?��>?K.��9q=�A>F��>y�	>{N-�S*Ŀ|���a��;��?�-�?�=꾐��>u��?# ,?W��|)��󬥾Nx*���:��@?g�3>��¾�� ���<��`���?��/?������]�_?+�a�N�p���-���ƽ�ۡ> �0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>eH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?b��>��?c�>H?p��=T���I��:���=���=!����?� I?Ѥ�>�%�=)\+�.��>�F�I�K�T3C��-�>pMh?J?�x6>X����M*�t_�~h��{9��N�Z�S���ʨ���'+>"!O>NAN>��`���̾�E?7��Rؿ���}A$�@3?���>�M?u����u�k�ٻ��]?���>��������:1��.��?�?n�?��׾B���>�H�>Le�>P�ֽ����>���:>cB?1��a���/�n�S��>��?��@1[�?	i�y�?���5L��}��Q��4=����=;#:?��쾹�x>Z��>��=}�t��ĩ��Ws��E�>�Z�?�;�?��>��k?:�n�2C���6=��>�Ui?�
?�������H>9�?���񸍿�Q ��wf?�
@��@��\?�2��T��8d����پ%��b^�^z���'j>�'��_��a��=�6���ؑ��>�c�=��>Ɩ�>_��>i�>�,j>����#�Fi��"㑿-�F��+#�C���Z�����;������2���'����֖G��W��&�=�5���ݧ���2;q6�=�V?V$R?�Zr?�6�>3�^��>&h�&8=�,1�Jm�=�.�>^�,?��K?N8)?^Ί=���%/b���|�����D�����>lKC>9V�>0S�>�%�>�q�:�=R>�9>��y>���=G�=8�����"=w�T>P/�>�9�>�E�>��d>��>r���N��x�w�1��=�	?8��&LB��Җ��"�����>`�#?���=�P��RQϿ���H1F?Aؚ��9��s�[�!>�+?�'P??_!>ڵ����<%2�=�Oɼ�����=���*�3�FP/�5;�>�:?���>�>D��� :�}�y�Rj���|=O�?���y>ވ����΋����>q&|>�ھ���8����� ��ے�� p�vd?ħ>��5>Z�ľ��*��틾�,=eUc>I���D!�>�?�=óD����*�e�1��>{�c=��L>��>����E�,#�>�@۽�������>xy�>6M�>��0?S57?h�@��J�<�KV�Oq&����>k?8��>�Z>��۽%3<v�>�!�>�9�9��ݼ���p!>p��=�\����<QL?>�ᦽ�L>��>Ϲ��a�#Uk��~?���(䈿��e���lD?S+?] �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��J��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿnh�>5x��Z�����r�u���#=��>�8H?�V����O�w>�w
?�?�^�⩤���ȿ*|v����>I�?���?i�m��A���@����>.��?�gY?oi>�g۾W`Z����>ϻ@?�R?!�>�9��'�p�?�޶?ܯ�?g�E>C�?�t?��>� d�>l/�䳿3'���f=~�G<���>�>����bH��N��kw��i��Y��d>=�)=��>ų�b(��PJ�=͏��ޫ���_�q͵>L�r>��I>4o�>sh?��>�ؗ>�U=;�����
���,L?ᵏ?>��MHn����<-��=�N_��7?�<4?&�Z���Ͼۨ>i�\?ѳ�?^�Z?�e�>����%��*⿿4c��~�<��K>�>Zo�>ս���lK>�9վ/HD��Z�>���>����4 ھ��˺�t�>bT!?�\�>�w�=�?-J'?��k>��>�/<�[	����J��k�>���>�?J�}?X!?��  @��P��Y\���U��(G>��s?�~!?i�>{����ơ��6=��j�P�½4��?�ah?J�!���?{~�?�-?�+F?}�f>�Bܽ�A׾j����[>!�"?���RB�=5&�@c� �?�?
�>Tē���½��(��F�E�����?��W?��$?�K��^��K˾$�<Z�W�҄�;B�";�i��x>�>A����ǧ=��(>�m�=I�R��16�OM=<�.�=D>ϒ�=4S'��Z��,=,?�G��ۃ���=��r�<xD���>�IL>
����^?Wl=�
�{�����x��	U�� �?���?Zk�??��;�h��$=?�?Q	?l"�>�J���}޾2�ྵPw�
~x��w�\�>���>�l���H���ؙ���F��o�Ž���ݑ�>���>l�?;��>�{P>C��>s@��k&�_�����;V����J!3�B*��"��/����=�3�o�9sɾ兾�0�>_����r�>�?a�{>��x>��>}���y>?�;>pz>G�>@�T>L�>>r��=��z<�s��]VZ?6Ȩ��#*���þne��JC?��K?��>�D!�q5���T�V�-?�0t?"͞?e)/>w;z���,��� ?]W?�뀾BZ�>�=�~�=�9ݽ��Ͼ���<Nl��+���1��>��7�P�H��=��L�r�?	�?���/��ɺʽ�����o=�L�?�)?Y�)�;�Q���o���W��S�K)�Z�h��,��Ӓ$�^�p�xϏ��_�������(���*=�*?5�?I��m��;/��k��%?��f>>��>��>x�>�LI>��	���1��]�-E'�*����Z�>�+{?A�f>��V?�-A?X�W?�,?/[�>�V�>�j޾5^?�?P����>P�>oe?��	?P@?Ie�>4�?]��=C�=.���P��h�?��> �>�?�(.?>2��+�c��<��+���V�(He=B���=�b����<�Z�{f�>+(?�Ǽ��@����3
�>B�A?럪>!��>�i��\s�����<J	?4�>�x�>b;��o��ʌ����>OP}?��Ϧ �k:>y,L>Ih���8��{M>�j߼��;�$���=�{_������>0+�=P����~���=!=�=[�>��?"��>1B�>`!��^� �ݓ��=��Y>h�R>a>l'پ�}��t��p�g��Ry>s�?�~�?��h=��=�9�=Rw���8�����㽾m�<v�?�A#?!HT??��=?D<#?^> 1��H��^f��{좾�?G.,?�;�>V����ʾF�����2�1�?��?�Qa��$� O)�I���_�ؽ��>��.���}� ǯ���C�y`����q���}�?��?f�@���6�����_���֬�
]C?7��>���>e��>��)���f��$�fj>>]��>�yQ?\��>'�Y??�g?�~E?)�f>O5�~����������%�=%V?R�}?�C�?�x?��>��>i
[�LkȾ��A��\�h�/�m���<��u>���>���>v>�>YrB>�������d4��w�<j~;=v�?D�>칵>��[>��>�lG?�6�>`�Ǿ���A������%FP�e�v?r>�?e�)?��!=����^9��������>\ɦ?Y��?@W+?3U�b2�=�w��R��H�i��~�>�q�>��>��=��+=G�>��>��>I����*<��O���?�>?�*�=#ݽ�ġ���������ġ�=+����BF�ۻ2�?����n>#ӽ�*:0�.'���u?��ľj���n�Ӿ��I��i���>�҄=�`�=���=�_�=F(�WJ�z1={���y�>�;�����<ef������P��(=I�ʼ<%�=�%=[���� |?�N?�y=?��2?r��>\,>���=�>�O뽞w?C!S>N��xe��^3�]դ���b��۾�۹���i�;��E�->��(��=vV>qy<>�A�<
>�� =��=kt�;e3=C s= 9�=ދ�=F�>ɀ�=�I7>�2w?���.���2Q��T�}�:?=J�>K��=�tƾi@?��>>�1��钹�
b��+?W��?�T�?i�?tRi��^�>I����ӎ��C�=����)J2>���=|�2�\��>s�J>����G������2�?;�@�??ދ�*�Ͽ�K/>2�<>�P�=;KT��.���S�h	f��[H���$?�E3��-¾�L�>oχ=��پ�
��Z{=�8>��g=y���Y��Ф=׻��28=�u=M�>!<>Xj�=��ٽ��=���=LJ�=4Ma>HE�;�_.��g���={I�=�D_>��
>��>�%?D�-?�3O?sH�>�vj�d|�*��>ZĻ�/\�>�9#>Q�z>e �>y&<?�#2?h�X?$��>Um>�-�>��z>��%���[��������jk|�I��?��?�8�>`��=�0�_)�|@>�$⧽�?�O)?d�?�ӥ>�U����nY&�c�.����G��+=-lr�NU�I����k���e�=Zp�>c��>,�>�Ty>��9>|�N>��>7�><5�<�q�=�������<�������=����$�<;|ż\[���.&�Q�+�����!�;Ȗ�;��]<h��;���=U�>��>+t�>y�=�f���.>w���� M�8�=�����sA�ad���}�
�.��7��8B>uVT>����B0���?�T]>�	?>k��?�~t?�3">���Ӿ�2��Twg�i�S� ��=g>�|<���:���_��}M�.�о�m�>+r�>å�>3bl>^+�
�=��v=�⾠06����>O�����d^�M0o�~����ӟ�چh������$C?_���M�=h�~?�I?�
�?���>�ǆ���׾޷5>\S���=0��in�$⓽��?N'?�>X��! C��G̾16��ѷ>�@I��O�����8�0��J�����_��>�몾/�о� 3�f������(�B��)r�� �>D�O?^�?�?b��W���PO�?���Y���k?�ug? �>�N?.@?����o�f�����=a�n?J��?09�?��
>n��=mX���>�z�>�Yv?���?��?���x�?��G�zAo>k9��0'>Ph6>���=l��=<�?V�?!/?�v���h��������"��*�=>.=,w�>L�=>Mh�>*��=�>�H>Z�> �>�>�r�>dܶ>'P�>��������X?� ��
�>dc?g,�>��=2�%���>Pn��F%�	g������Ϩe�1��G8����������jj>�	ǿ�P�?�-?>~�E���>'S̾�<�={�>�¤>�"����q>'j�>�~q>3�A>L��>�P��2	?,t�>3Ӿ͋>u��Rd!��C��tR���Ѿr^z>H���&&��������II��_���l�=j��,���9=�~��<�C�?�����k���)�d�����?0b�>�6?t㌾�"��L�>h��>۱�>w9��M����ʍ�Kkᾒ�?���?�;c>	�>A�W?��?�1��3��uZ�S�u��'A�9e��`�X፿�����
�!����_?��x?�xA?1U�<H9z>:��?d�%�ӏ�%)�>�/��&;��?<=,�>*����`���Ӿq�þ/8��HF>y�o?R%�? Y?�SV���M�`�V>�%@?��2?9�`?�j@?�'G?��4��,-?�K�=��?B;?hT0?�-?�
?��+>]S�=�9�7�_�=!Ε��/��aj��7�X���?a�<H�=T��=�����Y<;�.;�X<H��=�M=":��H;�c=��=_�>�̌>4�V?���>��>V/?��H�/	�ô���F?1r��ɦ ��T=�Sw����޾�c7>s�U?�I�?>\h?� �>�nD�Ac�{�>�5�>��>�C>�y�>��<�E��U�=N�I>Wo�=p�Ľ��/������W
��';���=%�4>>j�>ɀ>�b�g�'>�Ҡ��u�T$^>�`Q�nּ�*QP��YF�&�.���n����>� N?��?��=^�꾎ʓ�^+e�t�%?��=?��N?��~?-{�=��־LT9��OJ�4���>iS�<���j��KM���<��/<�b>X���������w>��:��QC���*t��c����=�!޾���G�޾S��y���>�g>sa���2��C���Y��/�g?�'�����+�����p��>�:ǽ���>�\I>���a�"��#�TUP>��?�b>߷���.��_�'��+�vKT>�*E?�vX?,:r?V]�c�_�+�>�Y����ȾM~Ӽ�$?D��>K�&?�v>U��=rȊ���rB��9����>~�?�*��:(�N�~�J��Q�$���>e��>���u?�S?�	?/�^?G@?8��>ʛ>3�=��㕾�G%?�K�?�/�=O�ѽK�P��7��E��>�>�u&?W�E��,�>�?��?��&?NQ?�,?5m>�U��:O>�5(�>��>cwW������b>-�I?s�>��X?'�?K�3>�Q4�#�H��(�=M>CA1?q�#?9?�{�>���>p��� �=�P�>Ia?-�?��o?L��==?Z$2>��>K�=k�>!��>�u?��Q?�|u?�M?��>�y�<������Ci���
��&P<Z�2<�;�=���`i��&��x�<Ұ�c����ʼ�m�H�"�mc`��R�;L�>�6�>��K�M�>w�W�l�̼=�>�4��|d��y����T�L�X=�s>�\?�4�>@n	�t�=y�>i��>�u9�v"?�%"?��!?�.0��:���\���W���?Y5?L͔>�q��<.��G�l���-��ی?WU?l�Żվ,�b?*�]?�s�=�|�þ߸b�����O?��
?��G���>��~?H�q?���>��e�5;n�]���Db���j��ڶ=�b�>R���d�\D�>Š7?�B�>`�b>&�=|e۾H�w��g���?^�?���?}��?%*>��n�H+�p���ZN���^?Gg�>�?��< #? �ӼϾV������k�������N���j��{�$��탾�ֽ�Ǽ=v�?�s?�Qq?��_?=� �h d�10^�����pV��$�w���E�uE��C���n��^�F$������`G=jR���A�;�?Q��>�]�����>�6}�ǵؾ5����C�>����Ž,�V>����C�=�>k'���P�������?J?ކ>"�B?;5��6���8��V��"����<���>�X�>=?P{�= ,��m�ꈼ�� ��P#��Ev>`rc?�K?J�n?�5�51������!�H80�p��ݷB>��>��>C�W�����=&��P>�S�r���r��d�	��~=��2?��>��>�L�?y?��	��[��lTx���1���<�?�>M$i?]"�>qֆ>�нR� �,��>l#l?Z��>d��>r���b���{���ѽs�>�P�>���>]�t>G/�i�[�i|��Uq����7�4��=��h?<���U�a���>�lR?\A$9f>8<,��>��n��["�K�3�'���>O?+��=@?>>�ƾ�z���z��戾q)?j"?�ْ�O�*��N|>�!?E��>t��>�҃?��>��¾�]k�� ?�_?t�I?�EA?-�>N�%=x=��<�ʽ��&�O]/=N��>��Y>��l=�n�=���	@[�O��i�?=���=@��
�����7<*Q��C�H<��=�h6>1
�/)>�*ھ��������=�sC=\֣�.ؾ}��F�E��_�a"��8W��J�$mB���D�\�������W�?k��?C�Sq�0����Җ��s��4g>Y��:�>M&���C�ͼI�¾=�8���4���|�q$l��c��P�'?�����ǿ򰡿�:ܾ4! ?�A ?9�y?��6�"���8�� >`C�<�,����뾬����οB�����^?���>��/��l��>ޥ�>�X>�Hq>����螾�1�<��?7�-?��>ǎr�0�ɿb���f¤<���?0�@J�G?��Ԁ��Y��=�I?8^?�p7>}�k�$��?˾��>$&�??9s?_6���)Z���ӽoc?�&���(������P�=֍�=�n�=)_��D:>#��>ے	�Zei��ڽ�,>�tb>Ȗa<����:�R_��v>!N۽��Ӽ"Մ?E}\��f�o�/��U���Z>��T?@/�>�I�=�,?k5H�O{ϿϮ\��&a?f.�?���?�(?�޿�vӚ>x�ܾ�M?AE6?z�>!d&�N�t�:��=L��E ��f��}'V���=��>Bn>�p,�5��<�O�����U��=K�?�ƿ��$�{��X=�5ٺ�R[��k��ت�_rT�e ���io����.+h=���=��Q>�`�>*1W>�*Z>RgW?��k?�:�>��>�J����?ξJ���a��<������F��tӣ��R��߾��	�������u�ɾT�<�~,�=o�S�P���!��e��?C��e-?��>�[Ǿ/�K���C�m�ɾx)���}�����}�ξ�v1�
mo�ny�?�A?'4���T��A�W#��-ҽ��U?�l�%;���
Z�=tp��*=u�>���=I澺�0��gT��8?#�? +ɾ�Vj�/b�>�@|��z=�?H�>����M��>x�8?d�P�-��>c�=SU�>+Z�>�->�B��r���*�?s�N?J=׽?�����>���e�5Z= +�=��*��D<'�>��j=G1��lR&�qv���]=�uW?�]�>�*�����i���p�_<=av?�?O�>�Kj?5�C?ށ<�>���[T��^�l˂=;%V?�i?�
>�E����ξ����?�4?U�d?мN>-,f����I.�@����?��n?%<?e���ML}��ߒ��[�P\6?�u?��^��럿G��]kV��Х>�T�>] �>2�7��)�> �??�q&�r[�������R5��u�?2z@�|�?$ӝ<*K �=�=��?T��>�P��Ǿ�l������jf=L��>%�����u�*���Z-�}�7?xD�? 2�>��������v�=J����s�?QI|?�ã�F�<�9��d��R	����=��=#-�]s =�	ᾞ5�m&�����݊�b=Y��y�>�@B?�\��>�,&�(޿�̿�H��%s̾�߱�֦?���>>��&�c�b�a��<i���8�gC>�����ʸ>�>iu��9��Y����I��^���?�p�=8�A>7���u׾�g��>Y��>��I>W�P>�l�I������?T��c��UK���a��t}?/h?�1�?�e?k��=Sz�V���#R�=��T?�+@?,�W?��X=�
����>!�j?�_��kU`���4�)HE�1U>�"3?�B�>;�-��|=�>���>�f>�#/�n�Ŀ�ٶ�����=��?߉�?�o����>b��?ps+?�i�8��^[��}�*�nk,��<A?�2>#���	�!��/=��ђ���
?"~0?	{�D.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?ֵ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>eH_���u>����:�
i	>���?�~�?Qj?���� ����U>
�}?K%�>��?�a�=�a�>��=dٰ���-��X#>���=\�?�L�?�M?�X�>&��=&�8��/�$PF��8R�u�!�C�$�>�a?"xL?�b>���M�1��!��Iͽ�[1����@�]M,��[߽�\5>4�=>#>��D�c�Ҿ��?lp��ؿ�i��p'�v54?���>D�?j����t���_;_?�y�>47�,���%��A�l��?�G�?�?��׾�T̼8>��> I�>s ս��������b�7>=�B?��D��\�o�7�>���?�@�ծ?i�]	?�#��L���\~�$����6�� �=X�7?�	�@�z>J��>�Ϊ=�qv�����^�s�ں�>%C�?�{�?���>��l?�}o�e�B��1=�@�>�k?k?��o��
�^�B>f�?��n���	L��f?�
@,r@��^?Q袿!hֿG����M�������=���=��2>��ٽ�[�= �7=�8��2����=�>n�d>5q>�'O>-a;>��)>����!� r��H�����C�������Z�+���Xv�z�P3��~���B���4ý>{��2Q��1&��B`��&�=��U?�R?	p?(� ?-1y�wQ>���="=l#�<�="V�>؃2?��L?�*?.�=#���@�d�eA���㦾Ї�L�>�[I>�^�>��>a�>���:�@I>Y�>>���>�Q>��&=*��x�
=��M>�:�>'��>el�>�l�>ܽ=XT��{U���}u��\��˟��U�?K����%�e��������?w���>�i?���=�C����Ŀ`y����,?�#¾�N�W�G�)>08?�&@?X��=6^��=|m=�|�=]�����#=9&�|ʷ<�sC���>>�u?�)�>�ҽN%���o�Rto�������$�z&?�x��k6>��n�`�0��8���=;��>�L=n�\�����]�h���˾#�=s�_?x��>����H(澽���	�^ =Ma�>���B��=-�:=|���K��S����>��<KWy=�J?�,>��=���>[���N����>�H>ou&>�<?�$?2?ڼ<�ޣ���,���o>9��>�ˁ>�D>]�B����=���>��W>Fl�����J��i�=��U>����_�@xZ�z�G=u�����=���=ν�Z�;�(�
=�~?���(䈿��e���lD?R+?i �=,�F<��"�E ���H��G�?r�@m�?��	��V�?�?�@�?��F��=}�>׫>�ξ�L��?��Ž6Ǣ�Ȕ	�.)#�iS�?��?��/�Zʋ�;l�|6>�^%?��Ӿ�k�>+y�[��7����u�]�#=���>�<H?�L��A�O�->��r
?�?�Q򾎧����ȿ
yv����>��?���?��m��>���@����>ߣ�?�_Y?{�i>�e۾#QZ����>��@?�R?� �>B;�G{'���?c۶??�
I>���?��s?1g�>a!x� W/�5��#���s=QfY;e�>�b>���]F��Փ�>d��D�j������a>�$=K#�>�y��*���H�=O싽NQ���f����>��p>��I>�[�>�� ?Ym�>��>�j=G���π�������K?t��?O���2n��G�<ş�=#�^�'?�I4?k[�N�ϾZը>ܺ\?w?�[?�c�>'��H>��6迿�}���<��K>&3�>�H�>�"��FK>p�Ծ�4D��p�>�ϗ>����?ھ�,���b���B�>se!?f��>Ԯ=F� ?|�#?qHj>�-�>WiE�9��T�E����>Ϭ�>�=?��~?h�?�����E3� ��1顿$�[�3N>��x?X?Ӫ�>χ��\�����C���G�ꈓ�-��?�jg?�
彖�?�2�?[�??}�A?��e>�Z���׾譽�	�>��+?j�R�\�I�Dd9�Pd�h�?(�>��?l4���O��ȼ{D�n�۾|?KXD?�y*?k�<_�yW˾�W���͢��[=yս�����,>�W:>�&%�B=�HT>�{6=�S�z���'�߽�T>E��>����Y+���2�I:,?lUH��ك���=��r��vD���>�SL>u�����^?<Z=���{����y��U�L �?���?�k�?~޴���h�~"=?��?�? �>�N��6޾����Uw�5ux�]t�	�>���>F�l��ߎ��3����E���Ž-���E�>�>F�>	��>�>>�>U�����GѾ��.&V�K
��1���5���ꚞ�*V7�����P־c׊�rm�>q�P����>�
?ǫ�>
.�>�~�>^�ռyA|>@W>���>�-�>�Y;>��7>�>rx�=�މ�=)U?������!��à�FBG���F?��]?D�>���?���L����/?j��?�+�?7�>G�z�
@��,�>��?���??z�>���;�5�v��E����r߼�Tʼ���> �޼22^��"��aĽ2,?�}?��W��������,����o=�M�?��(?z�)�;�Q�
�o���W�/S�̕��5h�i����$�$�p�9쏿S^���$��+�(��s*=ˉ*?�?0������ ��x&k�^?��gf>��>�"�>1�>�vI>�	�ݾ1��^�RM'�����Q�>�Z{?�DJ>��Z?� 6?��9?@�9?I�>��8>�-¾�t�>˚��
��>�{�>�Q?�	;?�1?�\?3*?���>,�5�d��̴���?�0�>(��>i��>ч�>ɔ��f;Ƀ6��E��త�X/%�el��x�=AU<X�:=>v�=�Z�>7�-?�Z�C@9��ݾ��>ߜ6?pX�>ܮ)>	���/ʩ�L�˻\�?EP�>Wݏ< �v�d������#y><Ct?<J5��ɼ���=�>���:X��=b�=4����:>z��ʞ�R�@=���9�+>o�k�4'�s�M�k�R�a�=E��>�?}��>���>�&���� ��J���=�;[>��S>��>�پ�����0��\2h��y>���?���?�	q=ӕ�=���=�}���r�����i��`��<��?��"?�UT?я�?U�=?�)#?�>��R&��F5���
���?�a*?&��>��
���о�ʨ���2��?��?��^�,｠�-�Ӝ¾B���>D�-��|�L`��l�E��T��_[��P��k�?�1�?)�ۼ��5���ھ����e���t�??7n�>b�>tZ�>�&��bi�����YI>�>STM?�֢>�W?��m?�G?�
R>�a!�����BK���X��#d�=��8?(ey?�Ә?bc�?�9�>B�0>�;�M��35ﾓ~����$�no��t4�<K"Q>��>�>Vh�>��>d�Y��I��q>E��̨=�L{>&��>��>*��>�]�>�>)�G?ey�>����o����]����9�بu?L��?Ea+?��=�_���E�&���M��>�<�?��?�K*?��Q�U�=7
ۼL����Br��(�>�M�>�Ș> �=7�D=?%>���>���>R��Gj��c8�<�L���?��E?��=��ſ�zr�|g�RO��vn<������a��
���o\�q7�=ُ������H��r&^�9�����n�A��P{����>�҈=�=^�=�d�<-�¼��<�%I=�<��=��S�� t<��#�Sg�R���7���GI<#*J=�
��}˾ȍ}?�5I?<�+?�C?
�y>'8>��3�e��>7����=?"0V>��P�E����;�٭��N���ؾq׾��c�?ɟ��@>�RI���>�A3>zC�=�؇<�0�=#�r=���=ָP���=�(�=:�=za�=��=2�>}^>�6w?X�������4Q��Z罥�:?�8�>f{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��D����4�?��@��??�ዿТϿ6a/>���>�A>\�=�ۥ���=��M���4�'3?$C�M:ܾ��k>�1�>0����M��A=ht�=��L>^
��g3����=y�Ƚů��/<꼬��>'�F>
�q=�<e�Z`q=U�=�&�.n�>x-�|���hQ��5�;�~K>@�2=�Ӑ=QE�>-�?�0"?�=W?i�>�@�J���3����>�uW=B-�>"��=�ށ>X�>��>?go)?�Y3?��>W�0>z��>��Y>e�+�:�^����[���Ph=݋�?a�e?T>�F=�J��:/�G�9j#��]�>4<7?��?_�^>�U����,Y&���.����Xs3��+=�mr��QU����[m�,�㽥�=�p�>���>��>#Ty>#�9>��N>{�>��>�6�<lp�=����K��<G��u��=H���%�<Xużۖ���o&�o�+������;=��;B�]<���;#?�=�k�>�R>��>ۑ=�$��|�.>�����dL���=�����A�d� �}�T/�E�7���@>[U>M6���D��C?�]>B�@> ��?J�t?%m#>A����Ծ�&���ii�(S�Z�=%�	>�?�VQ;�J_��L�ADҾ��>��_>��>�3,>
0�#�;�!��=��پ�,����>��Ⱦdl��*�x>h��_��d��{e���Q�[ ,?R�����=���?��H?92�?��>}�y<߽�W�F>E���,l�����4J�(�-��9?7J?�f ?�y��pt;��I̾B&���޷>�BI���O�U���e�0����7·����>���о�%3��g��������B��?r����>ܸO?��?�<b��V���TO����28���o?&{g?��>K?)A?���y�s���n�= �n??��?�;�?f>˝�<��a�>e�>�}?J��?�?Qf�?��K�!?���7��>d�/��d?��I��5���%d>��'?$�?ˮ/?J�������{��{Ѿd䌾�����=Ts�>2�>�^J>T>��=�C�����=٫>1�{>�>�Z�>��t>�E־�g=���L?�m�=�f>�!?�}�>�e>SӖ;3q>�乾Y�-��5V�c���w�a��;�쾽��=~½T�>���:�?��=;����h'?eҾN1�<�EL=��>��S>:��>"��>Lm>�_�>˩�>�m�=��>���>RaѾ�A>��W���D��>S�}�Ҿxu}>���Y�'���7��tTG���G^�Ck��恿P=���<E�?���{j�G�*��o���@
?���>�n7?=���-��HW>�>�>g_�>����]���	��2޾�%�?���?W;c>�><�W?�?p�1��3��uZ��u�B(A�e���`�j፿ݜ��ȗ
����'�_?��x?1yA?�U�<�9z>B��?��%�/ӏ��)�>�/��&;��?<=�+�>x*����`�T�Ӿ��þ]8�YHF>y�o?7%�?�Y?TV�|�m��)'>��:?f�1?�Mt?��1?��;?G����$?�f3>�E? r?�P5?�.?~�
?%2>R�=�Φ�x�'=�/���튾�ѽ,�ʽ����3=ML{=�ʜ�u<l=���<p��w�ټF};#
����<	':=��=�*�=,C�=��\?�2
?sr�>�|?�|���u��i��G@?���	;�c�#���{��-&H>���?jP�?��?�Z�>�U�����">
��>(�L>��>k�>
�����"���>>�q�<D �=-ս w����Z��뾅���A
��-�=n��>Awu>����J8!>n����,y�Ȃb>�(S��o���I���H��1�I(z��#�>��J?�v?��=I�����|�f�x�(?�">?ߘM?�?<�=`�վ�8��H�����Ę>�@�<��������K��BS:�W<�Pw>T����y��~�>��!��}������l3�����7=Kh%��[�6�uC������\�I��=VK��W�6�i��������O?L��=����q���%��<�=:m&=�ޱ>��佮�q=U�?�N㪾���<�!!?��O>��=��5u����I�>@o@?�hM?[݃?o��ٜ��ec�j-��h�;�.`<ui?\L�>��7?�=5{�=�b�����g���	�|�>+#?�
M���O��m���$�*�~;�>b�?P��y�?�H?�Ae>��C?�Z?r�>�*A>����A����e?=Ƈ?I����@��%��-�d�N�`�5.�>�?^ꃾ���>v�?k"&?�<?8k?��?�<X������ʓ>� �>��^����Z�>^	?�S�>+.1?���?U�{<��L�;�|�Ҽ�vw>�F>�h?�O?l�0?R��=���>�+���d>�>,�??MC�?v��?1_�>��J?��>�M3?�������$�>��>�A?y?��\?G�?S�;�9U��(���ܽ)���p�<��>�j�<ކ�����*��%�%=Tv>Ӗ���=>����č�������=X!?��>K���*7�>}�r��\ƽR9�=�<&�^}��g��>r9�q�H>-[�>�*?W�|>!����>6�>��> ��z?��(?\H?Ee��]�D�
;���p�h4?�q�>|��>Ԙ����\��3�=Fsg?�n? ��kP���d?�`?�� ���>��&��?�j������V?��?�;n��z�>��z?�i?���>����Y_�$���}�R�yn�a>�ݓ>��*�5k��7�>۲R?���>��2>�.>�3��4���2l���?+�?�!�?d �?��K>9�V��������-����]?�F�>!�X�"?̖��BϾ8���K���x�_��1���镾P���f&��ჾ?Aֽ5�=�?�s?3�p?��_?:�Xic�$�]�_���|V�� ������E�OnD�b�C���n��%������I�<=,n{�*��v�?�?5k��8%�>�"־)����X���>�����1��c>�Z)��EV<�~�=^,��8Tr��C��C�?�5�>2Y�>�G?r�Z�uuI���;�Aa7�'��v�Y=^��>vJ>a
?�j�ς�EA �\�߾�J��{�8<� v>;wc?��K?�n?� �R61�����3�!���/��C��ʮB>�Y>"�>�aW�ͯ��1&�L>���r�����g���	��7�=5�2?��>a��>�8�?�?�	�bg��Jx�Wc1�惆<H�>q�h?p�>Z��>+zн�� �}S�>ۜl?F��>�1�>v��$]"��{���׽�l�>`�>C��>�bm>C�� gZ�@���)��[�8����=��g?gd����_�w�>VR?���9�v<�h�>�$���#�;>�y�$���>�s?i��=�,>\ƾ	$�L[{����>)?�N?���ƃ*��R~>�"?!^�>i�>�.�?��>E,þIT��?��^?4;J?VA?�q�>�h=gD���_Ƚ8�&���,=`~�>u[>�m=+�=���" \������C=�K�=o�̼����?<Z���e�O<���<�4>�bͿ�D��gξ���$e�ǡྥ��y9ؽUS�2����]�Z����1羨�������nL�Dxd�H5a���
��?%��?m��8d�.����@�8ܾ$pS>q�ܾ�C!�@,��"��� �ݽ��ﾇ����l��y�3�r;���X��Z�'?Ӷ����ǿt����5ܾ!" ?g? ?�y?���"���8��� >u�<�ޜ�z��������ο¦���^?F��>q�6����>9��>r�X>�Sq>M��2Ꞿ��<�?Ո-?ء�>9�r�f�ɿ���j�<S��?/�@�~Y?�ZѾC9,�NL�hL?��-?Q=�J���o�ׇ�&�=m�?��?�L�>xDb��+ ���/?�񉽎P@��D=���<��<�e$>�[���>�?��������V/��P"=S��> ��=���=r�X8���>�X����r�5Մ?,{\��f���/��T��U>��T?�*�>T:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=n6�牤�{���&V�|��=[��>c�>,������O��I��U��=�����ǿ*^�-�5����<����b����d����;�uh�]Qp�(	���;<��ȸ=,�=�7���<>E�>(b�>U�R?�>y?h�>��R>}t̽`̊��\��c2Q�ء[��M<͇����A����C��bH��;��+���.��l�3����=�R�`f��nn3���O�36���?�=���YeC����'�׾#>ԾO۲�54-���̾p�4�z2{�*�?"�S?�����]�����΂���M?�I�����¾��=h3=��=~s�>�5�=�|��'�2���h���1?��?#N�����{Q7>������<�-(?N.�>��<�w�>�(?ݔ&��7��x�Z>��#>�y�>���>�+>������ֽ��?ԾV?�G�k/����>i����g�W�]=�>J�G��\��W>�I�<�����ρ;@^���T�<��V?���>�D,�����̀�`KY�-�2=�Dw?�E?��>\c?1�A?أ�<bp��M�o+�ʒ]=��T?H�a?~�>:���ؾ�����n2?��i?B�m>�[��W��n.�Ī��E?��p?{z#?[W�m^~�S]�� ����.?�8k?��Z��l��0	�����B��>�G?Y`?�����>��2?�3�E놿<-ÿ(�"�u�?b! @g��?�>�ߝ�F6=��>N�>�`s�1��o.��1����=_��>�_����[��w���D��b3?���?f�?s�i�����W�=���aŪ?؋�?����ɏ�����]�{������=h�=!�-��^a=qﾔ�(��5��L���������ݐ�>z=@[�Q����>��\�zK迖�ÿ�b���O߾�h��,L$?�n�>���*m��TQ�Ζd��<�t�W��dm�H\�> �,>\꛽z����$k��?�(ݤ���>D�1��
q>^E>��.���菾�I;�>m��>ÂY>�����O����?\%쾜�ѿ0ߢ����L�a?�ś?ʣ�?�J#?���K��΀h���C�auJ?��v?0jS?g�� � �Xvӽ4�j?�a���T`�p�4�WGE��U>�'3?oM�>��-�m�|=5">̀�>Lj>�&/�y�Ŀ�Զ�7�����?K��?�g����>&~�?�k+?m�#7���_����*�w�.��2A?^�1>Z���\�!�T4=�{В�,�
?R�0?|_�$*�]�_?*�a�N�p���-���ƽ�ۡ>�0��e\� N�����Xe����@y����?M^�?h�?ֵ�� #�f6%?�>d����8Ǿ��<���>�(�>	*N>�H_���u>����:�i	>���?�~�?Oj?���������U>	�}?�P�>��?���=�X�>���=H����0�S�">��=�9>��n?��M?�@�>���=�8�72/��MF��=R�����C��>u�a?/�L?�a>[����1��� ���˽X1��v㼍A�p�,���߽eP5>q�=>,�>��D�B�Ҿ�?�b�6IؿA+��w�(�S�3?���>��?[��?�s����RG^?�t�>����ϳ������� ���?
E�?�?�"׾pDμm1>���>���>[�ؽ�#��	V����3>W@A?��� ��@Tp�樆>O�?+�@�ͮ?�Lh���?���L
���2w� \�m4���R>�#E?g�¾lLi>/��>J�H=�d�r����kj��	�>GB�?�i�?��?�d?��b��8�eU�m�q>�&W?��>��<]��^��=>�>� ��:��e��)UZ?
�@��
@p7a?�6���ۿ�S��� ־�0��@�=:>�7�>�c��2�<�ý���<nƐ�0��<�3{>~>G��>�(>�5�>fۍ>g���"(��_��NV����6��R澐}���(��^�iL9�������ٱ����>�~J���;����X�� ���"�=�@I?�#X?ċY?+c�>�`��ȋ�=މ�W;݌��'V�W�>'?��C?��-?��=�
���e�	]z�;c��d���f�>m>���>^B�>��><g�< ��>0�<>Jb�>�x�=J�h=o�e<�Z�P�X>.��>�)�>�>T�A>�'>���i��f�j���w�j��ӟ?���$J��I��#Ȝ�> ���y�=ol)?~�=a��PX̿﮿��G?x���c�><�>_�+?@Q?.�>#Y�������<�=����I�t���.>�]���S�Ѹ,���b>-4?۠�>O�Q>`[��pR��䄿��q�=�M�>��+��U8>��?\3�mg�04�=S�>��%hG�7䇿&���Zc�������b?T��>v�&>�M���J���?�N�0>E�>��W�⍰>2�L>������<�����o>�#�����>u?�_>A�k=���>�N8�v��>.ng>07V>q�>?;)?4�x��|���舾x�%��|>v��> ��>=]9>e1:��x�=b��>��8>H)��4Q½&�	'�YK>F⺽-~�͋H���e=�����=���=G�ڽj4���=�~?ߦ������sJ���rD?�@?��=}�G<�"������\��¼�?3�@�?-2	��{V��?��?!@����=6��>뺫>�.;��F��y?v�ѽ�ᢾ��	�/&��r�?	�?  ����� l�NH>�$?;Ծ�n�>�g�[��:��`�u���#=؝�>o7H?�Q�� P�5>��y
?�?�Q�Ϧ�� �ȿ�zv����>0�?V��?��m�MA��@�/��>]��?�kY?^@i>%g۾lmZ��{�>$�@?�R?s%�>�?���'���?�ڶ?���?)W3>F��?P�x?L%?��I=nHB�SJ��pꐿ�ֻ�񄼨��>�r!>��߽��1�S͟��5����l�;/��m>p�=ػ�>]�{�L ��Xl�=�սV(� #�F�S>���=ʯz>/$�>���>n��>E�.>@�W='�)�3�[��{v�L?O��?�,��n���<��=3`���?��3?��r�gWо�˩>�\?C̀?۽Z?��>�����������_���Ȓ<��J>M=�>~��>�Â��6M>@־�-C����>���>x��]dپ〾z��Pv�>�!?���>�,�=|` ?��#?z�k>˼�>��B�.���w�G����>�b�>�s?�w~?9�?���2�ݑ�K"���\��H>�#x?ق?�>����X{���}���&�H��M�? �g?�&轨7?�+�?�M;?�XA?EBt>��־G��{w>��!?tu���A�T�&���z1?��?6��>�Е��gսH�v�7����?}�[?G�%?D���`��þ���<,�/�V}����;��I��7>j�>$��۸�=x�>!%�=q�k�}6��k<Fy�=7��>��=;E6�Eݏ�=,?I�G�ۃ���=H�r��wD���>�JL>8����^? k=��{�����x��	U�� �?��?Zk�?w
���h��$=?��?<	?s"�>�J��W}޾��pPw��}x�`w��>���>��l���>���ϙ��wF��=�Žii����>s�>�0	?���>b�M>Yp�>W��L(��h�:���\��#��7��9+��:�#;����,�D�!���ľ,����>�}�Ő�>�$	?{�d>
@�>�z�>��W��u�>��V>�~>N��>n�R>:�9>�8>@H�<�Ǳ��d?F���:�:�K�������M?��4?��D>�9z�B]w�s
,���d?R�?L�?�L���x�dH,��f�>)*�>�+|����>�Z@>i��=��V<�˾��q��3.=P�\����>�G�j�6���M���]��� ?V��>���,����y̽Fc����r=wO�?�:)?hc)��R�)�o���W���R�����g����M$��Lp����G�������(�bv,=�l*?0�?�5�f�cɬ�!k�9G?�G�e>R��>bc�>D��>*K>��	�<�1��7^��'�<k��O��>~.{?�È>��P?Ϻ'?]?�@<?��(>��1>9�
���?9���]��>6vp>�-?�:?u�5??�>+?�>)�[@�(ָ���&?�L?�4?���>�z?�e���!����">��=@��<�}�=��<�J��Jk���b���� )�>�k0?<!���kM�e�޾�8�>�J?~�>-�.>9���c�����r-(?q�?/h�>O�"�U�|�N��(�>�[?�:,��`�/h>Δ>��=��b�z�=&���]S��P��=�
������	=1C�=wp=�(�G��m �;c1O=�G�>R�?Y��>jf�>"���b` ��D�p
�=&kZ>W�S>S<>!pپ����� ��l�g���y>k��?�u�?�j=��=�#�=k����!�����Z����S�<:�?�%#? T?Y~�?�=?�6#?uc>y
�*<��w`��� ����?/�)?i4�>�Q�6��.��K?1��X�>��>�"l�\	I�ͪ>�tm˾�-�Nq�=n%���r�ش��$9�]n+��	�K������?�ؗ?
��֡$���ܾ��״���K?�F�>]��>�w?��8��=�H���>f�>yaE?o��>DP?��z?��[?�/[>!U:�ܭ�3ٙ���d���>�??�9�?f؏?�>w?M�>�O>X�.��㾡����s�F�ｖ����N=�]>�c�>ŧ�>��>q��=G�ҽ#����8���=C^>�Z�>�+�>���>�x>�S�<h�??�q�>	����N�hc��+Yp��d.=�t{?먑?چ%?$�=r��{�9�$����>���?m�?+};?��ý\�=��>}��ށ��}�>A%�>1n�>�l�=�Q=?
�=�ڬ>�>i������1�C;�;�#?X�D?���=�<¿^p��
1�1�����<X���%�p�j5�u�]�Z�>64��:t�����yc�<���{���Qg�����t�|�uY�>�;^=��=��=��<,���+�E�ghX=��=�Q�<���kXc�蟼�r�B��2�5�G:��g��=J�B<+�˾ g}?QZI?�+?޹C?�y>��>�f2��y�>Y���y?qCV>�P�?x���9;�y�������ؾu׾B
d�Uڟ�b~>�H��>9A3>�r�=�׉<���=�Nr=a@�=ăU�0*=[L�=F��=�k�=6g�=�Q>w�>�6w?X�������4Q��Z罥�:?�8�>z{�=��ƾp@?��>>�2������{b��-?���?�T�?@�?6ti��d�>N���㎽�q�=L����=2>o��=v�2�R��>��J>���K��=����4�?��@��??�ዿϢϿ4a/>��@>�q>�_T��7�����6Ei��ef���?��>�|�Ǿ�f>˅=,H�qi��� �<߆!>2N
��P���d�N�=�?��j�=*�7=Ci�>��3>#W�=#�Ƚ1%�==��=t��=~?i>NDün�c���p��Q�=��z=�w>>�Z�>m�?��E?�yj?Ff>n�ͽr�l��"��b�>w�=�?�z; =���>2-X?��y?$�`?�ٹ>�5:>y��>@�r>�z�E(}����%�޾�^
�7�?��b?y��>�e=�Fѽ��۾��*����J�$?M0D?w��>�g�>� ������;��@X�;#��K�>��|>	��3��Y�ڃ;8��F��� >G��>�W�>���>�ŕ>�e>���>g[�=c�=^.�=䀛=�>U<�<���O"=!v:��^�r��=�T�<���<O�d#j<9�)�a��=�;�Hጽ���="��>D>��>���=j��$@/>����~�L��ٿ=K���*B�4d�8H~��/�GU6��B>.2X>���
4����?��Y>�o?>G��?�?u?��>D�D�վVP���>e�IOS�ɸ=C�>��<�yx;�Y`�@�M��uҾ���>}��>O�>bk>W/,���>���t=��d�5���>�Q�������#	q��礿ԟ�e�h�M�Q���C?4<����=�I~?w�I?���?>d�>���>�׾�B1>����� =���a�p��t��*�?�'?���>���-�C��!̾(z�����>�QI���O�5����l0����z��x��>�Ī�P�оL3�+j���=hB��r�-O�>��O?��?�b��L���ZO�E���ۆ�oN?jtg?% �>�?j	?�����j�T���sD�=�n?u��?�:�?�> `�=iؽ4��>3�?Iۃ?F�?g܅?�<��X?��=]�>M�2���}<�cK=:��=
�>�C?�7?h�?J�f��G��`���Z�������	���=ż|>>>>&>-�<Lb�=��%>R�	>���>�ʍ>�W�=28�> &�>�6�����D?%U|=+x�>�Y?�m5>'��= ��bqi>��3�9�߽=y7�n����084=��Ƽ�\>�����s��>�㼿��?���>�(��&�?ې��l��<<��>t/.>������>��h>��G>a�w> ��>ǯ�=QƸ>��>2EӾ;�>)��Hd!�,C���R�I�Ѿ�{z>����&����{��j?I�m���f�
j�3.��v<=����<�G�?
���5�k��)������?�Y�>}6?ی�J����>l��>�Ǎ>�G��u����Ǎ��i��?:��?-<c>7�>l�W?��?�1��3�uZ�I�u�L'A��e�%�`�X፿윁�u�
�O��V�_?�x? yA?&\�<9z>��?v�%�uԏ��(�>�/��&;�,I<=�*�>>)����`�t�Ӿ��þ�9�HIF>�o?%�?Y?�QV��'i��'>� ;?�V2?��s?M#2?�F;?M��?%?p73>�c?u�
?~4?y�.?�?�42>X�=1,����)=�ӓ�pJ��D�ν��̽�Z�^�6=�L|=��Q�h�<�=��<��g�ϼ���O��8l�<�@8=?�=���=�C�>2jL?�?ik�>��?�E����P2��S?��O>��{T��(R��D�þ�}>�n?[�?�]?,J�>{�V��]�*E>I��>�n�>�><��>���=F�����j>"�->��<=$��)+�%�ƾ�d-��蔾9�=� �=���>��}>�r���)>e����|��oa>�3T�c幾]$P��`G���1�qdq��J�>ϹK?�C?߱�=3��j��<�e�@!(?r=?_	N?��~?T7�=H ۾K�9�	K�z;��:�>Y߹<Bm�.@���N��;��~��[�n>X��AR���	a>z��PϾ�)t�'!L�O�۾�!1=�+��4,=���[^ƾ󕃾��=.&>�lľ������_�����H?�B=�؜�_�]�`��D>9��>���>1M����v�>�F������=���>��>.S��&󾌯E�	��c>O�P?�~P?��?����2���DG-��M�����>P�?L�e>�? ?"�>��:>�*��ko뾍4��x��z�?��>�w1�o=5��(���S׾m�G�҉�=��?)Bn>�r?�n�?��?{eZ?ˠP?�?���>�	>\�����'??ê=��w��Wj�
TC�N�e�"��>]?�U0>�O�><?_|"?��:?��e?B}/?z�L>{���RO�x��>z�w>��3��"��D��<3�+?6ĕ>�c?P�?��>K�%��i��<1����p=��[>DAI?FY)?�@:?�7�>o5�>�ĕ��.Һ΋�>Yd?�[y?2ao?���=M�	?�-[>�F�>ʄ�=)�>h6?��?�E?�j?_:?*�>��<=&\н�j1�ł����G��=��9���;��X<��Z���}�<�5S=�}�=�u^��}��C!ڽb追<
��:�>�rr>l�־�E>�w��sp�&?Y>A�<@�>�_�����0�#Q>�{F>$��>|��>�3P���a=���>;ͣ>�v�)�? �
?�>?gZ��pzc�����`��9�>lA?%16>]�j�{퍿�mx��c�=�Q?a�H?TV*�|��B�b?�]?h��=��þC�b�ԉ�e�O?5�
? �G���>��~?g�q?V��>��e�:n�!���Cb���j��ж=Ir�>CX�:�d��?�>f�7?�N�>^�b>n$�=�u۾�w��q��s?�?�?���?�**>��n�L4���۾�2���1W?|��>�on��cF?m˼�����'���#ƾ���7þ� ���7����ɾE{a�I�y�%���<��?	dj?��|?ן=?*�
��	d��_���k�ܡ]���	�����zF�Vn2�Cni�H�~���"�G������=b�~��jA��i�?a�'?��.����>yf��'K�_�̾1�A>�����m�ϭ�=�,����<=�"X=4�g���.��z����?�>���>Km<?�[��>��1���7�{����2>%k�>a�>j��>,�߹�.�����ɾ�儾�fҽ5�>h[h?��d?�]`?���u@	�^ˀ��x��M�Q�3�=�# ���>Y�5�n{P��J)�D@�O6��S<�W��1%ݾ�g��dU?tU�><IJ<���?k��>� ���I!��œ�B����=�?�ώ?SJ?M�>m�P��[���>�!m?=]�>^��>(�����AA��@��h��>�ï>1F?ݩ)>�.���Y�����֏�|^A�U�=�j?�_���"\�c<�>A�P?�����9#=�˝>3*�$���|�-�@�p$�=��?&�=j�x>@�������쀿o����?1?�e��4��pK>b�?��>M��>�r?�6�>�Ѻ�=�0?f$q?*qV?��<?��>�̈́;�
���N2�UW�S��=,�>=ӊ>��+> ��=���#)㾝 ��r�+��թ=&�=�q`���=|�����`�o�7��<>�n�ON��վ��$���޾ְ�س���?����B��}Z��!��Y���e����r<C(�� p��R�uP}����?oX�?j�ھhZ�������u�}. ��,?��Y�7��
�ȾB�<����{�|о�"�5G��U���g���@?��
�ο�����k���5F?H6?b�t?�h�Y#�
�0��R�>q�f=��Խ����V���п�h��m\p?���>d�"���7�.@�>�?���=��b>�����%ž!��>	=�>>�(?���>�3��ſ������>�T�?	p@�{A?��(�7�쾎V=���>S�	?�?>I1��F�����>O�>u<�?���?�wM=��W�
�	�v{e?�<��F�3ݻ	�=�K�=��=`��ϊJ>[V�>u���FA�)ܽ]�4>�Յ>��"�_��ˀ^�h�<͈]>(�ս`6��5Մ?,{\��f���/��T��U>��T?�*�>T:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=s6�����{���&V�}��=[��>c�>,������O��I��U��=B����Ŀ+0��(�q�<��H��
������m��>ǽ�����[��I��	�=�:#>=s>L�r>�c>�m`>�}a?��l?��>p@�=G���\����:����=5�B���\�It��P��Ԃ��z����Pྭ��UQ�h5��8ؾ��D�i�Z=v�k�/l���A(��U���)���T?M>.���v�2qs>�ɾ�x��`�<r$'��,˾'�	���]�⾸?]?�̏�� 0�};1��*2=�C��H�a?!�	��8�]�C�\�>�,¼`)=��q>/3���M��v $�$���Y,?O�?��ľ�i��ޗ�=q����8�<�M/?�?�`W<�\�>X�(?M�����?&{>�4>�T�>�X�>��>��o��8�?v�Y?'��.&�����>{�ƾ��~���=+F>%�9�9�ؼ�"@>u9�<�����ʙ������<ɀU?��>�&$�_���'���AR����<�w?��?�0�>��j?9^A?�3=Ι�ҰH�G+�Wg�=e�T?�qc??��=K}k�"�ʾñ���J4?cf?m�R>��O�l,��~8�0��0?�r?`�?m��}�� �����y�7?�~?q�n�����B��=V�I�>K?p?!�,�S��>�l?6�x�����Sſ2�'�p�?�D	@=�@�O��"�֑X>~�?
��>!'۾����)J�E/ƾߕ�=��?H�������f0�_�K��?��?�$"?����-*%����=�N�����?桄?�E����=�J��n��	��A�̪�=������c�i�����@�G׾�-�������$�+u>#i@�|���8�>Î[�Xv⿝5ο'~��e�N�e��?�L�>���x�Ͼ�`r�gu�zF��D��2Z��d�>��>��������� y��{:����`�>���|�>!Q����qd��w�j<��>B��>o�>�<��/{�����?�b����οQ�����|ZX?�Ϝ?[�?�?' O<�m{�ܒx����G?��p?
tW?7���a�<;;�T k?�e��X�`�6R4�HTD�u�U>�3?(�>v-��;}=>��>P&>�.��qĿ�ʶ�F;��^Φ?Q��?�꾶1�>~�?�9+?4^��K���R����*���:�XA?��1>c���c�!�==��h���7?��0?��S�X�_?�a�E�p���-�|�ƽ�ۡ>��0��e\�lL�����Xe����@y����?I^�?f�?���� #�`6%?�>a����8Ǿ��<���>�(�>�)N>'H_�v�u>����:�i	>���?�~�?Hj?���������U>�}?�>�,�?ՙ%=�Z?��#�\F��`
=/��=1�2>
�a�w?��R?I��>z��=]���.���?��D����»>���h>�If? 1N?Gc>l.�0��ߡ"��[����7��Lb�M�P��F������>W$>���=^<8�Z�߾�g>?�[�!EͿ/׃�p�=\�?DI�>b��>I ˾�������\?,��>���d!�����H�I��j�?Q�@S2�>�;����'>U"�=���>V��<������U-�Ӗy>+�A?�mf�n����x���>^��?��?���?P�D�� ?cn'�����el�k=��Q�j��!>��C?v�þ�>C�?��=�=z�H﬿�`���>��?/��?�c?u�E?1�;����#��Q��=D�a?��?r�=�c�h55>��/?�2#�����^��@f?"�@x@�p?����~Tտ�	���������`��=`�=�9>�׽n�=$B=}�1���w�Qi >�ט>~�h>�`r>�YR>�=>[(>t4��?!�#Y���t����B��F���\XX��
�>�q����R����ڿ�#c���~ýP����R��L*��e���=KNS?��N?8�n?��?t�!�?N+>F%����=����c=Xh�>q�1?y�L?�)?w��=T5��>4c��Ҁ����鷈����>ChL>���>���>N��>9^��vD>w�8>ͤ�>���=^� =���T=�N>�ت>���>���>b*>�>����\㱿Z/r���Y�#�ʽ�ئ?��>M�4����Z+��ѳ��E�=u*?��=�����ſn"����N?C���0&�l�#�\&=��-?DST?�
�=p��'Q�`�T>^��-`�?��=��0������n"?>�?�c>�1u>o�6��8��T�L��[0z>�/8?4A���~@�w�t���A�'�ܾ}M>�<�>'e��(	�xO����{���]��_u=��8?1�	?zZӽt����i��y��)6]>�d>`�Q=��=�H>�=w����%!N��0=:j�=��V>lu?t�->�?=!��>U����^�;��>Z-/>�UB>��;?��#?�iN��+��q��"���Ah>K6�>SW�>�,�=09L����=��>��b>�͸������\���=���L>�c��5�Z��z��۽}=�ͩ�Bܿ=+�{=��9�;����<�~?���(䈿��e���lD?S+?U �=X�F<��"�E ���H��G�?r�@m�?��	�ߢV�?�?�@�?��I��=}�>	׫>�ξ�L��?��Ž5Ǣ�ɔ	�/)#�iS�?��?��/�Zʋ�=l�|6>�^%?��Ӿ�U�>fKV��՝�u���V�}�`��=�T�>��V?OԾͪ/��Qe�)�?�>v������r�ɿ
9����>���?��?u.��R �� �F�oZ?S��?�;E?�k>����!��� q>=1?(K?���>!0�dl>���>/��?�,�?eo�=�Ë?*@�?<�/>�˼3Z��÷�8���-Ī�6	����>CǗ�e��u�c�Y������킄��e�~a�>�N��O2�>]V=�ƾ[�A<(�A=�⦾]�=|�>��>�dm>O��>��>���>�l�>u�=Sl���r���8���K?I��?S���0n�/��<�Μ=�_�Ŵ?��3?;�\��gϾ��>o�\?�̀?A6[?u�>Ռ� �����f���r�<�L>K��>[��>w��K>�<Ծ�E�>�k�>S���ھ���,8�����>B!?�@�>��=�� ?��#?�j>q)�>�aE��9����E�1��>H��>�H?��~?�?�Թ��Z3�����桿��[��;N>�x?V?2ɕ>���񃝿�ZE�7@I�����u��? tg?�X��?�1�?��??,�A?�&f>����ؾ����
�>�!?�����A��5&�u.�\�?�e?�t�>YJ���Խ0�ܼj��d���;?�\?�"&?q��a���¾iX�<�A$�,S]�YW�;4�I���>�a>���Vݴ=��>�W�=�pm�~|5�A�p<�8�=��>�]�=�7��Ŏ�"d/?���U*�nI�	 �� T^�2ΐ>bo>/�_?��ν����A��� ��2����?���? ��?��?�~�T�`?�kx?'�!?j��>��3��$�ⶩ��־�c���r>�?�7>y���eǩ�,���'좿�3������>��>~?v�?.M�>|�>}��7�f	���ؾS�V�g����8�%�=�.�`ݢ���V�k�9��^��O���=�>���;*c�>�G)?�	T>��>��>U��<���>�>��|>U?���>R� >��>rf��O�ֽ-�P?ɾ�:�)��4�����A?c?|��>g�U��]�����x!?XO�?ʆ�?L x>�h�A3*�k�?���>��y�W	?Q�@=Ǳ*<���;�ᶾ������p[ڼ�;�>Y�ýk*:��ZL���i���
?;?;L��R�ʾ��+ߌ�J��=n��?�&?����N9��Er�pP[��kg����́u�6�ྷ5��Ix�4g����G�|���.��9�=9�?1�?C�۾�2�х���%��f�I�2�B>C@�>���>�N�>��=j���o�@���^�)R%�e#�����>FA�?�.>>U�F?�:D?6K?FLD?�P�>�h>� ��v�>z<�<�o�>��?�K?I?a�U?A�?j
(?��>	U�=��-��ž��?G?�?���>��D?���P����{�8m=ӱ3� ���P�p�*��D��Џ�<��=��<>�?6i�ɻ8�bb����l>��7?�+�>
!�>x9��-��f0�<���>s??�>�G����q�c���*�>J1�?�d���=�j*>��=���4 �:���=	�Ӽ%^�=줊��A���<�c�=�u�=)9��	w��T ��9;�x�<�t�>(�?m��>
D�>A��H� �8��}e�=Y>�S>�>�Eپ�}���$��R�g�X]y>�w�?�z�?d�f=�=���=�|���U�����0���m��<�?!J#?�WT?I��?W�=?`j#?��>-+�eM���^�������?!�+?�p�>J���ɾsg���"3���??�_���'�(�E����׽	�>�V.���}�����ZC���»#����_\�?��?��F�<7��k澀�n쪾tWC?h��>�У>���>�*��3g������9>;�>�P?�$�>E�O?�:{?�[?�^T>՜8�11��@љ�� 2��">l@?Ӱ�?A�?y?�w�>H�>��)���T�������\߂�d�V=lZ>���>�'�>z�>P��=�Ƚ`a��~�>�'h�=+�b>n��>��>o �>�w>���<�bF?H��>S}������J���l����꽫�q?���?�C?��=g��gs:�4�ξ]�>< �?C;�?z$?�"f��K�=�Β�����|)�����>S�>� �>t�=��;��N=aƵ>�"�>��ҽ+���8��੽#�?�hG?[�>��Ŀ��o�(�v�:/���Z9�9����]��o��@�R���=a���v��l���i]�$���𑔾ߓ��פ���~�����>�\w=�>��=g�<r'Ｊ��<i�C=��<83�<oxk�ClB<4Q7��@�:������5�<��D=q.��˾`�|?��H?��+?�C?Mo}>��>r-;���>\����:?�WT>S�Z����d<������є���ؾ?�׾��c��l��eF>l_J��\>�4>pK�=��z<�&�=;�i=ю=�h�V�=���=�k�=W��=jc�=�>��>�6w?X���
����4Q��Z罡�:?�8�>o{�=��ƾs@?��>>�2�������b��-?���?�T�?G�?Gti��d�>>��]㎽�q�=�����=2>G��=��2�W��>��J>���K��5����4�?��@��??�ዿТϿ*a/>��6>�{>>S�i 0�	�c�"�c�$ W��� ?��9��O̾���>���=ڬ߾�ƾF�5=��3>��]=�����\�MI�=�{���H=L�w=.f�>)A>�D�=?��sj�=M�D=�&�=�`M>ϔ�7<��6���+=���=@|a>o#>A��>��?�.?f|b?Vػ>�[r��¾�����>�E�=*F�>��= �H>N;�>R�9?��D?��K?��>�n=���>n��>�3��qm�����(���?�����?�O�?�q�>�aȺB=�C&�.c8��<����?�1-?��?9��>�P��޿~m��5�o���*���=�����v	�y�(=a#���@����m>���>���>��>b��>�#>1�d>4r�>�L�=�,=p.�<�鳺� B=�&�;�v�=�z��!7�=b7�p����TƽvO弄�=�ݝ�<*���F;�=ѻ�=q'�=�a�>7}>[��>�B�=վ���=�G���2a��Aּ�}�4�7�"Rc�d4���;��?�s> >�U'>ӝڽj��Ӳ?�v�<*�v>h��?�ɂ?��=��X�����H������s��v�>}�=<rn��U��X�K5l�i��y��>�
�>�J�>m�l>�,���>�yot=/�;k5� �>�A�������*q�<9��8���vi������D?y;��_f�=O�}?6�I?NΏ?9[�>�/��Rؾۘ0>,8����=A�z<p��V��3#?�'?'��>�^��D�}H̾4���޷>�@I�>�O���J�0����ͷ���>������оe$3��g�������B��Lr�V��>�O?��?E:b��W��UO����%(���q?�|g?E�>�J?�@?)&��z�r��0w�=��n?���?F=�?g>��@=��b����>�7?░?Qz?���?��8���>%D=W_&>��Z�pX>�I>�1>�>��?r?��>Ph@=d�7�/�JP��C&-���=mㅽO��>u�>Q,�>�ć<'ʌ=� ;=.`�>�P�>�H>c�>�C`>�=>�ᘾ9���(?,�L>$ت>�lF?��u>��
�Pͽ�ּf�û��`��94��h��i�<�<X-P;i�<"����>����PҔ?�B<>ʤ��?[�羾��{�r>4>�綽P�>��>=͠>�|�>$�d>��>�:d>Ю:>�)��~X�=�����Un�ΎL�y8��Tm�>>�	�΅�����7u=/HN��к���龳�s��Ԁ�w��HZѽh��?e�վb�_��O�_�<k(?B�0>��X?�����Չ�Q��<t>���>"Ҿ�4��6���c��ֱb?>��?�;c>��>I�W?�?��1��3��uZ�.�u��(A�8e�<�`��፿����
������_?��x?yA?rR�<�9z>Y��?��%�cӏ��)�>�/�9';��?<=:+�>�)��f�`���Ӿn�þ�8�=HF>[�o?"%�?\Y?�SV�_̽ݚ&>"�?S"?��m?��8?):z?�����?�6>_��>e�>/�,?�4=?0?G�J>��<>(��9���<�.��o����i�zŻ;�H��Jr>^w=���E�^<0N>��S!��U�耉=�K<+�=�>q�=��>��_?���>|�p>*�,?Z1���:�X����<?��=�f��������Cݾ�>�n?*�?��V?\�W>vM��4���>��r>��'>(Qo>�3�>�˾�;p�ܱ�;�>�C>���=�6����:,�����r��<��8>lS�>� |>���ER*>�����J{��f>��R��*����S��RG���0�X�w�bw�>��K?�K?�d�=��辊��=f�?�(?��<?�HM?p�?�z�=,۾w�9�VqJ�\����>�-�<@��������s�:����8�Qs>3����~�ZR�>�<�nO���K��&U�xͶ�gؽ�������v�	�gj�����j�=�m>Dh־�@5�\쁿"���22:?�������(XC��&˾])�=���>�s�>�� �|3P�h�9���{�F>�D�>#S�>Z[�'�Ծ+NH�א��ύ>_�Q?Jf?�6�?�"��ɸ���������@�㾭�n�A=$?��>a��>7q>�c>WѾ�f�gȄ��9o��>/~�>���B�;�Z���(�ľ%�a�c�=*'?��>W�+?��?H�?�q?�CD?��?=֎>��B>+����0?2�?x��=
��cՎ�'NZ��2����'?b�*?�A=?:x?�� ?�Q'?�Aj?�$?���=�X����w���>]�>��_������>A ]?�e�> u?��?��>zt4������i	=1m����=,�l?
�A?�@?�>�'�>�~�F��=���>~K}?ǲr?�dm?g�i�� ?W�>e��>�>[�> �>L"?8TD?Ӽm?�x/?~g�>乫;�Ħ��������.�<�5�7,�?�=Y�G�T�-��+�8Oo��d=*@���~r<�)���L0�����"A�>Ft>T�����0>G*žTq���3@>{����������:�#�=�$�>�?߰�>�f#��>�=v��>��>����
(?��?�G?!��:1tb��ھ�L���>��A?N��=�m��|���u�.Jj=�m?�]^?��W�@����b?T�]?�`��=���þP�b���K�O?-�
?��G���>z�~?��q?u��>�f�M<n�����Db���j��Ͷ=q�>�Y�+�d��=�>��7?GP�>u�b>/"�=N|۾R�w��q���?��?��?���?(4*>��n�m4��/�2����c?���>5Az�)??R�=�Ҿ�`��R������܌˾f���QЩ�Rɲ��@K�˛W����M_=�t?�d?4�w?�yK?A�8h��T���{��.^����\��0�-� �6��&V��z^�����P(ƾ�P��"N��E3��~�?�>8?��I�b�>'c<[��ƾ��>�M��5셾[?�>(��<��ͼ��I>�v��OZ�}�z�2� ?�dy>p��> �X?�3?�c�D��׭"��K�V��>%�a>�2>��?%J>��e���žM~��� ���q>�dm?$NN?t4m?j�C��
4��z�,
��������!��=�5����H>����`L�@=F�b�I�@������÷���Gھ(2(=�O?9�>9���݋�?+g-?�i.�G�v{B�g�Z����2?۪�?��	?O¯>w�l��xT���>�oo?D�?n�q>"y��i\�Q(��jY9�N��>-��>x��>eT>>W
�9�l�Ֆ�D^��t�R�=�=oi?8�o���M�g�>�rb?����5i�5��>�Ж<��� ���u$��]>��>A`�=�>:5���վ�O���̾h�1?�(?�_}��95��>�M?�>��>�?�>���V�>��??I�V?��P?V�<?ƽ?�:j�0��>��0����&=w�>]��>?c�<�/�=�����f��В��o;�֣�>!�����=�P>~r�L�e=��3��>�vڿ!8I��߾�����㾜e�􊉾-��� Af��K��о�<��|�}�"q���*��?��b�j���B�x����?���?����r���W��a}������Z�>��P�Ioڽ3Ǻ�x!������d�׾�Ƿ�̳$�}bO�J]��.b�f�O?1�"�{�ҿ��w�Iʾ�a?��$?���?D�;���:��6�N�H>�&��,�=�����颿�ѿ�8���g?�w�>ת"���r��>�"*?��>N�>
S��T߾o�!>�p?SL
?�!�>�l��CտLy���=��?Sv@	h??�a(�+�����=i��>$?)l�>�2�j�"�M�����>v��?�ݎ?�=��X�k�_;�c?��w:��>�ȩy;"��=��=�==i�g�6>�L�>���jCo��Ua�R�7>D��>����v'۽N<r�б=Y7Z>TT̽��w�5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=L� �2A¿��&�z�-�yid=4<�������нc�r�B�<�Pʾ�q�����wQ=^��=�Ђ>�]y>��>*�$>�3a?��?�p�>ҵE=�dL�Ѷ���;�H=]*��W�(�����߽�O��D��y������W
	���ž��5��V8>�]\�8�������Z�A���'?%q�>	���H���+�>�8�����phM��҅�
q�`��^����?M�G?I1��F��D��G[��Vp2��� ?p8�� ���b��7�>�W���=�a��>������'dƾT���-?|*?0'ɾ�ґ��>����}˻�'?a?��;�ӈ>��0?��������ŀ>�7>��>q �>`��=l���c����?�w\?H�y��� �>�?оךs�#�?==�>S3U�����hu>'l=�܉�o׀����|<"X?���>�Q$��!�e���{��9W�<�.~?$,	?_x�>�c?!�D?��= +�&�F�������=ԦU?_�^?]��=�Ɋ��}̾MZ��؊3?�
e?��^>g�w��v羽�4�I-�f&?�n?�b?�м"����2��ٝ��T=?0�?�]����=�jࣾ�g�>&��><	?�aR���>��~?����ls����ſ9�@��8�?9�@�6@��>��-��.�>��@?�6�>!B��Ὰ��>b��Z�V>:�?�F��<k��y�4����4%?e��?�?X�Q��s'�@J�=��9��?"�~?"ۉ�Ϙ>M��?k�(����PB&>���-F���+�P-;��D������;0YýWŃ>�@J̽�E�>~�{�(M�TiͿ����Pݾ���n�> ��>���Y�վ�Cj�'o�o\�|�A��KV�O��>�K�=Oޖ��W���s�R�<��z�=;5�>�t����>�]������ck��>t=�!�>4��>j�>ɤؽWZ��Ơ�? �M#ȿ�ѓ����#O?=�?徆?|� ?l'�=%n��8�=��J?�|a?�U?��@��S��_��I�k?�J��J�a��?3��A���V>�2?�N�>��.��{=�X">�=�>Q>	�.�J6Ŀ�������?C��?��v��>`��?,�(?`��_���������'�I�ۺz�@?H.B>��¾�%%�dA��j��	8?�4?�+����Y�_?(�a�E�p���-�k�ƽ�ۡ>��0�f\��N��գ��Xe����@y����?G^�?j�?ɵ�� #�g6%?"�>f����8Ǿ��<���>�(�>.*N>ZH_�a�u>����:��h	>���?�~�?Fj?���������U>�}?b��>�ӄ?��=\��>9��=*{���W@���>/��=M�E�6?Y1M?��>j�=A6�A�.�U�F�-{Q�K��G)C����>KOa?��L?�y^>l���.!�$�!�!iɽ��0��
��A���,��#ٽ�?7>s�:>P>0LF�UcԾ�@?�T��UٿЊw�x=��9?��>x��>�#�վ���L=��A?�6�>ڷ������4���L�mպ?l��?C�>"�I�k9�=�g�<��a>��L=;���m(;eBE��t>�w?��e����������R>W�?Q�@m��?�e�z?d�	�B ����z������(�V��=�8?xN��#u>�N?�t�=�	u�iê�lt����>���?A��?��>i�c?�`�X�3�2��<�y}>��e?i?7�D<��ŐF>?�������
��Nc?U@�@B]?q9��p9ܿ�z��]������%�79����d>Kﳽ�� =��=A�q�0:�'F">���>o�>r�>��>9�=�k
>&������奔=|��4?���#�n�����g�m�侔!p��w׾廵���>��� �>n�=SQ�	K�y��:���=3�U?�R?%p?�~ ?_w{���>,S���Y=�#��Ȅ=pچ>[L2?�L?��*?ǎ�=ˢ�� e��`��P/��ɇ����>��I>X�>a�>JA�>��8ȔI>s�?>V��>d� >�d'=5����+=1O>6F�>��>�J�>�Q>��>攷�!˥��s�NM��Yu���?�?�����"Y��A��y�f�')��Պ�=�C0?��=Z=��Hɿ|]���T?ՑɾL���@�	��=�<C?DLM?,�>p�־f�m���>�1�H�[�|�=���⁾�d*��rT>+�?��b>&�z>;��22���V��h���g>�,?�����D��do���@�(澫c@>�[�>Ù����!�iO���4�p�b��ki=�5?�7	?;��	��VO����X>��[>*� =�Z=UY>>l��lɐ��U���=�[�=��7>�v?(>D�=�̢>�D���3M����>��=>�6>.�@?p$?�����&��M"*�@'~>D�>6�{>��>.�B����=Ly�>��m>��_ɖ��#��kB��(J>�G��tl�R��k��=�������=q�=o����?�w0=�~?ƈ���숿3�꾬����D?R.?��=~�=<�"�����D'����?3�@GU�?\�	���V�b�?eP�?h����t�=�v�>�ϫ>��;A�L�_�?�ƽﯢ��	���"��A�?�
�?V�/��ϋ��l���>�u%?�oӾ�j�>׀�[�����a�u���#=���>U<H?�W����O�E>�Lv
?w?�]�"���t�ȿn}v����>q�?���?U�m��@���@����>ߣ�?fY?�ni>Al۾KXZ���>9�@?�R?��>�:��'���?�޶?J��?�1f>�:�?�x�?��=��9�����!���M��v�ν����D,�J�s�9@ľ��z�sɦ������G��[9ƾ��?��p<r�>�߭�ĉ�공��p=������b%�>ce�>��%>D�@>���>�C�>-�O>T)ͽX�t��J�� ���K?��?	��Gn�Z��<���=*'_��.?�i4?�iW��Gо/��>��\?k?�[?Az�>�z��*������3����+�<k L>��>Qy�>�܉���J>�վ�C���>�{�>7o���vھt���>����'�>L!?�K�>i�=�� ?�#?�j>�'�>%aE�r9����E�'��>
��>�H?��~?t�?AԹ�[3����硿�[��9N>��x?�U?9ʕ>P���>���yE�GCI�6���:��?Mtg?W��?2�?��??ߤA?i*f>g���ؾȯ��b�>l@!?�����B��~%�Q�Q?�<?���>I�����ٽ?�׼2�������'?"�[?�&%?�(��`�Jľ�A�<R�(���B�+�U<�u��>�u>R���}D�=�c>K��=��p��6���<#��=x|�>�Y�=��8�eZ���/?��!�K2O�~k=����1I���A>��a>�͸�)Kj?[kW��y��˿>��m���7��?���?��?`d�)Kp��N?i�?�C?���>l�Ҿ��޾��̾hlY�f��n=����=W��>�u==�Kﾻ�����ᕿS;3��"���?X��>�?��?��>�*�>D���D���	�p�־*g~����8�(�^I��}�RD��T������Ę��p�>ɦj�1��>!3?¶V>D��=X��>-��;�_�>�>�i�>��>?��>S)C>��>4��=��� LR?o�����'�q��ޯ��83B?�nd?/�>{;i�Љ�����?Ճ�?�q�?�2v>�h��.+�uo?�C�>���
n
?sL:=bf�lC�<~W����S^���
����>�1׽�!:��M��gf��f
??,?���ق̾�/׽k&��v.�=þ�?c�$?^3���3��e��1]�o��Ȇ����}i���)�R����C���܆�iS��x�6�R�Y=t ?�0�?�-
��RѾ
���~�{��f�B�'>|I�>5�>�[(>F��>�����(�a�ʐ���x��#?���?oj�>��7?S�E?ޠa?F�B?�$C>w�6>�1����?��=��=�60?e�<?G2b?IW?��)?0A?{�>y�?����Ͼ�6?�5?h�?�\�>YG?S7�Eo�,ݔ<��^>����.�v��=ɴ���ݗ� Cý���=��>Z^?C����8������k>�7?]��>X��>�%��p5���R�<}�>�
?WT�>t �C�r��h��c�>!��?����[=x�)>�=�=���U��N�=�pü/��=�CD;�V�<pÿ=���=���ӎ�+;D͍;�L�<�t�>>�?ē�>�C�>�@��-� �t��ae�=�Y>$S>(>�Eپ�}���$��}�g�u]y>�w�?�z�?¼f=��=��=�|���U�����.���g��<�?@J#?*XT?W��?a�=?Yj#?��>+�gM���^�������?� ,?���>����ʾ[�6�3�E�?BZ?�;a���~:)��¾�Խe�>rZ/�k-~����D��f��z������Κ�?�?�,A���6��r辗���a\���C?Z!�>�U�>��>?�)�K�g��$��0;>��>�	R?�!�>�O?�;{?�[?7{T>��8��-��/ԙ��2���!>@?�?*�?My?�x�>��>��)���fM��������삾l W=FZ>���>o'�>�>���=��ǽ_R����>��J�=C|b>v��>���>/��>�w>�R�<p�J?Y��>y����o��_��(���|J��F?��?�V8?�v=���0�+�ݘ辳 �>�֪?�ߨ?!-?Rfw����=����ݛ��Et|�po�>���>��>��+=$=k��=��>�>].�����7B<��諒��?,47?�<>z�ſ��p�r�s��;��l�A<4_��2�e�g���X����=�
���w��?��*�[�П�*)���t���7���}����>�T�=2�=���=�w�<@�ʼ�o�<C=8L�<tP=��n���M<��>��Ȼr�����_���N<9�D=�8�)�˾��}?Y9I?ד+?�C?��y>�C>��3�t��>�����>?V>�]P��|���~;�Y������ͳؾOv׾��c�ɟ��I>�{I�W�>H=3>�P�=]D�<�(�=��r=)ǎ=V�S��=34�=^V�=�_�=ʻ�=��>{I>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��4>B8>FRY��(.��z���n���h��?�s2�U�Ҿ*��>U��=)�jƾ��S=r�(>A�<�]�Lm[��8�=p���1=���=�_>�@>88�=����L�=*�m=�3�=��>i�ϼ����ȅ���<��=U�N>�>?��>�o?�80?LPe?���>1�l���̾ þ5G�>1��=PJ�>�4�=5�C>u(�>�$8?��D?X�K?�˱>Yh�=�ٺ>d�>�-�fWm�B���X����<Q�?�#�?H�>��Z<O�A����9w>�@vƽ�'?0�/?��?aq�>����^ؿY�4tR�3���gID�$�=��z�'�<P�=(�/��?�Q$�=J�>&��>%l�>���>�M�=�?�=q��>�$>��F��m�;U\�=p��=;E��w=��=�FP=�p�a�m=�\�( ��!���ν̼�<�ej��ѹ�� >���>L�>$�>p�}�{���v&>��/�c�]LS<w&��GR�]�|�x���_O���*�Ei>��Z>�?��54��Ʌ?���={b>7��?`�?�>�)ü��
��	��?1x�N����>��>�0u� kG�*U���b�踾v��>^�>��>��l>�,��?��uw=	�`_5��>z��B��r%�J;q�@������;i��PںG�D?�D��p��=n~?'�I?$��?$��>`����ؾ�70>�Q��J�=���(q��U���?�'?���>V"��D�}H̾����޷>�@I�-�O���Z�0�*��ͷ� ��>������оk$3��g�������B�Mr�V��>�O?��?]:b��W��UO����8(���q?�|g?�>�J?�@?�&��#z�r��9w�=��n?���?C=�?_>��=�T���r�>��?.�?X��?>^p?��r�	l�>b� =��(>��n��d�=S�/>V��=��>�?%�?1�	?w�������r-���A�� �<&��=��>闂>Hcu>m��=�=<iI=�)>�]�>qDr>H�3>�؝>u��>�ړ�B���+!?�?D>���>��e?��> \=�#�R���Kz>ĚȾ���>��_�m�a��<�"�=�0�=b	�<ʤ�>�&ʿ���?��!>�F��K+?��ݾT�*��R`>��=�?l<(��>v�D>7J�=��>�>�SI>Vj�=���=cد��A�=Mh"�|��W��O��˭��D�>����F����%��p������IھO�m��߄�.�?�!!ɽ��?]����f��A0�֋˽�%?û�>?<[?�����3��� >��>��>F���'��!L���l��?y3�?�;c>��>I�W?�?ƒ1�.3�vZ�+�u�s(A�1e�N�`��፿����
�����_?�x?&yA?yS�<-:z>R��?��%�\ӏ��)�>�/�.';��?<=�+�>*��Q�`�u�Ӿ��þ�7��HF>��o?9%�?{Y?TV������=�?2?`��?��.?�>?��ʾ�YD?�x�>2L?`1�>�*?��"?��?���>O��>�~b���F=�ս��Y�i}ֽ��~����!S=��>o�=r��=&z�<If�<h���*oc��� �������;��<��<K�=Mצ>6�]?�@�>�Ɇ>��7?/&��7�m����.?s�B=ߑ�������ѡ��^�i�>vk?��?�6Z?�od>ҍA�T,C�R�>R��>�i&>��[>�α>��N�F��S�=�>1�>�ߦ=A�I�;��1�	�N`��b�<�>��>/|>@��1�'>)z���1z�U�d>+�Q�Vʺ���S��G�w�1�)zv��[�>i�K?��?���=�^龴'���Gf�n.)?s]<?�PM?�?��=$�۾9�9���J��1���>�(�<��������#��D�:���:��s>F0�������O^>���#�̻l�tT��㾄��=+���1{<e/��}ž�B����=�>A����'$�����(���zK?�C=�M��qY	��*Ǿ!U>��>"K�>E+��k���3�.�����\=�=�>�C>}b¼꾔sG�w��{q><�G?֣_?n�?���tk��<!�x?�\Ǿ����L>�>�ؙ>uq�>�(弆�s>�S�TQ&��Ȍ�Vt'����>�o�>����E�E���]�޾AO9��č>�tM?���l�>�֒?$��>:�K?w�1?�3?O�F>+���͹���Y&?,o�?Ԋ�=:Yӽ��U�?J9�_$F����>�)?�'B��j�>��?��?��&?vtQ?}f?��
>�y@��d�>lT�>�-X�[_����^>��J?-*�>wY?F߃?U^@>5��n���v�����=�>�p3?�#?Ƚ?<{�>Ή�>'���~�=��>�c?�.�?c�o?s��=�?�52>���>�R�=���>��>�?�XO?��s?R�J?\��>�<xZ������us�\O����;�H<��y=�L��s�,\�*N�<��;d��6x���򼏫E�g���O�;td�>H�}>�����5>����b��	)E>��#�������u�"�_C�=<�>)?w��>`�[=⩼>Ŏ�>����"'?$u	?YH?X�;�c�(�Ѿ�k����>��??u��='n�����
�o��BU=�,m?1`?��X�w�[c?D�[?P���)8��	ɾ�y{��쾀�T?��?��<�k�>��?q?�\�>�9T���i��Ĝ��e��8n�'�=)��>�P���f��/�>l�6?���>�/c>�g�=�|þŲw��Þ�Y�?��?ܭ?^L�?�->�f��G߿i9�f|���lk?d�>�k��3@?�G;�Ծi�P�����OپC[��DȾeS���ȑ�<c!��jx�!�&*7�X ?��k?+�c?�E??)����n��>:���~�z�l�%��O����5�*eA�T�5����X"�4���ȾuR�<4uw��F��5�?V�)?2�@��w?!������%���=>sޠ�Ĩ��Z=�ݣ��Hu=8�m=�Z�I�4��.���j?��>/��>�u/?�([��^=��i)�8;�<;����>pj�>�n�>;�>~����tE�����۾�|��@򽅫W>ei`?w�K?>�w?B�M�
-�s5f�:���R�W���I�k�~>l�a�P�>G�?���]���C�>�B�vdx�k྾�/�����=n�H?S��>���=D�?J�4?]����#J��y��Ɣ=��N>�	�?E��>b�k>�8���B�:d�>��h?��?��^>e꺾���m��(�C���>3��>���>G��=����v@�����(����=��a�=8�?r�g���a�WJ>�s?�5���ͽ�y?G�>
�"�xq��"N<m�=:�"?)�=Ꝛ>Cþj��ͨ���Ɛ��"L?�.�>gH��7;����=t?%j�>�c�>a��?x?L���w�8>�H9?0�w?,GV?�Z?~2�>}kH���Y�T��$����?>��>�4>�ڈ��F�ڤ��&�S5Q>0'�=�\�T��������֨>@\R>_�\>�{߿HK�t��/j1��Ѿ��h���Z���<Xf��P�"���`]��lD��~�8����E��T�&_j�%v��*�?�"�?�����&�������������E��>(j4���ݽ����׽��ԾOn�xn������Q�� S�߶i��&?�0����ǿğ����3�?�8?~y?;
�F<$���3�P�>�8�<�!ļ��������οSǘ���^?���>��� ��=c�>�O�>�_>��f>����柾:�=N?��,?���>���Nɿ[ź�^��<���?=@փA?.�(�`��8�U=E��>]�	?4�?>o*1�H:��װ�FX�>�;�?���?#�M=-�W�k�	��{e?x�<�F��g߻�P�=�\�=7"=�����J>�A�>�K�(A�>hܽf�4>ׅ>�-#�#���u^�2��<��]>fս�m��:̄?E|\���e���/��u��:�>�T?���>��=�t,?�8H�,�Ͽ7/]��`?��?w��?��)??�����>�#ݾ��M?g6?P�>��%��u��N�=�����э�$�V��U�=p��>|>�X,����7vP��m��J�=���ſc"�w�-��`T=.I���n��c�^��V���3��Z�M�����S�=[B�=��a>�`�>�N>��L>�a?
r?��>s��=�Z���6��D̾� ==�h�5��N���! �̼��b@���ZѾE1���l
�uhҾ"F�;�=[�Z�����tO�����l5���.?��Y>������l�Nv�=c�۾R<��2�|<��<���ྜྷ����s���?��D?hS��$!�x)�^$
��"��/R?ؙ���_�%�j�)w�=��y�"L�<�>L�s<����4��a��l=?H�,?@߾����E?>�)����H<�qP?���>��)>�?�E?��<���=.��>�,<>ϯ�>`U�>Q�I=�پ�s�� �5?��t?��Y���<�>��������f��@!>e��&q���p@>dO�=O���N�=������= EW?���>�*�(1�C��e���?;=X�x?=�?�ߠ>�mk?�C?v�<����S� �
�Y�x=�W?��h?8:>�4���Ͼ�{��z�5?[�e?3WM>�g��Q�Y�.�R��-?�|n?�7?�Ο���}�V���&��W6?��}?�v��������["�.��>�>C�?Q�N�,/�>��l??V5�����(Ŀl$"�_�?��@}��?rߣ;�䎽}��=���>
��>�;���n�����&��H�<*��>|������8Q��L��t/F?��?�?�:��Ȉ����=Kɣ�B�? �?��eڎ=t��a@i���6BϽF��=uT^�E��������:��x־����̾�۽ip>�8@�r��R�>)Q'�9俸�����m�+O���Ǿ�?�ŉ>CU��h���Z�~���z�մL��uR�?*��2�>xf>�������Μ~�G�L��� ��?�=>hK�>���Z罓|��tC.>��>�C�>N8�=dr��yᾌ,�?)��A�ο2������b\?���?�[?D�)?X!�>��������_:�>qЂ?�n?��?��=ϮȽ��N��j?�a���U`�d�4�oFE�OU>_"3?fB�>G�-��|=�>��>�f>$/��Ŀ5ٶ����s��?��?2o����>w��?�r+?�h��7���Z��8�*�A%-�d<A?N2>݌����!��/=��В�`�
?y0?�x��.�`�_?)�a�L�p���-���ƽ�ۡ>��0��e\�M������Xe�	���@y����?M^�?i�?ڵ�� #�_6%?�>e����8ǾJ�<���>�(�>
*N>�H_���u>����:�i	>���?�~�?Oj?���������U>�}?���>F�?J2�=P�>�d�=摱��g�n%>���=��5��j?q�M?���>�=Έ5��z.�|E�({Q�S���D�_�>��b?M?�Zb>B���$&��S"���̽�1�n��YC���+��'ڽ"�3>q?>�'>�#E��Ѿ`E?�0f�tӿ��q��3%>Z�?U?6>R@�><����dw���q���Z?��>.��f���P��SP����?�f @���>�6�ml>�
�=��?�%>$˃��EN=�d����>7�,?�eJ��v�!�F��N�>D�?�&@�ȡ?7Y��[?��(�z<���gf������S8��_�=tbB?��ݾ.}�>?H�>!�j�4���j�d�F�>�Ա?���?�y
?	WL?��K���"�e�����>Ii?��>��>cn�LQ�=h6$?N�n��<��i�R?U	@fC@�kb?�筿ۿῐ>�����߀Ҿm?�=ڥh=u�'>6����=s�<�c���=�N>��>�i\>�t>GD>}�6>6vI>[����r��a��L�����7���'
���8�ɿ����[�=��a���jr��1�RO���Z�dQ�n���H�=�U?�R?zp?�� ?�;y�~
 >����_"=�A#�`Q�=j#�>Lk2?t�L?;�*?f�=���U�d�*W���=��������>9KI>u�>I�>;!�>KLy8��I>�?>�{�>.&>@�'=~F���
=��N>�G�>���>8c�>�Q.>3�>����� ���h�5����Pͽ�{�?挾K��ᕿW�|�"5��(��=��-?��>�M����˿
�����G?��������5½5��=�/?��O?"z>^���W�W��J+>'���Lh��>�㽡�e�0"���6>�<?��1>LK>��A�g,$��#`��i���P?>�^7?�[y�G+��k.n�С(����|�6>}L�>�\׻$��玿<�����'���<W�)?�[-?�����`� l<����5�e>lG>R>k	?<�z>��h;DU���W�{[�<���=�I�>I[?p->҆�=� �>���8�Q�h��>�}C>�;*>\@?&�%?���*y��v����+��Hw>~�>;�>6�>mDL���=���>�?d>�/�8ֆ�/��=�D��hW>�-~�<=`�R-~�j�x=W��DB�=�;�=����r =��s*=�~?���'䈿��Ie���lD?Z+?� �=��F<��"�E ���H��G�?q�@m�?��	�ޢV�7�?�@�?��=��=�|�>�֫>�ξ�L��?�Ž1Ǣ���	�)#�fS�?��?��/�Wʋ�3l��6>�^%?��Ӿ[��>�DY�'�����a���n���=:'�>�7?gN��㨽)� G�>���>����T��PLĿ1n��g`�>�g�?�m�?�������(U6�W�#?H��?�n7?޵=��Ӿ��2=��>��??�}S?Z;;>�)�B��!?�S�?ls�?���=8`�?B�?��(>��#���ֶѿG?������&=Խ�I=:�2�q�߾�0�zn��_����Y��߆��?�v9=-��>N	l�_� ��#A=��=�禾2潂_�>�
?״�<��>���>���>?kQ>ߥ�ġ2��V=�l����Q?�B�?z�r��Չ<���==a�U�
?��8?��k=�����v�>(Ma?C�?�Z?�0�>>���+��*B��%���.a=��7>P��>RY�>l;J��8>� þ��o�Iuq>wN�>�T#;�sj�����q҃>5�?2��>6�=K ?��#?�k>s�>�OE��Y���(F����>}�>0b?h�}?F�?�
��� 3�"��	���?�[�/F>K"x?�?�֓>�ҏ�m���Cb�9yF�����M�?�yh?�~ݽ�?�U�?��??lD?��c>o��C+׾�Y��N>%�$?����"A���%�ѹ��?+9
?��>�>�ę��h'�t���뾵q?�P^?)?|m�>�a�K�Ⱦ���<��_�꒼\�-�GD��R->��>�m��3z�=!U&>!�=vo��2���]<K��=�ۖ>/'�=�",�9{����)?�׽Y&��6/��}�v���=�p�<>��	>9 Ѿ�7?2���� ��s������89I��Ȕ?sQ�?�a�?��%���o���O?���?X??x�?
��?.�<��VA���&���r��>y>��?�e���9�ڲ�����6���s�̽0)U��Q?|�>8��>6?	��>w�>�˾)�E�E���:���A�n���KHG��8��1��Ƌ���E����-���\Z��>P�=Kr�>��?���>�\�>�`�>���=�g�>8>E�>%�>&�P>fH1>]�>�x�<ߏ��&LR?`���,�'�Ƿ�Ӳ��83B?�qd?�1�>i�ɉ�������?���?]s�?x>v>b~h��,+�9n?�=�>C��=q
?S:=�5�3>�<�U��ݼ�04��O�몎>�B׽� :�|M�*nf�Rj
?p/?v
����̾U:׽�����4�=���?�/B?:C+�rB��S`�J?���W�M���C �#��w�5�5�g�����(���LM���I�_�=�V?���?�~����b����S���m�ǭ8>���>�^>��>ʭ�=&ξ�.��Zd����FBi��?�-�?�E>Ҽf?�g4?��O?w�J?��>���>�b�����>
f�=���>1g�>�D?�-c?�C?�?��F?���>�t����~u����J?��>�E?��?�&?��f>�I�Iq��L�g
x�LB�=eL<0�3:�v%=�=ġA>0Y?J��K�8�	����k>�7?�~�>��>R��o,�� �<-�>r�
?rE�>�  �w}r��b�zW�>���?��b�=��)>���=t����Һ�\�=	���"�=:���f;��\<��=���=Rt���}�-��:I�;Tq�<�t�>E�?��>jC�>�@���� �����d�=?Y>KS>�>%Fپ�}���$����g��\y>�w�?�z�?��f=��=���=}���U�����������<ݣ?"J#?*XT?F��?Z�=?Qj#?�>�*�cM���^�������?C!,?B��>�����ʾ���3���?�[?;<a����:)�	�¾��Խ��>[/��.~�m���D�������z~����?���?xA�"�6��w�����M[����C?�!�>�W�>h�>��)�J�g�%�c2;>���>{R?�#�>��O?�<{?��[?sgT>L�8��1���ә��I3�>�!>@?ⱁ?��??y?*t�>��>a�)���$T�������Ⴞ*
W=,	Z>k��>�(�>)�>��= Ƚ[����>��`�=��b>Y��>���>��>ޅw>)M�<�YU?~_�>�оG������J�b.�d>v?�ݕ?�9F?�|�<=��������r�>5ڪ?N�?��?it����=��4=h�¾�Ď�T8�>���>�z�=�H�=�Լ>�>���>!��>I�>����!�<��d½$�?��N?< �=��ĿAp��w�b�����;L��5d����e$S�+o�=�5�����}W���Y�2A���������d1�����iO�>i�=N�=�6�=j��<y5��c�<@AC=%��<�=��O�H2<X�(�[���L����!⻸<niQ=��:/�˾yu}?�*H?�++?�gD?{�}>)j>�A�ۊ�>�h��	�?^�P>j�R�0ս�`�=��F���o��ɧؾHrؾ��c�c柾��>��4���>�5>j��=k�<Խ�=N�=z�=�v��)=]y�=�ʽ=�=��=�>��>�	y?8󄿅����Z��7t�=�>?��u>h�>�վ7Q'?E҃>�đ�N�ǿ���L�w?�=�?��?(? �����o>'gA�i�c�L-�=�U�/9 =�y�=i���8o�>	'<>BJ��ۧ�U=�'�?��?��1?5n|�~ο-^�=\b$>]��=��U�b!�a,�������S��o ?��'��a��s>l6�=i	�R����9c=�+>�4<�&�8u_��l�=%u��?.=�*�=�G}>e>fK�=���c8�=�|�<�n">ʤ->�_�</��������<X�x=�r>5�c>Ò�>f�?�a0?;Xd?6�>in��Ͼ?���I�>�=	F�>>�=lsB>T��>n�7?��D?��K?х�>���=I	�>�>S�,� �m��l�5̧���<���?�Ά?Ҹ>"�Q<l�A�����g>�50Ž�v?SS1?�k?��>�r��߿�"�A�;���+���V�K8=�C���4K�^��n�R�������>ޭ>��>�O�>q�o>](>��G>mN�>qN.>k�(�-;�;W�H�&��lر��>P�r��h;�ذ�mǦ<F^�`o{�h޻�u�<}a��a�<n���E��=���>�?�=䴨>*�>BՈ�h�=�d���q���/�}#���xN���`�Ө��tE*�ߥ$�*�o>�(>�7��w����?_>[TG>>��?܇??L>�\� �t�����<����t>� �<�M����J����xX��d׾�S�> ��>x��>hSs>�n,�j�>�;tx=σ޾��6���>Z����=K�Fd�c�o��⤿�w��Qi�?_�ĨD?�~���7�=�|??7K?-L�?��>(�~���ξB�&>lZ��a=�L� �j�gy���?�'?9��>�0�B�F�5<̾V���ѷ>�1I�L�O�m����0�����Ʒ���>P�'�о!3�Zg�������B�scr�l�>a�O?v�?�Pb��R���UO�U��� ���h?�og?��>0U?6?���h�q��+r�=��n?y��?�>�?�%>^`�=J���0E�>�)	?���?��?��s?ֺ?��|�>��;�� >r������=�>+ǜ=_\�=�v?��
?��
?w����	�-����C^�qq�<�ϡ=ă�>�t�>�r>���=�g=R`�=x\>՞>��>�d>b �>�K�>���V���Bt?��>ʰ>�so?fi>N�<*瓽���.=>;���\�X�ůQ�iW��A�=��
>�r��2s!����>(�Ͽȕ�?/̀>��7�9!
?�_��vt>�"�>g�E>�|��g?P �=��>�?�ۜ>h�>��V>�w>Rư�z�=��+�{�ݾ&�]�4�F�#����>��ܽWþb���5����Tp��x��0����b����<#�Lв<�t�?�8�2(w����ӂ�X� ?usX>r)?[���o5�<@݆>^z�>���>�o�%���Z����n���?�[�?m9c>�>��W?H�?��1�*3�qxZ��u��'A��e���`�8፿����~�
� ���_?�x?�wA?|��<�8z>���?��%��֏�*�>!/��';�r1<=�*�>\"����`���Ӿ�þ3�IF>E�o?�$�?c\?�NV�o���mO�>�Q?��?��?�c�>�ڃ?b����?%�>g��=��?rL?��b?�8?34�>�'>�ޔ<��<Kӥ�4׷��^��ǽ���r&+���=�u�=o b�;�>�K=�e��|�<L�㽊��h'������i]���;�>�]?�R�>Ė�>��7?����r8�IҮ�*/?��9='������o�������>1�j?k��?�cZ?med>{�A��C��&>jM�>�t&>7!\>Qb�>�|ｋ�E�-�=�>>_`>���=��M��́�	�	�����\�<n">4�>��{>䎽��&>و���z��jd>Q�ݐ���R���G��1� v��T�>
�K??4"�=�1� ��Gf�eO)?37<?uM?��?�_�=<Sܾ��9���J�����`�>�ͯ<���񴢿,)����:��43:�s>����<���Gu>.4
�N�Ǿ1iw�aX��5쾼p'=3� �;o,�[���,������=�s>��ɾ8�!�W��<��gyC?j-9=�e���F��p���>u�>0@�>����񑽯�<�����3ه=�$�>��>~�p��4���%G��V羨��>ԕ8?i?|�?�Ȝ��t��i�]�_�������]H����?�$�=X?��Y�Cdx=	�-�3�/t���G�a�?��>u���<�����H�#�S�f���>�Cc?�˭>8��>&�?]�7?�@?(�5?x?��x>�w�<�>n���4?Jt?���=w�^�|��:�^����$�	?W�c?��7�87>�D!?�4?l�`?��[??�v>���'��@@��%�>g�:>$l��H��5n4=r?L��>r�,?�a?,�?/9����&��\�>�>�D?'�4?[�?��w>:%?}i�EF���q�>km>?Z��?��u?d"�a?l��>U\Y?�|�>�>�w?���>^�C?��K?�<?�MX>�\-���s=�{9��̽��q��6����2�<�s�x6�}�޽9�&�M ݽ�΍�� 	='�< �ݼH�[<3>F��>G�y>�H���@,>oǾ���/=>	h����y���d7�(U�=.�>�?d��>��"�R�=;�>u��>����&?[�?��?��h�V�b�+c׾V�]��Z�>@??w��=;7l��W���s�$ف=�!k?f�]?@Z����f�b?;-]?~�쾙x9�V~ž�~�0�����O?�q?� F����>��?�s?RX�>��W��k������lc�/�n�S��=�q�>Y�C�k��>N�7?<D�>~�Y>�I�=n�ʾ��w����	?���?��? C�?=�,>m�l�E�ݿ�5�}�׆i?�A�>�C��2?B�>׍�N7���a��P(��񦾑�ܾ Ǿ���	��#R��WI��a��	?o�c?��p?u�L?�2���`��5^���l��_M��?�l�B-�ߛC���F�$�l��V�+��9��I��=��{��\A��;�?�(?�p,����>QR��4����Pʾp�:>����Y5�bd=|���(�5=;9`=��d�3C<��X��t�?g��>ٌ�>��9?��Z���=�a�.�1&5�z����S >BΙ>���>���>Zr�O'4����0NϾ+F��Q����->�Y?)�^?d9l?���m�wm�s����K�G?�J�^>�B��x>T:?�[��3�I�\�L��}�#�����v�f��w=�cG?F�r>���y�?[q?�
�0�$%��[�0�n��=fA�>��M?k��>�BH>/���=�	��>4.l?[
�>Y͞>䬌���
O}�����>��>f��>W�K>��)�]Z�p������I�:�f��=U�e?�=����d����>��S?�-���t�@�>W�,�/���������=ū	?���=��4>D��G0���y�}����)?rh?~��KA.���z>�h!?ق�>5��>��?'��>�e��s`<
?e�^?H?)??z��>��l=�A����߽�,�YH=FY�>qk>�4=��=�1��Nk��8<�3L?=3�=����ý]U�<�y����;�4!=��C>Q�޿�E���ھ��)�p=پ&�	�������:��1h��7L�9����>���e.���M+��}5��`����`�X/���?���?����u־Q=��5�}��>ݾ��>��&���Nbپs��ӗ�� ��詾^��2�Y�Ub��W�+�'?Z���ݽǿҰ��<;ܾ�  ?�A ?#�y?��D�"���8��� >&A�<�,���뾲�����οF�����^?��>��1����>C��>(�X>mIq>w���螾9�<��?�-?_��>�r�"�ɿO����ä<���?6�@C?M26�x>����=)��>�G?��T>�d3�Q���j����>ø�?	�?���=�nO��J�B�`?ȯ=��G��Ui=q��=� �o\��k����z><j�>�_�OA������->���>�~��x����^���<r�Y>ʪ��ɳ��*^�?�Z�aX��4�M���Ɗ>��e?��>���=U�2?o�h��[οr1x��[?B@��?ܨ:?Ⱦj��>����k$T?��??��>~��W�e�qI=�Z��jD����E\����=���>�|F>�YZ�U�-����� �$GL=����Ŀ������宣=̰ٻ�H���޽-��s�i��颾 �a�ǫ��ݿf=���=��Y>:�y>�eq>��b>��^?�u?���>c�T=�'�#[��mPо�b^=I]R�g�O��;�����_���*־8���T��%�ٲ�y:þ��C�;��=\�X���+(���_���,��X?��>���z*b�s��=�����~�~�1�6q��h#�!���K�Kg�?\�I?����ʂ#��=�w}����͔N?�/��}پD஽� z>7�V�_<"��s�>�bv<����|���F��T-?~�@?�u��u�����>"#��[*_?��?la�=���>|�Q?'a�=Ɖ=��>7�>�\�>]? �>�������$?|�~?��4��"ĵ>r���ä�_ފ��z(>_b���E\a>'�>�;��1�l��P�@>�(W?fF�>�q)�����}��t����=�y?sI?Un�>Ij?�C?6$�<�<��'R���	����=�X?��f?�W>�?i��;�֣�J�6?f�b?C.O>
�^��V�1����?��m?\�?~����}�􅒿���C(7?5�y?�f��Ο���
���	�@f�>J�>M- ?�?�TL�>�??�$3�]������*�9i�?Z�@�e�?(��<�1Y��Qn=�>�>$�>� ��������*�t������9
�>�ѯ�Oz��D5�����!�M?��?��?������
�={����?&��?z��\w�<�  ��vo��
 �A�� t�<^�B������8�i�ɾsK����i���C�i>|�@Κݽ>7�>�.��ؿ�տ�ʀ��۾������?A��>G�����/fn�?�y���I�d�6��bV���>|�=6!q���[���h�H3!�B<�*�>�;ǲ�>�U�=���#x��F=�|�>~��>�C�>�:����¾�x�?~��0�׿����&i�v�h?�Z�?@��?G?���/����V�X,�;=�H?}�b?.eL?�6��� �s쏽(�j?�_���U`��4�MHE��U>�"3?�B�>D�-�L�|=�>���>�f>�#/�s�Ŀ�ٶ�"���^��?��?�o���>n��?fs+?�i�8���[����*� ,��<A?�2>���f�!�G0=�:Ғ�׼
?v~0?�z�.�]�_?+�a�N�p���-���ƽ�ۡ>��0��e\�N�����Xe����@y����?N^�?i�?ҵ�� #�g6%?�>c����8Ǿ��<���>�(�>*N>hH_���u>����:�i	>���?�~�?Qj?���� ����U>
�}?Р>S.�?0==w��>1�պ޾XL���I:>2R>X������>vR?� �>��k=G����,��>�iJG�M��k?����>��f?PZ?�'C>�� ��Ov���4�u,M�ڃ8�yGh�/,L���v�|�ɽ/�%>�>NW�=~���˾K^5?|�4���տ�!��5��=\?]ă>N�>�A����<���,�F?� �>}a��鬿������0�?�Y@%��>d
�LC�=W>;j�>�i>��b�1�ݼ^l��L@>��/?_�a�������t�(��>8��?�"@T�?r�y�c+?�i�ۄ��#�}�F�����[��=��6?pU����>Yn�>(��=�vt������m�o��>䟰?���?H?:�R?V�^�U'�X�	=�8\>{�c?c�?S�=~
��� >��?�9�Ԝ����5Bc?{@�1@P�W?����"hֿ����@N��S������=A��=�2>��ٽ�`�=��7=��8�C6�����=��>��d>\q>�(O>�a;>Ւ)>���1�!�Rr��<�����C������Z����Xv�Hz�H3�������=���4ýy��mQ��0&�QA`����=׬U?�R?�p?� ?�Qx���>�����=�y#�E΄=��>�`2?y�L?��*?>ד=���#�d��b���?��"և����>�I><w�>GH�>).�>��J9��I>�??>w�><>��'=1޺�=7�N>lM�>���>pz�>��;>t�>)ʴ�xA����h�#�w���̽��?�Z��ޮJ�����y��H���$��=�;.?�/>�����Ͽ.ѭ��AH?p����)�Mh)���>�[0?IW?ײ>$���R�J�>��ok��) >c����l�O)���P>b-?s�,>ї�>�s=�#S+�y�g�
b�H>�"7?�V��0�z�v�g�?��6�ݾ)>dA�>S<l��a��뉿dq���b�b�=�l<?�?%K�q�Ѿ�w�g-ܾ��s>��6>~ʣ<:c=s�>�z��iýN�x����<1�)<�F>f?�U*>�t�=ާ�>���{M��ҩ>"B>��,>7@?J�%?���Q�������#-� �w>
L�>�b�>:�>�fK�[<�=�d�>�b>������6l�&�@�~yV>���3_�E'q� Ct=�i���#�=�Ӓ=�� �>=�1o*=�~?���(䈿��e���lD?S+?_ �=(�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�-)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ��>�����.�p�	xe�v�q��>�R;?���?�a��! �Қ?���>�F޾W9��Φ̿�r���>G��?Z��?�y��Q���D�/>)?C��?]�V?s�9>���V��<Hz�>"1!?�j?��>&���G%���?饼?��?6��=J��?�/�?F��>�D�<����j��쥛��1w�D�����Q>ot��9쾎�V�q���+n�������j"�+V�>��<���>(
�X^�����MIռ7���I��Ї�>C%$>�Tu>���=2�?S��>y�l>=v��qy<-q�J�9��NM?�W�?���Ӻo��v����=�"i�YN?�l8?���<JҾ���>��]?Ղ?��Y?���>8�������m������wЭ<�?>0��>��>|��XU>��ѾI�I���>�~�>T�ڼo0Ҿ�͉�+�Fĝ>�'?���>jʮ=�� ?x�#?İj>eA�>�aE�~>��� F����>���>X9?Y�~?��?����b[3�I���㡿��[��N>L�x?�X?Rƕ>⎏�ᆝ���E�.�I�iv��"��?L�g?~��y ?v<�?֋??��A?Ef>[���׾䌭���>��!?��M�A�PM&��	��~?�P?���>�-����ս�%ּB���|��� ?(\?�A&?����*a�t�¾�)�<ͤ"�� V����;��D��>��>�������=�>�۰=�Nm�G6���f<{g�=��>�	�=�*7��q��'=,?�hH��ڃ��֘=��r�dsD��>?CL>.����^?��=�h�{�����s��4�T���?h��?<e�?����٢h��)=?��?�
?�2�>�F����޾̠�̖w��x��m���>���>�n��-����n����E��/Jƽd�p�A�$?��>ݸ>�$?^��>t=���"�R��t��#t��'�*�W�Z�V���E��ҿ���~1���վZ����׹>�6��yy>�9�>�[�>u�&>�^�>Y.>��>3i	> s�>
�>�q�>���=������Ѽ�0b��KR?�����'�C��H���3B?Sqd?2�>�i�؉��?����?���?+s�?s=v>g~h�3,+��n? >�>���q
?�U:=i�&;�<�V�����4��M�ѩ�>�B׽? :��M��mf�fj
?K/?���Y�̾L9׽�˕�M�=�	�?��.?��M7�$�\��If��vQ���*��K��m4���U5��|�a���!��j��o/*�e�<�B?�?����(��P x��rR���l�q�>>L3�>lht>�g�>�?>{�־҂�QP_��+*�l(����>�|}?�E$>ga?�U?�_?#�??��=�t�>��[�p?.\�M)T>j��>�7?�[?�a?Β?�E?=��>�����<"���Ҿ:�A?�5	?��?`	?�}�>8��!��<�|�=����x���V����0�����@N�;@H�<9�ѽK�=Z?�����8�����k>��7?*��>&��>&
���!���n�<_�>!�
?]L�>�����sr�V\�:Y�>���?�+�ù=��)>���=�Ņ���غJX�=�¼7�=t>��-m;���<�`�=�=�Us��o�$��:�'�;쭯<�t�>6�?���>�C�>�@��.� �c���e�=�Y>4S>w>�Eپ�}���$��v�g��]y>�w�?�z�?ϻf=��=���=}���U�����H������<�?=J#?(XT?`��?y�=?^j#?ε>+�iM���^�������?�+?(��>$�P�ʾ�����3��}?�l?5a�'��')��¾!oս�8> -/��~��ﯿ�C�懍�(��iј���?�Н?�8B���6�c��Ϙ�<��<lC?|��>*�>���>��)���g�3%��#;>��>��Q?�#�>}�O?�<{?��[?gT>F�8�{1���ә�@I3���!>
@?ʱ�?��?'y? t�>��>�)��2T��	����*ႾXW=�Z>ڑ�>�(�>��>���=+Ƚ[Z��$�>�@b�=��b>��>���>��>��w>�F�<�<S?V��>�\ʾx06�+���'5F��,�P@p?��?��q?��/<x�� 7�k,V��f�>Kߟ?�
�?�S?�g���I<��=Kߜ�q����:�>d��>�э>:N�=��ʽxR�=� ?���>��� 6�M�0��eֽj,.?�{?�\�=c|ĿJ�m��7x��q���U"������h��S��q�U��(�=#p��{�	�W۪��kZ�����̘��Pط��'���~�@.�>"�={��=���=nV�<���Pq�<�P/=�ٚ< %=F�U�3��<]�O����":��H�*���V<d2=:LP�ȱ˾�}?�I?o�)?��C?-�y>��>h�M�H�>x슽k?-LM>��h�Q�� �D��b��c�� Cھ�*վ�f��Z��˜	>P�U�4�>�2>�3�=��<��=�h�=�4�=ߌ���o%=p��=S3�= �=>P�=,�>�>��{?%������aq\�=V�Wo-?b��>�>?v�fH?G�=�Ʌ��]¿ǲ���?�`@u�?�'?,y,���L>�bX���x= 0=x�þ0F=>M�W>�Q�]��>2�K>b�N��֚���D�BA�?�@��^?�%����Q@>��->�u	>H�T��73�m�s�CCu��b^�<:%?�7�,�Ͼ�~>T��=�X߾��ľח:=��,>��4=��{�Y�1��=`�S�]8=mf�=?�>��.>���=�սYk�=ؠM=7b >lrP>��~�+ke�w���=7��=v�U>�J!>G��>P�?p`0?XXd?7�>Xn�FϾ�>��pJ�>��=�H�>��=uvB>���>��7?6�D?b�K?���>��=\�>�>�,�մm��k�(ɧ���<o��?�͆?Dи>��Q<s�A�ɠ��f>��0ŽUv?�R1?l?��>�3�7����Z�$�h�4��J<N>���K�0��<KQ�`9���Q>sG�>��>2��>�|�>ӥ>�ƃ>�q�>x�=�1����">�3н�b���Z>D�=�3
<O�p><Yu���H��(<��<`�;�.һ���;�B�=ҴC�?Σ=���>r��=�`�> �	>K#���?>���!y�+�i����~�L��t�AT���<��17��9>yă=��i�x����?��W>V�5>�?[.l?jb�=M6�\���Β���T=����eV>��c����<8D�!Nx�T5�X����>��>��>��l>Y,��!?���w=.�a5�X�>Ez�����)�Q7q�?>������pi��غK�D?�D�����=�~?ƳI?dߏ?|�>E��yؾW:0>N���="�'q�Z����?'?'��>����D��H̾L��"۷>�II�c�O�;��0�V*��̷�H��>����R�о�#3��f��&���Q�B��Pr���>ڴO?m�?H6b�~W���QO�/���/���p?�zg?��>{J?B?K��{��s���{�=�n?:��??<�?�>��=$�ֽ�x�>5R
?�d�?rܒ?հr?�?��
�>�"/<"�0>1����C�=9>J�=��=�b?��
?m4?�b��Ț	��9���e󾥗Y��1)=��=�>�>��>��i>���=Kp�=OÒ=�bZ>ڛ>Vю>_c>���>sɆ>_졾;W��G-?pR�>�ݱ>4g3?冸>K�"�Fm��
S7>^�'> �<��������I��[4�=q��=�	�?#����?�ԿaMZ?�+�>3��^?�SJ�d�ܼ8��>r��={ԃ��� ?�\>�	�>pʚ>�&r><�>_�r>�.>�	ɾ��B>`���;�C�[��i�QӾ��u>+r@�r$���������uq������]�&�u�FG����=�]Ֆ=ʚ�?�6W�	�n�<�&����b�%?��>v40?f����r�;�g>3�>�º>��ܾKq���^��Iwھ�?}G@G:c>W�>��W?N�?*�1�Q3��uZ���u�q(A��e�V�`�፿$�����
�Y��*�_?8�x?�wA?�O�<7z>£�?��%��ԏ�|*�>)/��(;��?<=	*�><)����`�įӾo�þ,5�+EF>'�o?�$�?�Y?dOV����g>+�7?�??N\h?�9?:�C?]�1�Cm3?k�Z>M�>@�?2mG?�h4?��?�p>� ^>�|�=��~=�g,�A����ͽ�r+�Q71<�-=��'Ʋ<�� �
1�<썐=s���c�$��kĽ1����O� �ɽ�}�;T�>�զ>U�]?�&�>^	�>��7?Ii�zq8�86���</?zt>= �����������w�E>�j?5��?sqZ?��c>�qB�*gB�(^>�{�>�B'>�[>r]�>���&F��0�=� >�>)��=NO�`���^�	�e����a�<��>�	�>�OE>�<�����=s��/�U���>A`��R������h���:��3;)|�>�X?2�(?@ZP>�����ꀿ[{G?%7*?*�F?ۑ?�"�=C���L�\ǁ�:����>��p=��޾B���U��Y	t�C��Ѡ>���������O^>���#�̻l�tT��㾄��=+���1{<e/��}ž�B����=�>A����'$�����(���zK?�C=�M��qY	��*Ǿ!U>��>"K�>E+��k���3�.�����\=�=�>�C>}b¼꾔sG�w��{q><�G?֣_?n�?���tk��<!�x?�\Ǿ����L>�>�ؙ>uq�>�(弆�s>�S�TQ&��Ȍ�Vt'����>�o�>����E�E���]�޾AO9��č>�tM?���l�>�֒?$��>:�K?w�1?�3?O�F>+���͹���Y&?,o�?Ԋ�=:Yӽ��U�?J9�_$F����>�)?�'B��j�>��?��?��&?vtQ?}f?��
>�y@��d�>lT�>�-X�[_����^>��J?-*�>wY?F߃?U^@>5��n���v�����=�>�p3?�#?Ƚ?<{�>Ή�>'���~�=��>�c?�.�?c�o?s��=�?�52>���>�R�=���>��>�?�XO?��s?R�J?\��>�<xZ������us�\O����;�H<��y=�L��s�,\�*N�<��;d��6x���򼏫E�g���O�;td�>H�}>�����5>����b��	)E>��#�������u�"�_C�=<�>)?w��>`�[=⩼>Ŏ�>����"'?$u	?YH?X�;�c�(�Ѿ�k����>��??u��='n�����
�o��BU=�,m?1`?��X�w�[c?D�[?P���)8��	ɾ�y{��쾀�T?��?��<�k�>��?q?�\�>�9T���i��Ĝ��e��8n�'�=)��>�P���f��/�>l�6?���>�/c>�g�=�|þŲw��Þ�Y�?��?ܭ?^L�?�->�f��G߿i9�f|���lk?d�>�k��3@?�G;�Ծi�P�����OپC[��DȾeS���ȑ�<c!��jx�!�&*7�X ?��k?+�c?�E??)����n��>:���~�z�l�%��O����5�*eA�T�5����X"�4���ȾuR�<4uw��F��5�?V�)?2�@��w?!������%���=>sޠ�Ĩ��Z=�ݣ��Hu=8�m=�Z�I�4��.���j?��>/��>�u/?�([��^=��i)�8;�<;����>pj�>�n�>;�>~����tE�����۾�|��@򽅫W>ei`?w�K?>�w?B�M�
-�s5f�:���R�W���I�k�~>l�a�P�>G�?���]���C�>�B�vdx�k྾�/�����=n�H?S��>���=D�?J�4?]����#J��y��Ɣ=��N>�	�?E��>b�k>�8���B�:d�>��h?��?��^>e꺾���m��(�C���>3��>���>G��=����v@�����(����=��a�=8�?r�g���a�WJ>�s?�5���ͽ�y?G�>
�"�xq��"N<m�=:�"?)�=Ꝛ>Cþj��ͨ���Ɛ��"L?�.�>gH��7;����=t?%j�>�c�>a��?x?L���w�8>�H9?0�w?,GV?�Z?~2�>}kH���Y�T��$����?>��>�4>�ڈ��F�ڤ��&�S5Q>0'�=�\�T��������֨>@\R>_�\>�{߿HK�t��/j1��Ѿ��h���Z���<Xf��P�"���`]��lD��~�8����E��T�&_j�%v��*�?�"�?�����&�������������E��>(j4���ݽ����׽��ԾOn�xn������Q�� S�߶i��&?�0����ǿğ����3�?�8?~y?;
�F<$���3�P�>�8�<�!ļ��������οSǘ���^?���>��� ��=c�>�O�>�_>��f>����柾:�=N?��,?���>���Nɿ[ź�^��<���?=@փA?.�(�`��8�U=E��>]�	?4�?>o*1�H:��װ�FX�>�;�?���?#�M=-�W�k�	��{e?x�<�F��g߻�P�=�\�=7"=�����J>�A�>�K�(A�>hܽf�4>ׅ>�-#�#���u^�2��<��]>fս�m��:̄?E|\���e���/��u��:�>�T?���>��=�t,?�8H�,�Ͽ7/]��`?��?w��?��)??�����>�#ݾ��M?g6?P�>��%��u��N�=�����э�$�V��U�=p��>|>�X,����7vP��m��J�=���ſc"�w�-��`T=.I���n��c�^��V���3��Z�M�����S�=[B�=��a>�`�>�N>��L>�a?
r?��>s��=�Z���6��D̾� ==�h�5��N���! �̼��b@���ZѾE1���l
�uhҾ"F�;�=[�Z�����tO�����l5���.?��Y>������l�Nv�=c�۾R<��2�|<��<���ྜྷ����s���?��D?hS��$!�x)�^$
��"��/R?ؙ���_�%�j�)w�=��y�"L�<�>L�s<����4��a��l=?H�,?@߾����E?>�)����H<�qP?���>��)>�?�E?��<���=.��>�,<>ϯ�>`U�>Q�I=�پ�s�� �5?��t?��Y���<�>��������f��@!>e��&q���p@>dO�=O���N�=������= EW?���>�*�(1�C��e���?;=X�x?=�?�ߠ>�mk?�C?v�<����S� �
�Y�x=�W?��h?8:>�4���Ͼ�{��z�5?[�e?3WM>�g��Q�Y�.�R��-?�|n?�7?�Ο���}�V���&��W6?��}?�v��������["�.��>�>C�?Q�N�,/�>��l??V5�����(Ŀl$"�_�?��@}��?rߣ;�䎽}��=���>
��>�;���n�����&��H�<*��>|������8Q��L��t/F?��?�?�:��Ȉ����=Kɣ�B�? �?��eڎ=t��a@i���6BϽF��=uT^�E��������:��x־����̾�۽ip>�8@�r��R�>)Q'�9俸�����m�+O���Ǿ�?�ŉ>CU��h���Z�~���z�մL��uR�?*��2�>xf>�������Μ~�G�L��� ��?�=>hK�>���Z罓|��tC.>��>�C�>N8�=dr��yᾌ,�?)��A�ο2������b\?���?�[?D�)?X!�>��������_:�>qЂ?�n?��?��=ϮȽ��N��j?�a���U`�d�4�oFE�OU>_"3?fB�>G�-��|=�>��>�f>$/��Ŀ5ٶ����s��?��?2o����>w��?�r+?�h��7���Z��8�*�A%-�d<A?N2>݌����!��/=��В�`�
?y0?�x��.�`�_?)�a�L�p���-���ƽ�ۡ>��0��e\�M������Xe�	���@y����?M^�?i�?ڵ�� #�_6%?�>e����8ǾJ�<���>�(�>
*N>�H_���u>����:�i	>���?�~�?Oj?���������U>�}?���>F�?J2�=P�>�d�=摱��g�n%>���=��5��j?q�M?���>�=Έ5��z.�|E�({Q�S���D�_�>��b?M?�Zb>B���$&��S"���̽�1�n��YC���+��'ڽ"�3>q?>�'>�#E��Ѿ`E?�0f�tӿ��q��3%>Z�?U?6>R@�><����dw���q���Z?��>.��f���P��SP����?�f @���>�6�ml>�
�=��?�%>$˃��EN=�d����>7�,?�eJ��v�!�F��N�>D�?�&@�ȡ?7Y��[?��(�z<���gf������S8��_�=tbB?��ݾ.}�>?H�>!�j�4���j�d�F�>�Ա?���?�y
?	WL?��K���"�e�����>Ii?��>��>cn�LQ�=h6$?N�n��<��i�R?U	@fC@�kb?�筿ۿῐ>�����߀Ҿm?�=ڥh=u�'>6����=s�<�c���=�N>��>�i\>�t>GD>}�6>6vI>[����r��a��L�����7���'
���8�ɿ����[�=��a���jr��1�RO���Z�dQ�n���H�=�U?�R?zp?�� ?�;y�~
 >����_"=�A#�`Q�=j#�>Lk2?t�L?;�*?f�=���U�d�*W���=��������>9KI>u�>I�>;!�>KLy8��I>�?>�{�>.&>@�'=~F���
=��N>�G�>���>8c�>�Q.>3�>����� ���h�5����Pͽ�{�?挾K��ᕿW�|�"5��(��=��-?��>�M����˿
�����G?��������5½5��=�/?��O?"z>^���W�W��J+>'���Lh��>�㽡�e�0"���6>�<?��1>LK>��A�g,$��#`��i���P?>�^7?�[y�G+��k.n�С(����|�6>}L�>�\׻$��玿<�����'���<W�)?�[-?�����`� l<����5�e>lG>R>k	?<�z>��h;DU���W�{[�<���=�I�>I[?p->҆�=� �>���8�Q�h��>�}C>�;*>\@?&�%?���*y��v����+��Hw>~�>;�>6�>mDL���=���>�?d>�/�8ֆ�/��=�D��hW>�-~�<=`�R-~�j�x=W��DB�=�;�=����r =��s*=�~?���'䈿��Ie���lD?Z+?� �=��F<��"�E ���H��G�?q�@m�?��	�ޢV�7�?�@�?��=��=�|�>�֫>�ξ�L��?�Ž1Ǣ���	�)#�fS�?��?��/�Wʋ�3l��6>�^%?��Ӿ[��>�DY�'�����a���n���=:'�>�7?gN��㨽)� G�>���>����T��PLĿ1n��g`�>�g�?�m�?�������(U6�W�#?H��?�n7?޵=��Ӿ��2=��>��??�}S?Z;;>�)�B��!?�S�?ls�?���=8`�?B�?��(>��#���ֶѿG?������&=Խ�I=:�2�q�߾�0�zn��_����Y��߆��?�v9=-��>N	l�_� ��#A=��=�禾2潂_�>�
?״�<��>���>���>?kQ>ߥ�ġ2��V=�l����Q?�B�?z�r��Չ<���==a�U�
?��8?��k=�����v�>(Ma?C�?�Z?�0�>>���+��*B��%���.a=��7>P��>RY�>l;J��8>� þ��o�Iuq>wN�>�T#;�sj�����q҃>5�?2��>6�=K ?��#?�k>s�>�OE��Y���(F����>}�>0b?h�}?F�?�
��� 3�"��	���?�[�/F>K"x?�?�֓>�ҏ�m���Cb�9yF�����M�?�yh?�~ݽ�?�U�?��??lD?��c>o��C+׾�Y��N>%�$?����"A���%�ѹ��?+9
?��>�>�ę��h'�t���뾵q?�P^?)?|m�>�a�K�Ⱦ���<��_�꒼\�-�GD��R->��>�m��3z�=!U&>!�=vo��2���]<K��=�ۖ>/'�=�",�9{����)?�׽Y&��6/��}�v���=�p�<>��	>9 Ѿ�7?2���� ��s������89I��Ȕ?sQ�?�a�?��%���o���O?���?X??x�?
��?.�<��VA���&���r��>y>��?�e���9�ڲ�����6���s�̽0)U��Q?|�>8��>6?	��>w�>�˾)�E�E���:���A�n���KHG��8��1��Ƌ���E����-���\Z��>P�=Kr�>��?���>�\�>�`�>���=�g�>8>E�>%�>&�P>fH1>]�>�x�<ߏ��&LR?`���,�'�Ƿ�Ӳ��83B?�qd?�1�>i�ɉ�������?���?]s�?x>v>b~h��,+�9n?�=�>C��=q
?S:=�5�3>�<�U��ݼ�04��O�몎>�B׽� :�|M�*nf�Rj
?p/?v
����̾U:׽�����4�=���?�/B?:C+�rB��S`�J?���W�M���C �#��w�5�5�g�����(���LM���I�_�=�V?���?�~����b����S���m�ǭ8>���>�^>��>ʭ�=&ξ�.��Zd����FBi��?�-�?�E>Ҽf?�g4?��O?w�J?��>���>�b�����>
f�=���>1g�>�D?�-c?�C?�?��F?���>�t����~u����J?��>�E?��?�&?��f>�I�Iq��L�g
x�LB�=eL<0�3:�v%=�=ġA>0Y?J��K�8�	����k>�7?�~�>��>R��o,�� �<-�>r�
?rE�>�  �w}r��b�zW�>���?��b�=��)>���=t����Һ�\�=	���"�=:���f;��\<��=���=Rt���}�-��:I�;Tq�<�t�>E�?��>jC�>�@���� �����d�=?Y>KS>�>%Fپ�}���$����g��\y>�w�?�z�?��f=��=���=}���U�����������<ݣ?"J#?*XT?F��?Z�=?Qj#?�>�*�cM���^�������?C!,?B��>�����ʾ���3���?�[?;<a����:)�	�¾��Խ��>[/��.~�m���D�������z~����?���?xA�"�6��w�����M[����C?�!�>�W�>h�>��)�J�g�%�c2;>���>{R?�#�>��O?�<{?��[?sgT>L�8��1���ә��I3�>�!>@?ⱁ?��??y?*t�>��>a�)���$T�������Ⴞ*
W=,	Z>k��>�(�>)�>��= Ƚ[����>��`�=��b>Y��>���>��>ޅw>)M�<�YU?~_�>�оG������J�b.�d>v?�ݕ?�9F?�|�<=��������r�>5ڪ?N�?��?it����=��4=h�¾�Ď�T8�>���>�z�=�H�=�Լ>�>���>!��>I�>����!�<��d½$�?��N?< �=��ĿAp��w�b�����;L��5d����e$S�+o�=�5�����}W���Y�2A���������d1�����iO�>i�=N�=�6�=j��<y5��c�<@AC=%��<�=��O�H2<X�(�[���L����!⻸<niQ=��:/�˾yu}?�*H?�++?�gD?{�}>)j>�A�ۊ�>�h��	�?^�P>j�R�0ս�`�=��F���o��ɧؾHrؾ��c�c柾��>��4���>�5>j��=k�<Խ�=N�=z�=�v��)=]y�=�ʽ=�=��=�>��>�	y?8󄿅����Z��7t�=�>?��u>h�>�վ7Q'?E҃>�đ�N�ǿ���L�w?�=�?��?(? �����o>'gA�i�c�L-�=�U�/9 =�y�=i���8o�>	'<>BJ��ۧ�U=�'�?��?��1?5n|�~ο-^�=\b$>]��=��U�b!�a,�������S��o ?��'��a��s>l6�=i	�R����9c=�+>�4<�&�8u_��l�=%u��?.=�*�=�G}>e>fK�=���c8�=�|�<�n">ʤ->�_�</��������<X�x=�r>5�c>Ò�>f�?�a0?;Xd?6�>in��Ͼ?���I�>�=	F�>>�=lsB>T��>n�7?��D?��K?х�>���=I	�>�>S�,� �m��l�5̧���<���?�Ά?Ҹ>"�Q<l�A�����g>�50Ž�v?SS1?�k?��>�r��߿�"�A�;���+���V�K8=�C���4K�^��n�R�������>ޭ>��>�O�>q�o>](>��G>mN�>qN.>k�(�-;�;W�H�&��lر��>P�r��h;�ذ�mǦ<F^�`o{�h޻�u�<}a��a�<n���E��=���>�?�=䴨>*�>BՈ�h�=�d���q���/�}#���xN���`�Ө��tE*�ߥ$�*�o>�(>�7��w����?_>[TG>>��?܇??L>�\� �t�����<����t>� �<�M����J����xX��d׾�S�> ��>x��>hSs>�n,�j�>�;tx=σ޾��6���>Z����=K�Fd�c�o��⤿�w��Qi�?_�ĨD?�~���7�=�|??7K?-L�?��>(�~���ξB�&>lZ��a=�L� �j�gy���?�'?9��>�0�B�F�5<̾V���ѷ>�1I�L�O�m����0�����Ʒ���>P�'�о!3�Zg�������B�scr�l�>a�O?v�?�Pb��R���UO�U��� ���h?�og?��>0U?6?���h�q��+r�=��n?y��?�>�?�%>^`�=J���0E�>�)	?���?��?��s?ֺ?��|�>��;�� >r������=�>+ǜ=_\�=�v?��
?��
?w����	�-����C^�qq�<�ϡ=ă�>�t�>�r>���=�g=R`�=x\>՞>��>�d>b �>�K�>���V���Bt?��>ʰ>�so?fi>N�<*瓽���.=>;���\�X�ůQ�iW��A�=��
>�r��2s!����>(�Ͽȕ�?/̀>��7�9!
?�_��vt>�"�>g�E>�|��g?P �=��>�?�ۜ>h�>��V>�w>Rư�z�=��+�{�ݾ&�]�4�F�#����>��ܽWþb���5����Tp��x��0����b����<#�Lв<�t�?�8�2(w����ӂ�X� ?usX>r)?[���o5�<@݆>^z�>���>�o�%���Z����n���?�[�?m9c>�>��W?H�?��1�*3�qxZ��u��'A��e���`�8፿����~�
� ���_?�x?�wA?|��<�8z>���?��%��֏�*�>!/��';�r1<=�*�>\"����`���Ӿ�þ3�IF>E�o?�$�?c\?�NV�o���mO�>�Q?��?��?�c�>�ڃ?b����?%�>g��=��?rL?��b?�8?34�>�'>�ޔ<��<Kӥ�4׷��^��ǽ���r&+���=�u�=o b�;�>�K=�e��|�<L�㽊��h'������i]���;�>�]?�R�>Ė�>��7?����r8�IҮ�*/?��9='������o�������>1�j?k��?�cZ?med>{�A��C��&>jM�>�t&>7!\>Qb�>�|ｋ�E�-�=�>>_`>���=��M��́�	�	�����\�<n">4�>��{>䎽��&>و���z��jd>Q�ݐ���R���G��1� v��T�>
�K??4"�=�1� ��Gf�eO)?37<?uM?��?�_�=<Sܾ��9���J�����`�>�ͯ<���񴢿,)����:��43:�s>��������/z>��
�w�����p�dL����WQ�=�d���=����ƾ�������="�>L�������8��>D���G?�"%=�畾��W��D����8>Cp�>8�>�{��������<�y^����=�0�>��">_�z�����=��	�s�>��A?7�[?>5�?�_[�W�j�-<����q���R�<���>9��>��?b4>p�:��u���b`�+E���>���>)? �I�L�`�~��Q%�(��>p$!?`>s��>��>?8�?Y�`?v?L=�>'>R>�(T� 쓾=#?	�?�=���ʾ�X�4!O�V?VIj?�N�;��/�>�E??��?Q�>���>�g׾�)�o@�>�s�>�'Q�%㷿wf�=h�1?m�>��e?�BG?� �>�(��V���S��l�=�=>k��>�� ?J�"?�@?b]�>�]���.�=���>+c?靂?=o?Q��=�L?��+>�d�>iC�=/�>`b�>�%?��L?��s?�,J?��>���<�ݭ����}-r�8SR�P;�l<z�k=�E���k����҂�<���;�F��ݣX��ͼ��C�Я���,;z��>��v>�����/>�Kľ$͈�
j?>D�ü�g��s���>;�e%�=�s�>�a?ao�>�V$��:�=S�>g��>���r�'?��?��?��;�b��پ�#K���>�FA?�n�=WAl�P��)v��q_=C�m?k^?�OX��|���b?� ^?*k��=���þ �b�w����O?��
?��G��׳>��~?I�q?���>��e�j3n�&���;b���j���=�a�>�L�^�d�SC�>#�7?�A�>T�b>e��=<@۾n�w�Ln��?���?|��?��?� *>�n�>0����m����\?��>�Y��QX"?�]���Ͼj������1��
���)���������%����FaӽR�=q ?ar?�p?eh_?u�� #c�9]�T ��9�V�7�S��:G�L�D�B�1�l����/��V���M�J=XtV�ޑ/��6�??�"?�у����>�t����ɾ����h/�=����J��Օ<�L�<�p%�Y�H>�ҽw8���ѾrL?���>@J>�#?��9��g9�����B�~��M�/>f y>&�5>���>� ˺�T�gg`�5����$�k�=^~>^�Y?O�W?� c?�IL�N//��������E9������KVX>F�=��y>&E/�џ���O;;�U$k��9*��a��(S�_�r>�3>?�IR>�x�>' �?(��>�t�����rE���Z=��>��g?T� ?!��>V��.����>��l?�|�>��>pn���g!��?|���ý��>4��>�,�>K�q>KJ/�G[�=���/����8��=��f?�ㄾ��b�/�>b�R?7B�:�rN<��>ݪ��Z�!��g��$�*�>�d?5^�=�?;>?�ľ���{��ӊ�8�2?��?�Y����$�3�=�N?���>��>Ww?QN�>��u1��?{g]?s�?V� ?�?��=C�R��n�yNڽH,��;�K>�3>���<, m>D����9��xSz�m!>��=�?����Fi=�������F�G=3��=�bο��8��7�����x��l��vᇾTL
�d�O���	���6��%��x�޾c��sg>���@_ھ|M��`=���?(r@�컛.y�����ʠ�#�F��=�>v�=Y\������[�=�e�#	��'������̾>O��5��t+'?�ē�`Tǿh렿�ؾ.%"?�"?��w?�
�Wv���5��� >�>�<@��(G�Y3��͔οp�����\?�I�>s���"����>N�>�P>�lk>r����uQ<c[?D**?vi ?��c��Dɿ���<���?N@��3?}Q��������>q&?�F"?���>ţ4�V�%��Ҿ�*�>��?p��?Mx�p\\�h���3H?��v��{+���8���9v����yP=	μ#�>Y�>�Y�!��z8 ����<��A>/�<c�<�"?��?��i�>S�e��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=s6�����{���&V�~��=[��>b�>,������O��I��V��=dK���%�� Ri��z#��pd>}_=�t>?�ὖ��������[=�Q��Nu�}����>n7�=�����9�]��>4 1?�I7? �>7��<g(=q��E����8�|��	>ʄA>s���ֿ��ƾB� �.u��b�h��
Zྭ(�bȍ>^�;�_'���@F�����`[� �M?}�>J��B�o�[>x��2���YN$=�L��w�K��>]k����?(�a?�7>��NM���C��?��fVd���?Z��;[h������Ç>��>�=���=���>1����F־��%��B?4�/?�����\ľ��:�x��1�<��C?Z�>B>�V>a��>2zl���߽&q> �E>�>WD�>d�\�ќ��(k0�ֆ)?n�_?�pݽζd����>"毾-Đ�Ǫڼ��[>��ټK��㽕aw=��;��E��(1�_�c=.;U?���>��(��q�Υ��Yo���|)=mR{?�	?��>��d?��C?sc<Al��\P��
�ළ=�uT?�d?�j>����;�о�O��T5?�Rg?vV>�j��t�Jw$��f�P
?�Sg??�ѝ��Lz�����>.�ؖ3?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?p�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������'��=ix��/ �?�L�?�ح��&H<����i��W��	|�<���=�<l�3���羓�6�;c��$��FZ��1�s�>- @#� �}��>kN4� ��QEͿ�Y���о�.i�$f?Lo�>$꽽����c�k�v��D��_D�񀂾{4�>��\>N�ֽ5)��´��,�P�����	?y�o=1�p>;�~�1i��b�������ǔ>)�>�>}����պ��?�_��%N����� ����k?��?�w?�?I>�\�{����I?��g?ΥL?�>۽ѕT�6Ɇ��j?�_��~U`�ˎ4�HE�]U>(#3?�B�>��-���|=q>D��>f>e#/�K�Ŀ�ٶ�i���'��?���?�o����>P��?�s+?�i�8���[��\�*���*�^<A?�2>w�����!��/=��Ғ���
?l~0?y�'.��N_?�`��1o��t-�O-Ƚ���>��3�B�^�������e������x�ݭ?�?bM�?9���!��%?���>�����nȾT��<�-�>>`�>6�L>�l��u>v ���;��]
>���?��?��?f���u��Sc>��~?
��>���?�
�=�>���=ձ�=���|�'>��=�1&��z?,M?���>`x�=:��'.�eF��/Q��
�N�C�ǡ�>�]d?�N?��_>�v����6�H�!�Caͽ��5�xR���I�tj����m8>SB>�>�J���Ҿ��?�p��ؿ�i��Yp'�I54?���>��?��e�t�����;_?�y�>%7�,���%���C�?��?�G�?��?��׾�O̼k>��>�I�>��Խ ��5���{�7>1�B?#��D����o���>���?�@�ծ?i��	?���P��Va~����7�a��=��7?�0� �z>���>��=�nv�޻��X�s����>�B�?�{�?��>!�l?��o�O�B���1=8M�>Μk?�s?Ro���e�B>��?#������L��f?�
@u@a�^?*��ֿbQ��#�۾XgϾ/����+����=�	:�%r>\��=�At=��>��=�0�=�Zp��=�ݡ��v3>z��>����1!��𩿸���ț-������%�x᱾_!��(���������V�Ⱦ�l���r������8~��ɹ�س�=.-�=��)?���?`�[?m]>JL��i���/>��&��=�7½��e>�{�=�'?�cB?��?��>mDZ��aV�
��K=þN�ľ@��>��D>���>�O�>!9�>Hqȼ�TY>��,=&ݜ>�e=��&<��<F䀽-X�>�v�>���>0 ?,I>EoG>�K��ѳ��m�u�����Y[�?�p���WA�:���[z�gxʾ��w=��+?l�=tb����ȿ'��h�E?'���KZ
�~S�ߩ>D$A?�M?�">Pžp@!=Kz>Q�����*d.>���`�a�;$-� �L>�I
?�+n>�A~>�1�6f<���Q�F���S�g>n:?���� J���u���A���R�W>���>�y�Q]�ۑ���_���Nf�rpT=Ɨ;?��?�p�����Jz~�d���2DG>W[>��=ͻ�=�YS>@�^��Gѽ��D���=�=6�N>]�?�܋>��4>J��>���B�'���>%�=>'o=q?݄?v��J`(�DC�S6����!?h��>}H<�Ԓ>�jj�7�~<+�?|�>�zd>I�λ����4��f��=g��kv�����=y�(=E�d�_>�Z�>��0���I��%>s<~?�b��U݈����`�����D?x�?O=�=�{<n5"�̦�RN��p��?A�@��?H
�-V���?8ԍ?V�����=�9�>�V�>l�;�pO��?��ƽ�	��4"
�M�&�0�?�9�?fI��j��y-k��F>X�%?#ӾXh�>�x�{Z�����r�u�ȹ#=���>�8H? V���O�>��v
?�?r^򾾩����ȿ%|v����>�?���?<�m�aA���@�I��>��??gY?�oi>�g۾`Z����>��@?�R?��>�9�~�'���?߶?���?�hI>m��?��s?��>p�v��/�-�������z=���;�	�>\�>�J��_F�����-K�� �j����Uc>�v$=<�>�&��񻾘z�=�׊�18���e����>=q>�YI>���>�?��>��>!�=4��Y������[�K?ⲏ?���.0n�=-�<�z�=��^��'?�C4?GG[� �Ͼè>��\?@��?{�Z?D]�>;��b9��)㿿=w��ã�<��K>|/�>�3�>�&��{�K>��Ծ�BD��`�>9ٗ>Y`��DھD?��ރ���E�>�[!?���>î=`� ?�#?3{j>���>xgE��<����E����>���>D?��~?d�?!繾�S3�����$᡿"�[�y9N>�x?�T?���>U���􂝿��C�Q�G�;�����?�]g?���M�?�+�?3o??�A?Qf>����ؾ7}���ހ>&'?�ž�5S����i��=*uZ?l�F?�1>.s���Z�=м�>��a�1�B�>�GM?.P�>.�w�u�#������<�Dg<@s���K���
��:>9>l>=5���7�>(1�>��=%�Z����"�=%q�=��:�a��� �F��==,?��G�Eۃ���=��r�:xD���>2KL>�����^?�l=���{�����x��;	U�� �?���?0k�?���h�d$=?#�?�	?�"�>�J���}޾���Qw�;~x�;w�1�>+��>Ưl�h����������F����Ž��`��>M��>�n?$�?�W>�U�>���|I(�
�� q���mW������6�.�����%��L0��%l�����GŁ�K�>
*�����>[_?Q�g>��p>Y��>H��7�>��L>e�>8�>�o8>��%>��>���%��9Q?��¾6�'�C �����:vC?f=e?{i�>
�[�Vㄿơ��4?đ?�X�?Wp>�h�1�)�	j?!V�>~��1?#.!=!T��<u����������~ �u9�>2�ٽ�8���J��A_�.�	?�6?lZP��"Ⱦ8�˽E���e�n=%M�?=�(?��)�U�Q���o���W� S� ��0(h��m��m�$� �p��ꏿ�^���$���(�^^*=�*?-�?f�����H&��)k��?��`f>��>�>�־>�{I>��	���1�/^�M'����TR�>Y{?�G�>
�D?��@?�]?&�L?zZ�>��>�|վ޾�>񋘼T�P>���>�HE?��?� ?B��>�M?��>�Ԁ������<�?�H7??O_�>DJ ?.d���Ͻ��#=%=܏��,�̽gH=��2�/�����u����<��9��?3(R��Y2����r��>��=?x�?]=]>0i����Y�m߭�s/�>gu ?�)?�T������G�߾�?�[?wo���=JD*>+��=���\�齷T�����1I =:콽��ؽ)l=4�[>_5>n��;�I^=U��=vt�=��y<'k�>�?���>�E�>WN��=� �������=
�Y>�Q>{Y>Q�ؾ�V��.��%�g�Cjy>4w�?;a�?B�e=���=�c�=^���!z��+��r���a�<[�?+#?qT?*t�?М=?B#?��>���,��_���G����?��,?�s�>�X����l��'�7����>��?��W��P���2�ĝ��m�I�Q�0>�/�/�r�ڭ��-.�َ��������n'�?q-�?��'���%�~���鷙�����)?���>��h>`J?R)�[U��D��>��>3�;?�Ժ>�+M?�?��S?�D>,�.��5��j����9׼o*(>�T9?Q�n?�?�	z?~��>>�>�������,�a8��8ؽ�G���hJ=�d>���>� �>��>���=�sʽ$-����<�q��=,Q>)��>��>�j�>H�|>�#=AF?�H�>�Ǻ���"�8cǾG\������Z��?��?j�/?Y����zJ��:׾�|�>O�?��?c�!?zf���>̱9��|��4������>u��>��>y��=]���^n>���>%X�>w�]�S���0�
�E���>Y�C?=2?˿�S���u��F㦾|�<��j�b�-����a��J�=|8p�v4��[4��u¾����'(彀�����ɾ�9E�^)�>�7�=��=��>��r=:Ä���<�d =��:=�-�]����ϼ[(�9@�=C}R>��9�7,c���=>�^�<�ʾA�|?��I?e�+?�PC?��y>�x>d25��>j���?�ET>Z�J�5w��=�p%���ᒾ �׾{ؾq�c�]���N>r�E�h>ڲ2>�P�=��<\o�=r�k=.B�=�.����=�n�=dc�=iI�=�!�=�(>�|>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=J����=2>r��=x�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>
�_>�<>!KH��~I�h���J��Z����9?�*��~��47>�>C�����Q��<�>�	=_GŽ�a�3P�=r�ȽЙ�=��=�S�>[ZU>G;3=R�ɽ�S#=���=�a�=��n>(�Z��些w����T=㻚=@9v>bB�=�[�>^�?��:?��e?��>]lz��5��0aq>FA�=lCb>�p;�}۔>Z��>]I?��7?�O?MŘ>ڍn=�E�>(*�>�"6��n� ��!���������c?f?�?,P�>t��M����J���I��%I����>p;�>���>%v�>a���Oܿ��/�)�!�F��޺��]�X=�+m���)�2 }�����=7��%��=3�>EC�>V�y>�>S�>Z�> ǿ>�" >�!=��=SUS=Z:��5=e��=S�<����r��Γ�*��=<��=X=5:3�w��ˍ�<-��=�"�=�H�>;�>��>|�=����r3>�ȕ��L�4Ⱥ=�?���b@���b���~���.��v3�ѬB>��V>}��ߑ�9�?�V>}O>>iX�??�u?�a$>.��n(־���k�e��Q��9�=��>��A� �;���_�irM���Ҿ�M�>/��>$�>�;5>�35�>W>�deŽ�t��ǌ5��, ?����e6��=�{�R�� ������h� �;Ђ
?�V��+h<8��?��e?w�?��>���z���1�>#.���8>��4�R����׽� ?>0?��>���}=��̾I7��6�>T?J��O��֕���0�B����O�>[���ŨϾ�@3��S��쨏���B�Qnr��:�>=�N?�?��]��ʀ��O�����W���r?� h?O۠>�??�ޝ�!���?���=no?���?��?5
>?�K>m���+�`>2�/?㑡?�ԕ?Rt�?�}����r>�Hf��Q?> �!>�	�>��>��k�(�`��>_^>��\>��ҽSd�[������������W=%&)=��H>�v�=�>��	=�ox��A�=�>o�@>�,>�M>ޓ�>y�Y>a���#�
�#-*?�'�=r:~>F.?|h>�Ƃ=������
=o��l3J�M2,�@����N׽�=7��5�=	Ɋ�ƒ�>iPſ�Ӗ? LX>�I�+Q?k���\�!�V>��?>������>j{A>�r}>��>6�>r�+>RA�>ڒ7>2<Ӿ�>���c!�)C�|R���Ѿpz>�����%�P��ό���MI�Q_��j^��
j�!+��<4=�I�<E�?܍��d�k���)�ʤ����?,T�>B6?�ӌ��숽��>���>oÍ>�3��?���PǍ��lᾑ�?���?ke>��>�=e?�]?Ga��k6�p;\�|Sl��8��S�8�?��X��"�r�b���A��Q?��w?־8?B[�<�"�>�?��1�����n��>�����3��V��K�>}㌾�f��lM���X��X<ͽͬ�>��C?`}m?G"?�����+A�>-N8?�W8?R}y?\3?��;?L���Y ?6v>\�>T�?ӷ8?,?Q?�>�>�8�M}<i��|���zf޽Z�ʽ+����9=�yK=��<��<���<���<��4��à���g<5�3�D�<��=_�="�=��><�c?�"?Q��>�n?��;(��h2��� >n�>�+����۾S�=��\�(j5>+�
?T�o?��?Zr?�L�3�C�p=jI�>���>o��=&�>n��<�e �f�ʻI�i=���>@�q>ӧJ���ԾU~��ΐ8��-���ͽ[:�>Fh>�f|���3>�ˢ��px�?�j>GLU�_����QU��yD��-0���t��6�>05K?�"?�4�=M�뾮�����d���&?�e<?�FM?�g�?p��=�۾�'8�<�H��w ����>q��<'�����T��
�9��w;�x> 4���ܙ�z�n>���g꾼?o�uWI�3���=){�dt=��~�̾�r��?�=�p�=4!��yV��L������+I?11i=�5���4]�������>�ؕ>[��>�4@�v47�B�>�CO��i�=�V�>'�9>�aG�/V��d^D�w �'Ș>�:?��I?�;�?���]�}��-�;���&�.�R�G�?H�?�?�F�>�	�;ɾ�������U�13�=�?�4?΃-�Q� �־���k�F�q:>G��>Msh�r��>v�^?{6+?@h?�?L��>Ns�>a�]��#���b.?�t�?p���F������?�W}Y����>de%?��n�l�=�v?��L?7^?�?�M�>a�><�;SR1�'j�>�0�>�_E�ZԴ�S�L>�3?!��=�V?HT?I�>�=�/���>>={��=���=V�5?V?�F,?�Z�>V�>y���?!>j?8�?�L�?q��?�o1=Mڻ>��M>��>[��=ф��t�,>�'0?r�?t;S?�I?L�?A�p�U8���^F�����cK>��7>��=���;�ps�ib�����۟��
t;�㱻zPJ��n�<x��Q����,�=�i�>�u>����0>BmľV����?>7}���k���ቾD9�..�=9�>H�?Y�>
P"����=G�>X<�>����'?1�?qf?��{;&�a��VپR�L�_s�>_FB?ϵ�= �l�ΐ���/v��}q=n?gq^?ޅU�je��K�b?��]?Qh��=��þ��b�щ�k�O?3�
?�G���>��~?d�q?-��>@�e�:n���Db�I�j�vѶ=[r�>JX�T�d�w?�>k�7?�N�>7�b>�$�=Eu۾�w��q��b?}�?�?���?�**>o�n�F4࿾^��tP��/N^?�>�>�R���5#?C����ξ���|Y���⾁����H������Ӧ�K�#�TɃ���׽r�=9�?ls?Kq?�_?`� ���c��0^����4qV���������E��E�.4C��hn�_y�Sr��c��7�F=9=^�kmL�K�?�?��N��{?�ӝ�.d��.k��V��=GH��`���mq�;+�ͯ����>[�Z�F�_��ھ�b?���>��>)z2?�#R�%iE��l6���S�3f	�#�I>Z��>�q>�o�>6]�=f^���|T�����2��A���68v>9wc??�K?�n?GN�/+1����Μ!��K/��O��x�B>�C>�>��W��u�M=&��R>���r���<y��D�	�Qs~=)�2?��>���>MQ�?F	?�t	�gV��fx�p}1�ݙ�<�>�i?)1�>S�>�нV� ����>��l?���>�>_���pZ!���{��ʽ�&�>}�>X��>��o>Y�,�g#\��j��Q����9�w�=#�h?������`���>\R?p��::�G<}�>�v���!�Z��S�'���>M|?���=k�;>�ž�$�y�{�*8����4?H ?ꥠ�7�.�e�S>r��>+��>5	�>�i�?�#�>�^ؾ�A�C�=?��W?'Q?d�8?��?V��=��Y�V?��U5�.����F>�hF>t͕=(� >ow�ti:�ׇ���>F�<�Xt� ɿ��G�;���=���Aj'��~)>'�ؿ�`��r�5rپ�e�����4��}�:���K߽�&�VQ��� �8Ĝ�xو=+1��
9[�a�m�ǎ��%��?���?���=;�=�����S )���l>Y����D�����f>d5�8����.޾�P�g���T�����O�'?�����ǿ򰡿�:ܾ4! ?�A ?7�y?��6�"���8�� >XC�<-����뾭����ο@�����^?���>��/��o��>ޥ�>�X>�Hq>����螾m1�<��?7�-?��>Ǝr�1�ɿc���w¤<���?0�@G�A?3�'��쾔�O=� �>��?�?>>S0��T�ػ�����>2Ξ?�$�?^P=z�W�I���e?�<��F�]Bӻ}��=1I�=��=	s��KL>v��>�U�R�A��ܽ�?7>%��>�,��k��d[����<��Y>�?ֽ����4Մ?{\�|f���/��T��U>��T?�*�>y:�=��,?D7H�\}Ͽ�\��*a?�0�?���?�(?/ۿ��ؚ>��ܾ��M?bD6?���>�d&��t�"��=Y6�q���o���&V���=;��>I�>��,�ދ���O��I��d��=� �+ÿ�5�x
�;#�$�@����<��S�V4<3�>_������TJ���H��d$>Y�#=���=��>�w>�e?k*S?/�>��>��h��q������&�X�0��U��'��=
پ���[$k�+J��<���' ���������\>��H��#���E��x��[�7�?.�=�`�gX]�Ep�>�)��!��_*.�%��^wz��px����v�?5>j?�t��Յ��u�8V�8�����#�?����!���+N��[򯼟?�>W\)>(0��B�>"�y��;&�^!a���G?�2?}���������?,��	ȓ<q�3?�X?Q�޽��?��>˂j��y����>~\?6L>���>�F><ؾU�Q���&?-Yb?-�N�y5���>�þ�p����=l3�>T�&�^d��A%>�&>��7�O�߽�� ������*W?r��>��)�Z�0^��8���<=��x?��?�!�>�kk?��B?X��<�P��V�S�3��Hx=j�W?�!i?��>F���Bо.�����5?�e?�N>�Mh� ��[�.��C��?��n?�P?g~��%^}���	���h6?��v?s^�xs�����N�V�e=�>�[�>���>��9��k�>�>?�#��G������yY4�%Þ?��@���?}�;<��R��=�;?l\�>�O��>ƾ�z������)�q=�"�>���~ev����R,�g�8?ݠ�?���>��������>Ӝ����?jy?� ƾT��=�*���?�����bC��Lz>~Mm��;�O����B������ND�m��|�R��ֆ>G�@���V?�yj�]���[¿Z���ݾу��'I?��?ۢż�D>���J����gq��NF�����>��>�諒
c���\z��q:� �漛n�>}亼�H�>��Q��G��Kڔ���<��>6�>79�>-����q���	�?��8˿UԜ��'��Z?+��?�8�?�?+�<��b��w�Ν��>?�v?T�\?$ᄽ�PY��x��j?�_��vU`��4�_HE��U>�"3?�B�>@�-�ϲ|=�>���>Sg>�#/�t�Ŀ�ٶ�6���U��?��?�o���>f��?`s+?�i�8���[����*�ɯ+��<A?�2>����J�!�A0=�2Ғ���
?Z~0?�z�W.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�A�>!�?@}�=��>�"�=ʰ�b�8�6�#>
p�=�N>���?�nM?oN�>E��=��9���.�5:F��nR�CS���C�Y��>
4b?\�L?�b>�b���J/��!���ͽ2��߼�r@�/�k�޽��4>>�=>;>�D��Ӿu�?vp��ؿ�i���o'�f54?d��>��?�����t�C���;_?%z�>�6��+���%���B�L��?�G�? �?t�׾zV̼>��>J�>I�Խp���⁇�;�7>��B?���D��i�o�L�>���?�@�ծ?Ti��	?���P��Ua~����7�f��=��7?�0�*�z>���>��=�nv�ݻ��W�s����>�B�?�{�?��>!�l?��o�O�B���1=4M�>Μk?�s?�To���b�B>��?������L��f?
�
@~u@_�^?*9�߿"졿�(־�kξ"y�=�=�U>������=�$3���l�x��.�= Ĥ>E��>�C>'��=�=6>��H>k������ʜ��䊿�=@��������[O���fEV�	�U�˾�x�;9�� ���ܽ 4T��������z�=�U?�R?�p?�� ?6�x���>����n=�"��m�=��>�+2?f�L?��*?H��=�]����d�\O��am���߇���>S�I>J��>�
�>�F�>:Ο9��I>�?>%&�>�>��%=6캝I=�%N>�S�>��>V��>�F�>�+�>�H���?ſ��o�,������Vݭ?{����s龔˲�i^�{F�%���>F�>��{��ɿ<�>2?����&���![��>�)?��?:�>r���ȿ�=Ӷ&>*y��_�l��5O>�4��,+ʽ[5�jx�=i?�m�>0h�>~E�1a���S�D���I�9a�M?�.��������s��<��ė��>�v'>��=����ġ��N��fQ���Y��}'Z?L� ?!˟��x�vX���ƾ�ї<|j=�԰>[��;�>���=-����r��qI�=�l�=���=�?�J;>��=qO�>�j���lM�/��>��1>�w<>^�??k9)?�p��Ѯ����_���u�>Õ�>�u�>���=0�_�0�=�|�>��v>WC���L���d�%n@��P>o�J��dc�`�^�'#=���C�>��#=�=�J�+�(�(=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾIh�>�x��Z�������u�z�#=T��>�8H?�V����O�`>��v
?�?�^�੤���ȿ5|v����>W�?���?f�m��A���@����>:��?�gY?ioi>�g۾;`Z����>һ@?�R?
�>�9��'���?�޶?կ�?|I>$��?��s?�n�>$Cx�R[/��6�������V=WkW;�j�>w_>B���aF��֓��h��Q�j� ��Q�a>P�$=��>2V佀5��s?�=2󋽋G��%�f�{��>},q>��I>1\�>� ?Kf�>���>ub=OX��y܀������L?�$�?3G��r����;hY�=��v�Pk?/,?�+���־-b�>@S[?�D{?{�R?=��>���,x������E��1ɜ;�`>?��>_a�>�yt�U�O>
پ��W���>�}�>� �վ�bo��@�j$�>T� ?
�>��=�� ?O�#?ij>�>	E��:���nE��R�>�W�>�?b~?V?̸�CJ3��ߒ�־����Z��(N>{�x?��?�ޕ>e���Bz���Bm���K�z���av�?�#g?)�(?r6�?c�??�oA?=d>g��F׾D���!�>"?ݪ
�%B��a'�����?e�?yw�>�咽�н/g��&��bv��r�?u�Z?�'?�p�a��þ�U�<y�7�a���<�^�c>7S>�S���ׯ=d>~��=Zn���7�
mW<��=�Q�>7��=�	8��拽C=,?ѥG��ڃ��=��r�rwD���>�HL>���U�^?tg=��{�d��lx��hU�"�?l��?�j�?Q��`�h��#=?	�?�	?P$�>�J��~|޾���WQw�|yx�w���>J��>wl�0�U������fF���ƽb��u>�>�I�>Z?!� ?��T>���>������%����!���^����>�7�>E.��M������ �>����¾R�~��y�>9N��}N�>W�
?�Aj>��|>��>�֧��=�>�!P>=ց>���>�T>��0>�J�=kZ
<1*ҽ��Q? þ��'��澺Ԭ�1jB?��e?:��>��U��c������o?���?h(�?;Gp>��h�l�*��Z?#��>����T	?��#=��t�R|A<J��x��*��A�F̏>�ͽ�8��L� ng��M?�}?��6�9�ɾYNν?�����n=�M�?��(?�)���Q�|�o���W��S����N5h�=j��M�$���p��쏿�^��-%����(��q*=��*?v�?��Ֆ��!���&k��?�zcf>��>�#�>S�>RvI>e�	��1�,^�M'�a���BR�>h[{?3I�>� 7?�y<?5�f?��E?��>�϶>�D׾�?R?'>Q�>��=��>�:?�:U?z$�>*�?��>Bv!=)���O�??<�?H��>R?@W��FC=���=խc�\ͽ)ݓ�`��;���=�꨾�����=9#>��?�x��D<��_��<�>��E?�n?&G�>E�o���(����<hC�>:�?s�}>����`p���c
�>��?�v:��*�<>A>C��=a;�KS=�>�۬���I�pL������;0���^;xe>=Y={^e=Pj�<�'�;ao�<�t�>g�?O��>�C�>8?��w� ����^�=zY>S>�>�Eپ�}��8$��]�g��^y>�w�?�z�?A�f=�=>��=�|���S����S���
��<�?�J#?DWT?ѕ�?�=?�j#?��>$+�PM��[^�����î?IC,?4��>�>�Gξ܏����1��.?b"?��c����<�'���þ�˽��>*�0�12{�˧��&F��1���#��n����?�@�?@�D�X{4��~⾹x�������??�t�>���>
q�>�d'��g����<>(�>�O?�d�>�._?^r?�:/?]}>n���+���:��k@¾���<?�L?�{�?�y�?+:�?���>B+=C��^�f�������/�=ݥW�F���>�>?��>	�?�d=W<�q��>�i���U�Q�=�Q�!~?�O?�NB?˘�>�u>D�J?�;�>v`ľ`��ĥ�\y���~���q?-�?��$?�X=����2��1����>�ȧ?~�?�W)?��G����=�y��F��Ďi�\�>&��>�>�>�=��=��>���>-P�>'�D�4���#��;�$�>�r>?T��=�Ͽ^n��T����	��W ���b�Vr�!$��Kr�Z�>�7�	�#�۾����*��r! �Y���Z���W�����>XÃ=2��=�EZ=.%�=�ɋ=�3�=e�꺤�i;~u�r���hA�=��x��k��I��:Ť��gg���>n�K>��ʾ{2}?6XI?��+?�D?�z>y1>��4�56�>�ǂ�v?��U>b3W�Z��[�8����o��K�׾Q־�`d�v㟾�>7�H�w�>f�3>2Y�=Fƈ<��=NMr=-��=ʀZ��\=�J�=��=�i�=�P�=&�>��>�6w?X�������4Q��Z罥�:?�8�>f{�=��ƾq@?��>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=L����=2>s��=w�2�T��>��J>���K��F����4�?��@��??�ዿТϿ6a/>��@>�>��T�rI7�6�i��d�R�o��%?6�9��ľS�e>+��=׾��ʾ��<��F>�cZ=#t,��0_����=\t��I�0=X[=���>x�I>��=�������=>S=pz�=�?>�����f$��"��`G=M^�=l�]>�%>NA�>�?�+?��L?Z��>��^��Od�����>&��>Aj>���=��G>#��>PC?^�? N?���>��8>�>�
S>�+��T9�3���F���[�=�{?�|?/�>h7�=yY�<� ��@J�Ι�d?��#?��>O�>����$ۿژ3�S!�t@����?�W�=��zv�<H��=n{��ӹ$�ւ�<Qf�>�z�>vt>�&c=�y>>��>H��>�B�=�60=���=��=�[y��b���GU=*gw=%߆>`n�=�.�;�h=��uJ��t�꼍Ҁ<χ$�

ü
!�=��>(Z>׬�>2��=�ݳ��@/>t����L�s��=I��)B�%)d��6~���.�Q6�R�B>
	X>E؄�4���? 8Z>��?>��?1=u?D& >�$���վ�H��A;e�.`S�,��=�>7"=�Jv;�fG`���M��xҾ��>�+�>i1�>$�[>ɀ-�4�8� �7=M׾R�:����>�_���WV�����k�h0���e��p�c����o*8?]������=P-�?�M?<f�?!�>�P�W�Ͼp�P>�Վ��=�<��䄾����)J?��&?:��>��۾?�3�̾����a�>}�I���O�J���
�0���%��ѷ�%�>\���{�о�3��[�����ÜB�!�r��%�>ͷO?�?z#b�I��O����xʄ�i?.g?O\�>�?��?�����$�����=,�n?'��?;�?/
>�->t��?s�>� $?�P�?��?�)�?$S6���>�Y��D[>��<���>Fs?>X����|Z�B])>� ?M#?;rp��"���,��>�> ���ڼ���=|�>�0�>���>��"- >��I>@�%>0�F=�KC<��:>r�d>�"Z>��h������L?�݁=M�>sU?v�>R�>z6����x�Y������i��hyV��E�>��>׃=vн'�����!>?�̿�ڱ?��>V���X2?DG����'>�)�>ci>*��Iq�>�ٹ=�,=��>�>��=���>B�s>�ԾN	>���<!��pC�Y�R�@Ѿ��x>����x$��n����`CJ��派�O��Tj����p�<���<?��?f����j��)�+@����?��>�6?��l��7�>���>yt�>X��N1��-���bᾣ�?e��?��c>9x�>��W?9�?��.�C90���Y��6v�*zA��0d�8�_�z��h���	��0��=�_?�Xy?�%B?��<NRy>�?z�%� 9���>�/�:;��G=��>�W����b�"־�o��k�^
B>��m?;̃?)o?*S�� ��#>C>?�9?���?��9?ʉ9?^� �,q?�+>�}?�	?c�?v:#?@r?e=>"#�=�g�<���=�>��hG���s��OMϽ�DR��sH=�
�=�l+���p��a=�G}<��F�ac ��-I<�*����0=sJp<G|�=PP�=�մ>��e?�o?5�z>�38?`]`��i�:o���>è=��R�wѾ�W�v�E��g�>�C?��?i�~?i�>��I�\�a����=��>��y>���<�o>��K���.>n��<�R�����8>�׼��Y���튛���=O�C>�T�>Th�>]���p7�=.|���jT���>fB�b���bX��,���1��Da�-��>�"%?X?��=f�	��0?�
�q�P�>�c?��\?֔r?�>J���O�3�XY/�I�r�m�>�R,�(��	4��yo���&,��ů<���>Ɛ���]���E�>}��b���y��P�q�\��=�@�q��;���D���-�P��=)�=��)���������O?{��=�]���1��9���gZ>��{>s�>"���A)x<:�/���ƾ�@�=��>ŉ8>}s9=��R�5��a�s��>1$:?��g?�w�?p믾����(J���ߺ���+�5�;?�r�>�?���>Z�O=];�i.��kpb��}E�>�>7?�D/�-DZ������1��0��2G=�ǐ>��A>HP?��n?�� ?
B?��H?+�>QU>�+�yD���D3?Y��?��U={�)��)J�
E�XP��?O?�E����>-+E??A?ܰ?lQ?H?.e��+&׾���2�>3�>S�A�����n!>)Gm?]�]>AJ?�F?���>�)��ܾ����ͨ�=�v>�#+?i�>-�0?Wd>6��>ԣ¾wE�<�=�>cPy?9��?���?1�>p\�>�lA>qI�>�D�=��>GD�>t��>�I?s�e?ߤV?
�?�as���ǽ� ��q»��k=�3�=T��<{�&�1���C�==��=���=�bͼ�:�<[|�=
2������ӽ��t�Z��>jw>Ǔ�_�0>�sľ����?>Tͼ�\��d���y5��B�=�}>>�?��>�!�d��=�u�>���>ċ�յ&?��?�?��;�`b�Y&ؾ�aK�Ų�>��A?U��=�Tm�lR���u��oI=1m?�6^?pS�P����b?{^?�.���<�+�þX�c�V��O�O?b�
?GQH���>�/?�r?9R�>�e�g�m����Kb�]�i��շ=���>�\��*e�m'�>��7?��>�gc>/o�=�Xھ�w�����q%?vՌ?$�?��?Y3)>�Yn�1�߿����K���]?�.�>�����"?�R���ϾQ��e�������b��󡬾R,��`Ȧ�r>$����A׽P+�=�?Dls?��q?9�_?[� ��d��h^����lXV�B��6�A�E��E��]C��n�ԕ��S���J���E@=KT��J=�[��?�0?L��X_�>7���ެ�������=5���j{�z8;z=���`=ܛ>�7��m�s�Qj��т?�f�>���>��=?}�M��tb�D�E�.��h����>v�>�9�>�}�>�8C>
1��d��+���@xB��@ӽѷy>6ta?�J?�j?�����.��+��L��mK��;�����E>=/>|�>�X�'�`s��B�JKv�w�������d�7�=��2?6S�>榨>Ũ�?�0?�:��y��n�g��i8���C����>�e?_��>Tӆ>�Я�R�����>	�l?_��>��>4���vY!��{�*�ʽ�-�>��>���>[�o>ۉ,��\��h��3���9�Ř�=�h?f����`�4�>LR?�&�:�4G<��>�;w�0�!����Ե'���>~?Cɪ=�o;>�už���{��B��:*?��?F�����)�Ysu>�� ?�g�>YA�>�2�?���>"}��q�>�Q?W�[?�SI?��9?�B�>�K=c���=�ƽ�y&�K�%=S�>��W>AKr=���=���]���$��fb=Q��=d��7ȽZ�;����<���<��3>�Pҿ5G�����N�Y���TZ����%�ʽC���Բ��:|���F ���о�Z;9(8�h�K�Ɓo�ơ��E��
�?V�@]�g��]�����ֻ���W%�l�>#0�����|ܾ<,^��{��2��6
����2�A(J��k��+���P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >]C�< -����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾r1�<��?7�-?��>Ŏr�1�ɿc����¤<���?0�@E�@?y�)��X��V=e��>�7
?A�N>�1*�`��j̲��+�>;V�?���?��Z=fW�~:��)fe?��|<8�C�Ə���E�=��=y"=����P>�G�><��~B��?ɽcsC>�p�>��+���x�_����<J]>?Cѽ�����Ԅ?Ey\��f��/��T��BV>��T? $�>�+�=f�,?!5H��|Ͽ�\�%+a?[1�?{��?Z�(?bڿ��ٚ>��ܾm�M?D6? ��>�c&���t�Y��=� Ἄ������'V����=���>
>A�,����O��)��O��=+��]A���`s�{�(���4>Z��=Bj�=�E�=f�>4�꾏�����e>���<O���� �>���>)x�>m[�>�=?AT;?��i>LH�=�m>(�[�3�bK��퇾M�u��+��:=�KϾ��*��m�P몾��������վ[�*��@>�I�y�����3�.�C�P��?�=ݜ�oMZ���=��Ҿ�����S۽�����c�!A���8�?	�u?p�g�eUb�;:L��m��Ld�>�D?���[��Pq��n�<��g>�Б>g��>!H.>�Ǥ�~�a�lea�cSH?@�6?�uf�E/��B^�x���d,�Q�A?)��>��	>��>mn�>\�]>��2��>����v_>ڣ�>b(>
~���{���?$�_?Z��\T����>����������=�!>���:������=V?|��J��*>�X����W?uύ>��)����R���d'���:=�sx?��?��>{yk?�C?M,�<Z��1�S���
� �v=��W?N�h?z�	>3���IоA���)5?�>e?�L>��g���e�.�HH�DF?sCo?�=?[���Fv}�%%��_��<�6?��v?s^�xs�����:�V�l=�>\�>���>��9��k�>�>?�#��G������{Y4�$Þ?��@���?f�;<��Q��=�;?l\�>�O��>ƾ�z������<�q=�"�>����zev����R,�e�8?ܠ�?���>������j��=�M��.��?xف?DH��g9����őE���ϾS:Ͻ|>�;��V���}���,��N��l=��ϼ��j����>��@T�i���?�����ſ2J�����}�;,?ޤ�>�+�<�X�?�a����ʴپ�3�Ι��?L�>��>�ᔽ'����{�Mu;�@<���>f,�*�>��S���������3<7ڒ>���>��> ��������?R��;:ο��������X?�_�?�n�?+_?�:<��v��{�����.G?/s?�Z?A�%�N.]���7�!�j?�_��vU`��4�iHE��U>�"3?�B�>J�-�B�|=�>w��>g>�#/�u�Ŀ�ٶ�6���X��?��?�o���>l��?ns+?�i�8��~[����*�
�+��<A?�2>���H�!�@0=�RҒ�Ƽ
?V~0?{�a.�X�_?�a�>�p���-���ƽ�ۡ> �0�_f\��O����}Xe���Ay����?Q^�?f�?Ե�� #�f6%?�>d����8Ǿ��<���>�(�>�)N>H_���u>����:��h	>���?�~�?Hj?��������V>��}?B`�>N�?O��=���>O�=尾p_@��$>;�=D@>��z?ѥM?_�>�9�=��8���.� F��VR�E:�?�C�h��>�b?��L?�}b>�����7/�� ���̽C�2�~R޼��@�|b-��V�
�4>a�=>�r>�E���Ҿ��?K�`�ؿD5��0�$�`4?r��>�S?���j�z�0fN�c�_?<$�>�!�����Y�������H�?C��?��?gt־U��0>���>�̃>�ؽ����醾H]9>�3C?� �(���S�p��}�>l��?�3@ZQ�?��g��	?{ ��P��-`~�����6�M��=�7?�.�]�z>���>d�=�mv�����^�s�6��>dB�?C{�?���>έl?��o�+�B���1=�O�>��k?�u?��n��a�B>��?�������M��f?��
@u@
�^?1�{ڿ%:���վd���;9�f=�y>I)���=���=��'��B��R>ax�>-0>��<�_E>�@q>DbP>'y���H!�1���΋�l2Y�8�&I���#���
��s��c��%E��g����(��[��<��g�J�-�9���W��P��=��U?�R?�+p?� ?�z��>f���%
=�V!�ؽ�=���>�2?��L?�4*?�m�=����d��R��?J���߇����>�	J>~|�>CT�>���>����$I>bv?>�n�>�>-�&=�k:��
=��N>���>���>`��>���> %�>�(��e���(������Vt��6Ǣ?�j�GO�!;������������{<�C�>�&�>='���	ֿ�Ѻ�� E?�ٍ���=Q�@Uf=��?7?ˡ>�W�%�a>�<�������-��>��������45����>�p�>lv�>���>߈?�T�c���v����gO���H?%�!�މ�=mH��u}�z����>O�^>�94>\�\��G����z�R�Q���N/Z?�)?�^��2��K���̾�g>R�<��W>B�A>4�>�#6��gŽ�
ڽa_���P��ه>�7?��U>�m&>�j�>�:Z�H$t��͛>^/>�܁>��H?JQ,?
/�.co�Ѩd��*$�:x>)Q?.Ȉ>`�=-�G��xo=.�>t�c>�}<��<�ь���d��1>�H��\	d��iż�t�=�����=L�!=�}b�<?ѽeP�=�~?�x���ڈ�O������mD?�I?��=�eP<*t"�����t��m��?m�@GO�?��	�وV���?�@�?J���Y��=�g�>R��>�|ξ��L���?_�ý�̢�Ƹ	��A#��@�?M�?[0������k�i�>;G%?��ӾSh�>8y�vZ��x��e�u�[�#=��>�8H?V��-�O��>��v
?�?C^�ȩ����ȿ�{v���>D�?���?@�m�zA���@�r��>��?�gY?xpi>h۾�`Z���>�@?rR?��>�9�:�'���?�޶?���?oI>��?j�s?�o�>k�x��]/�!4��������~=OhT;ф�>ٍ>T����JF��Γ��n��5�j�8��	�a>��$=�,�>���Y���n�=�����B��фg����>Aq>�I>�f�>@� ?_P�>�֙>��=��������ӊ��J�K?lI�?}��m��6M<�t�=�h���?�?0?Ů7���о�>W�[?��?�aX?hΘ>���ԭ���Ŀ��䵾��h<|Y>
�>�j�>m���3QK>�ԾF2@�}��>��>I���Wؾ�h��Y��(N�>T� ?7=�>޸�=! ?k�%?�܀>[t�>/:���!E�RF�>�^�>Ĉ�>�z?�/?�w����(�C�P���SpI���%>��f?(a&?�~�>����3���?c��5O�A�^��=x?�)?^���'��>�X�?�7c?t�/?��j>�j �W������>m� ?O�\f:���$���Fj?4�?X��>��Ͻ+ح�X�7<�A�����? fd?��'?����2\��������<T��h�,:n=�<�l��Dy>�Q >{m��”=u�">��=��x��8��s#���=���>���=��'����49,?��F�ZɃ�@�=\�r�s~D�߸>qFL>�����^?�>=�#�{�����u��M�T�U��?���?�e�?�����h�&"=?e�?��?v�>�S��܌޾���kjw�?�x�}l���>���>�#l���;���ɜ��AB���ƽ�y�Y��>ra�>��?Bx�>>�^>"g�>�E��w�&�&���{��,`��/��6�/�-�������&'��,�Ř¾ L��P��>!Ԅ��]�>�?�Mg>�y>Lu�>�p;e2�>_�F>-}>I�>�8^>c�,>$��=I�h<)6Ͻ�L?d�ѾPG'�ڑܾ1/����A?H�m?���>�Rۺ�%��|���-
?���?.A�?�GQ>�4g�`t �:�?�?s�g�ą?<=���������Q�;�D� =���*-G>2O��&�k�I�0�n�Wz?:o?�f=�3��[CٽO����o=�M�?��(?8�)���Q���o�߶W��S�����-h��e����$��p��돿�]��$$���(�cm*=��*?��?x����%��&k�?�,df>u��>��>.ݾ>�|I>��	���1��^�2N'�޾���N�>'\{?�o�>��<?=v@?�ua?TJD?>'O>/�>����?A�\>UG�>���=tG?��?>#�>�?�6?~��>���Zn��q�پ2i?��?K�?O<�>���>����g#����B=�A%� ]�)��&�>Bi�ܪԽ]��=���=�+~>L�?��8���-��۾�;�>~�E?2@ ?P,�>�"D�1>��6Լ2%�>�3?�՟>�龑~�nf� M�>��x?�������<���=��;=�ﲽ��i�p�'>9���Ӏ=��P��볽�p1����<��=�x�<GW�<�=y�=�q�<���>��?��>�g�>�x�e���B�W�=+K�>��>x/E>�ƽ�)��������U�쮄>�O�?�f�?�=��>�>%j���7Ⱦ�o� �Ⱦ��uM?��?O�:?�&�?�>?�;?~*>����㑿 |���鞾��?)B-?���>���F�Ѿj��>�.���>.R?nm��	�g�%�����c4��!>��.�!I� ��)�Y�q��������?���?\ <���њ��6ʏ������;?�D?�}>ӵ�>�d7�.`����B>D�>��M?f��>��f?zhk?4��>�9L=o
�S���0Ӽ�0����Pr>v+t?6�|?8l%?ܐ?ڢZ?lT=����9��{Ə��R��&5��􀾈���l�A>�+�>��>9PS��=:iJ�=�ii�=���R�
y�=�\.?�?��>g��> w@>{F?��>̮���b
��흾b����!����s?�B�?�&?���<����F��������>�j�?���?+?AC��1�=��������f��L�>d=�>®�>�f�=�E=c>���>���>�6�]����7�~d��Z?��C?�=�=v0ƿ�r���t��w���n<d���ݴb�����YoX��\�=,���k$�d]���_�E���P��pF������`y�3��>[�=�O�=���=���<gǼ���<b�J=^��<-�=Ak���u<LCD��&��:���{D8f8Z<;�H=��ڻ]�˾g�}?�;I?ʖ+?Z�C?�y>*>>��3�O��>U���!@?V>�P����Ѓ;�ӫ�����7�ؾ�t׾��c� ̟�4E>?PI���>�=3>=L�=�1�<��=�s=�ˎ=R�Q�V=I&�=�M�=�`�=��=��>�L>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?��>>�2������yb��-?���?�T�?>�?>ti��d�>M���㎽�q�=K����=2>o��=x�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�;>-�>)>R�%2���_���a��^��8"?��:�!0ɾI�>ݜ�=��۾��žZ9=�F5>��T=�����[����=��{��?=��j=Mq�>�:E>Vl�=_����U�=�dL=c��=��K>�Ȳ���0�[�$��V=c�=��b>ʲ">���>�?H:?[Z?��>x�������9(%���y>��>5J�>9}û�����_�>V�i?��;?�vH?%1�>"��=�\n>M��=�d��ƾ+s�ZC�1�=��?�?�H>l�u�h�U�r���Uq�w����N�>�bP?;�>KzG>�	�GP�A�A�l�"�sf����=A$.>8<�%�=�=�����6�h u=�>�0�>s>�w�>:��>6��>��>F�>�a��=�<�e=��5<Y� ��ܯ=>*x=�+p�< ���j=൮<kT��G�F�ǎ:>��=х,;<Y�< ��=/��>jj>��>��=+���M6/>������L��%�=�5��d'B��+d��=~�j/�Y
6�DqB>�X>A���d0��9�?�JZ>�?>Ӏ�?NIu?�L >$�p�վnL��Ye�H�S�!f�=L�>a�<��p;�jN`���M�yҾ� �>�Ҏ>6�>�e>0�-��e:�T7=�I־�89�m��>�]�����n�(�m��񣿮[��Wn�J���9?�釿tT�=1��?ߌH?�5�?A��>�����վ16>������:=��i�߭��?>b"?6?�>Y�ھ�>��H̾����޷>�@I�%�O���A�0�W��ͷ���>������оa$3��g��������B��Lr�[��>!�O?��?^:b��W��CUO����8(���q?�|g?"�>�J?�@?&��%z�r���v�=�n?ó�?N=�?�>kv$>������>�9?ˬ�?ț�?#�?Dp&�5�>��=Ov=�ቾ�F>ǚn>/�+�ܫE�
��>V08?C�.?0�Ľ�I��� �N�E
��?N>#��>7�g>m�5>��/>�T�=��=���<H�N>���=���=Qͫ<�%>��6>�<~�����F?�5�=�3.>X�P?q5F>��>�HZ���)�KMܻ�����Đ�yO��O�9��l>鎾|#�jU'�:�>(�ƿ�"�?��C>�$��
�/?��H��&��>J8�>I���t&>�=>h�>���>�}d>
->w�>�er>+4Ӿ�>����R!�R'C�w�R���ѾIyz> w��G&�������I@I��o���`�j�)��!3=�O��<yF�?�����k���)�8/��,�?N6�>�6?n猾�F��s�>���>>��>S;��a����ȍ�^~���?���?�?c>�%�>��W?�?ލ1��73��jZ�!�u��A���d��`�8ڍ�����1�
������_?��x?�rA?g�<�z>���?�%����;3�>�(/�;�}�>=6��>�-���,a���ӾǴþȞ�k�E>��o?g'�?JT?�[V���l��'>P�:?'�1?�Vt?��1?ċ;?����$?b3>E>?k_?	I5? �.?(�
?��1>I�="䞻^�(=�^�����l�ѽ�1ʽb���4=�|=u�)�U<j�=<��<�]��ڼ2;MV��mi�<S�9=�I�=e^�=��>Z9?e_?e?�U8?�:^�0�Ѿ>׾�*U?Q��>��m˾���ϥ� �T>b&6?7�?��H?ޠ�>���~R���>ȃU>�Λ>^�=��>Cc<`�t��r�M�>?��>�	=�M	�����(���C;=L+=��&>���>��>��3��^>�й�T�u��">�I=��GھU�|���5�\�!��n���C�>�j;?a+?�p˼M6��/���e�I{?�W?լO?��?N�>[C���.��8���j��}�>��½o�����!��
Y1���<�H�>���-(���-�>N�
����,`��JJ�\9���W;`	���<R��K�Ǿܒe��9�=�Ĭ=s��E�+����%M����U?j�=5ѵ�ie��Ӿv�=jio>8�>^J���bS2����R�
>
��>��N>[$2;1߾eL��A���r�>)�<?��R?(�?[{��,�w�M�H��=	����@:�3�?��>\�?�:�>����(��H9�� S�"���>�}? 32��Q��ǐ�-����a���J>e��>��P>��>�eg?�9?W�3?�5?���>"�>���Z���.?6Xz?���;I�n��	=� �X�3�=���>��O?U��W�>p}A?0yR?�e�>�{F?�b�>J��=˛v�hپ�5�>�׌>)tN��Y���[�<Ѕs?��<>��X?9�3?#�>1�|��8M:>P���v��=�l?"��>��D?�;�>4��>�d˾M(=���>Й�?�b�?W��?K��=h�?K;z>�#b>#�н��+>���>o�?|E2?�w�?mZ?)U?�(�<.��Җ\�t��蓽X��;i�,>��=���<�R�k7V�bm�8�B#�ҿ�����Mf��2z�<3s==���<���>i��>���C�/>��ža����>>u������L��\$�D��=���>�?�L�>�|"��(�=�ɽ>
E�>�Q��%?\A?�?���8�\�%4Ѿg�Q��Ѱ>��A?C�= yl��(��ht�A,\=��n?Y\^?ݍC������b?��]?d���H=��Eľ+c��~�`�O??�
?�I�Z�>��~?��q?�]�>Xe��/n��!����b�
�k�E�=|�>�g�e���>�7?&-�> �e>�t�=��۾�w��@���?�ʌ?&�?��?V�)>q�n�U������#^U?���>(ǘ�_�"?��<��ξ�N��\�����澺0��cؼ��Ƥ��m���!A��돾nӽ�z�=(�?R|?H�s?�X?P	���<b���f���}��P����F���mD��A��]A��q��������&����R</Dk�m�V�)�?! ? �X���>���G`��ㅾ��.=����b	r���g<��E=��=�(>"�>�rp^��9��ł?Lq�>���>HS?W�b�^�F�s]@�p�R�6�ľ��D>�*�>&�a>��>�{T>P�d��4:�:��9�z��捽?8v>�xc?�K?�n?3r�W*1�������!�&�/��b����B>n>㾉>�W����U:&��X>���r�����v���	�֠~=F�2?�(�>9��>�O�?*?�{	�Fi��Rnx�`�1�A��<�/�>Y!i?�A�>�>��Ͻ,� ����>l�l?	��>��>	���_!���{���ʽ�9�>�ԭ>'��>��o>��,�\�qf���|���9�w��=u�h?H���
�`�7�>OR?��:�cG<�r�>�v��!�����'��	>�z?���=��;>�~ž�'�M�{�	7��?�#?��?33g� �*���A>�� ?_��>>#:>4_r?�H�>������V���?h�c?�ON?�xE?ذ�>MN�=Z���x�ҽ��!�n�;�U�>�>���<ܸ�=f����Q��Yν�Ͷ<w�C=�ꋽA�'�L�z=���%��=�6�=��>�{Կ]�?��vʾ��gq��@�ܾ�u��o �3��O���ݾ�$����̾���������s�˾6����C���|�?@*@�AS�������L��9>˯���ǽ�B���������ǰ��Q�>�CdR�ܐ}�}���P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >ZC�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾�1�<��?7�-?��>Îr�1�ɿc���}¤<���?0�@�tA?a�(���쾳�U=+��>h�	?}T?>�1�I4�l԰�F@�>�2�?��?��O=��W�?^
��ce?�f<�F�?L�G��=>��=�k=�����J>�f�>���-}A��g۽�4>F��>)�"������]�a+�<g�]>�Խ�C��5Մ?+{\��f���/��T��U>��T?�*�>R:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�߅�=j6�艤�{���&V�~��=[��>a�>,������O��I��U��=�f�<v̿�Z�����_m>fT�>�z->5Ӿ����h�>���<<�ƾP���G��M �>¹?���=�
�=2�>-G?z=?eg�>�>���~RL�������⥾HR��X���ļ�ŧ����H��������6��#��Ɔ޾�)�Ջ><�I������I
�mll�Y�q���>�i�=��x�K�nz�=�.�A_��}L�V����'�җe�m���2J�?
�,?���M�Y��L��ǘ�m_���ځ?��T���0���3>�K%>>�>�|�>~m��jlj��T�1�K?;j4?�6��:e���>�:���5���>+?��?������>Jq�>/�>�"���Q>X�(��h�>�3?�'>]�����H��>��^?뽄0����>#'���jH�V@Q��t�>�.�����7�>�j���
��3� =���;�W9,W?��>b�)�V��V!��,`!�H 9=M�x?��?$m�>Ek?�B?�ȹ<���}�S�j�
��v=�W?H�h?l�>e���о�����~5?Sse?e{N>8�g���龔].�]����?�sn?�>?�̟��<}�l㒿)��f�5?��v?s^�xs�����J�V�g=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?�;<��T��=�;?k\�> �O��>ƾ�z������1�q=�"�>���ev����R,�f�8?ݠ�?���>������k�=�w��i��?"�?�*��X��>���K��{����𽮨�>�s� |�����tO�_���-7&���ξ�	3�b>m0@�$��7��>8㎾6Ϳ��ο������������5?�"�>#�.>�M2�Yd������G��X@�4�@�i[�>ͫ>���J����{���;�g�����>;��;��>�#T�����N���M,<���>��>��>xⰽU轾�ę?F<��)#ο|���S���X?7*�?���?�*?��6<�w��|�'���F?ss?�%Z?c�&���]��u8�!�j?	_��LU`���4�VHE��U>�"3?�B�>�-�2�|=�>��>�f>�#/�J�Ŀ~ٶ�����V��?���?p꾚��>���?hs+?�i��7��	[����*�Έ+��<A?�2>K�����!�,0=��Ғ�̼
?w~0?mz�i.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?���>��?���=/m�>��=�{��="���#>���=�F���?�dM?���>���=i8�:?/�#F���Q�*��)�C����>��a?	�L?� a>�B��W�+��� ��c̽e�0���qoA���-���A4>�a>>ӷ>uC�
{Ҿ��?Lp�9�ؿ j��!p'��54?.��>�?����t�����;_?Rz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?\��D��t�o�x�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?rQo���i�B>��?"������L��f?�
@u@a�^?*��޿�%����׾�ž���=6��=#�D>N��YU[='!&>�AJ=D�&�_�=�P#>u�7>��n>J�$>��3>��/>�R��3<�9U����,�+�/��� ������M�YtP��G�T���I��݇1�u�ͼ(�q�w�7 |��M�	��=¯U?aR?xp? � ?*x�x{>ɼ��	=�p#���=1�>�i2?g�L?x�*?��=L�����d�EU��@D��!���~�>�KI>>z�>D�>�&�>���8e�I>N-?>k��>�� >�d&=:���=�O>�S�>���>퀺>ߜ>Y�>kt���һ����
;��%.��	R�?rդ��U|�����X<�!X�qW�
�E?w��=�h��Y�տ<v��z�D?{9��*��G�b�X
�y?g��?���>�qѾ�,�=QQ=+5�<v��j��=���
��<2ﹾ�	?|*>S��>�I�>��:�XoT�v���Ҿ��,>T�U?n�����A���}�!4��[�+�>1ͱ>F�<�a"�c	�����^X���.���E?��?�픽o�̾ ���ٛ���|>��>�&>d��=PT�=� D�i�[�=^=I��=H00>B?��p>q� >��>�Ś��r���r�>J�O>�J�>nI?:�'?5�����/\l�7�����>��>љ�>o�>D⧾~-��8�%?�u�>��x��<�=��ɽߗK��+>++f<eT��K�y�3e6>�� ��H%�\#�=������+�Z�$��~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾRh�>sx��Z�������u�]�#=N��>�8H?�V����O�i>��v
?�?�^�ީ����ȿ4|v����>W�?���?f�m��A���@����>;��?�gY?woi>�g۾,`Z����>ͻ@?�R?�>�9�{�'���?�޶?ԯ�?�J>��?�s?��>���
,/��賿�u���ǉ=�����>�V>κ�\oB��e��=ш���i�D����`><,=c�>�W�奔�f��=N	���e����p���>�2v>0�;>S��>�?v��>�˛>��= �����:@����L?�;�?����]v��E��N=�\[��?��%?�C� ��L�>�YR?{%x?�[?��>V������gÿ�����:;�\>Q��>VE�>����JO>,�Ծ��e����>7�>Iͼ��߾k�6�_b&��y�>m?N�>�p=s ?;�#?e�j>�w�>J�D��s����E�R�>�&�>��?�;~?�?"����2����}a����Z��L>�~x?�?�z�>ڦ��蕝�{���b�>�x���5U�?�f?��ὅ�?��?�b@?�V@?;�e>b��ՙվdl��3�>,�!?�1�ζA�-�&�@���?��?�Q�>[����ս:��4������?~\?�2&?N����`���þe�<9�*��=/��j<F�J�Ͱ>#m>5\���=��>=@�m�/k7�a�<޵�=� �>D%�=�'5����;,?��F�҃��#�=P�r�'|D�w�>z?L>������^?�z=�l�{�^��u���U����?���?�j�? ᴽy�h��=?�??�&�>�X���t޾����w�=�x�Zq�0�>^��>K�m���^���ޜ���C���ƽ6���q�>l��>N�?���>�lM>��>
󖾌&%�Ǔ��~�^���7�k|/�@>������l���_ž���Z�>������>�5?�}f>��w>}3�>��ٻ.c�>I%Q>�s�>��>�jT>S�5>�\>��<}:̽�CR?<�����'�W��i����0B?�Rd?���>�xi�}�����?���?gx�?�v>�ph��+��]?eN�>s��t
?M�:=�i�ɏ�<4���n�"����Z�T��>�ֽ�:�oM�Ukf�N{
?�G?a���YU̾�ֽ�奾
�=�u�?�!?�j#��O�p���X��DP��2�+@{�%"��J�"�0�n�𜐿$I�� ̅�C7*���;3!2?�U�?d��c�-���2jn��D�\>k4�>�j�>nݼ>u>Z>l��K�&���U��$��������>�(p?�>	\*?��T?]�q?�F+?r.j>a��>�����?��׽�l�>�"�>�@4?wB?���>'x�>�$?r��>O�=Wn�ʂ��?�X?��C?�<�>���>�ʁ�#tv�r�g��)���?.�<c.��Ż�L>:Ky=v�1�nX>���>H�?�����7������f>�*5?5��>���>�]��P�j�n?�<ox�>�?�4�>� ����m���B�>�h�?;���B�=��>b��=��k�@�u;���=?��H�|=�t��� ����:U��=�#�=�6�j��,�D<�Cv8g�G;���>��?���>�ŋ>����w�/U�KЬ=��`>N>��>��վ���������f�b]}>���?<�?v"t=^��=���=-���P���E$�����<�(?�z#?b�R?�y�?3>?pH#?��>�N�P|���8��4���Ke?İ/?lq�>,��Ew����G2H��T�>1:#?�ш��*�J�)���w\�uW>����^��?����J��甾�<"�4�A�?vʖ?�Ԕ=�r�����>��.r��r(?���>qׁ>���>ܩD�e�P����e>)��>��O?;��>�[?��c?��?�u\�<�־m���ԝ��;B�$�9>u�.?�.l?ub�?�/�?z#_>���=�ȕ�S־/K?�!ѻ�
Ύ=�~f��S����a>��>���>7*>��q���>=�]����;������|=�82?�a?��?���>�#�>QI?���>�쾾n������m��sn����r?�6�?D(.?�Ɩ<�S�˪+�q��ܬ�>��?z��?�T1?��9��8�=�X���|��d0��tѳ>�y�>P�>i��=���<�W>�w�>!��>�l���=9��V'��?gD?l2$=�˿�}|������m�=��d��A@�,��"Mf��f>��r�pm+�J�ž�����꓾��~�_$���_��C-]�U��>�s=�c�=qL�=��=Էm<�f�<؁2<��h���<.w�{?�������ͻl�V� �h=�q<�U<�(=�˾W�}?<I?��+?V�C?��y>e=>̔3�ᚖ>����@? V>`�P�ɇ����;�M�������ؾov׾��c�Oʟ�}I><ZI�7�>i93>�H�=xB�<��=s==�R�=�!�=vU�=�k�=��=;�>_X>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>ºB>�>��S��05���s���h�XZ��5%?�a;�g̾��s>�6�=m�ܾ�z¾��R=H9>>:7=�p�ն`���=�燽�_=��=
;�>K9>q�=^<��=�=��=�%�=�wK>�u���xa�|�$=M��=Ci>��>��>�?�8)?eO?�+�>�7l��ؾ'O�;��>�W >o��>&*�=�<S>�.�>�C?�=>?Y?^M�>��>�ި>VV�>�&&�iG�v5��q������<_��?]�}?��>������� p��G�-���8�>��1?��?/�>R&�vZݿ��=���'��O�;���=��o=�����j�.�<>��$��%z��'s�`V>q?��>��=>�[�=�Hc>��>���=�ʥ=�S�=�[̼#�����a�<>���=j���du�b<��:=����@�J�u|��xs <+	��ح�����=nS�>��>���>��=�³��T0>���)�L��=Mা��A�69c�gg}�HR/�ql6�J�C>L�W>����1T��ee?9�_>{�@>i��?œu?�3 >v�@Ծ)ם��3e��V�k�=d�	>.=��x:�S�_�GjM�}Fо!��>�`>�ַ>�1�=m�7�n�1��J=�ⅾ�#f����>ாo��<? ���X�RY���ҋ��U��
�y�>A3��߼����?�Z7?v�?�?� =5����ˠ>��O�E�<+�]�%���K����?��+?x�>�Ծ�y���H̾���޷>�@I��O���g�0����ͷ����>�����оH$3��g������0�B��Mr���>õO?��?z9b��W��>UO����1*��hq?�|g?D�>�J?�@?�$��gy�5r��Lw�=��n?���?=�?R>�k�=�Ԉ�T�?.?P?'��?O��?sP�?L}�b��>%��>u�'>ӽ-��?���_��T��=�7G?{Z8?o?��<�����$�+�M�伹�*>�r>�m8>-��=�7�>��<|F�=�Z��1۸=>>ň>��>���=�H�=U�z�y&(��]?!#o<�+>�3?6>+z�>����,Ͻ6����O˾��%�C�û�[̽�XF>�t��������ｎ>(�ÿz�?)��>v	;�3?��� �ڻ��0?*�,<M�=��>L�=ڷ�>�#�>X	�>�1W>B��>�s�>AӾ��>���F`!��C���R���Ѿ�z>P���d&�J��������H�i���o��(j�s1��B=��U�<=O�?)2����k���)��=��9i?�>%6?۷���$��T�>^��>���>c.��T}��4���H�'�?��? @c>s'�>*�W?U�?ߑ1��3�tZ�ܱu�%"A���d�"�`�Eݍ������
�/�����_?��x?<wA?B|�<�*z>���?��%� ����6�>�$/� ;���<=�0�>@'��Pa�s�Ӿձþze��=F>܈o?)%�?�W?�LV�	(l�((>�:?\1?��s?p�1?{K;?�#��$?�t3>ya?DE?[*5?3/?��
?��2>���=񯕻R�,=2̒��Պ��9ҽ��ɽ����2=�{=f�����
<�M=�j�<K���5⼁˵:����]��<�==��=`0�=��>Y�V?��>���>ț?軾�1$��_־��8?��<������� 2p�=����>hX?���?@�P?͙�>�L�� ���-�=c��>�ؚ>��K��R�>G��=�#>��򽜳i=�q�>�i=���q���ﹾ��������b=���>t�{>�B��F%>yȤ��{�'�b>��M��ｾYS�h�G��0�(Jv�[�>_�J?GA?# �=��������f���&?;�=?�M?@M�?��=0پ��8��H�f,�j��>��B<$��W`�����8L9���*���r>��E(����^>Jr�r߾��n�S�I�g�4F=VS�ھ_=+��Ծu�~����=i> ���	� ��	�� ����'J?3Yq="ޤ�v�W�pM��'�>���>=O�>Kr+��J{���@��Q���l�=�|�>ɏC>����ڌ�b�F�ts��6�>gX=?(�`?KD�?�����2z���Q���$L������ED?+)�>�r�>�h�>&�4����c���-Y�L5���>֝?a'��TA�]�-���>&�ZhZ=��>�5>K�?�V?q]?f�l?��?o��>3��>CM:�Lξ�M*?\ׁ?ֲ�='F��<�>�1�z�L�.[�>/�(?+�ν���>���>k
?b�(?��N?��>��>�žȞ��4o�>�>4�M��E����%>@#:?��M>x�L?�G]?�&�>��7�9Y뾤n����K>�=�{?�?�c9?�Y�>|��>��c�9,>��>�O�?;h�?�/t?�`L�-U�>0�>�x?��A������۶>�`?�/l?�)o?�(H?���>r�û;����ܽ�)�<+n�=�!�=�u.>��>j'<R2P��W��#O'>%i�=����[���$�Lv�=���=���<S�>�M�>�j�)f�=�ԾD0p��~>�/��(��Hm�A!ҽ��=5��>u�?��>s,��Ƴ=�ݽ> �>s��F�?/^�>�R?O���!�L��C������s�>.XG?_�Q=_�g��/��\\��W�=��d?:�|?��_y��b?�]?j�=�+�þ��b�ݏ���O?o�
?��G�w�>�~?�q?���>(�e�C9n�����Fb�k�-��=�v�>+\���d�V>�>s�7?JG�>V�b>��=�r۾}�w�4t��O?��?� �?t��?j!*>��n�c1�^���aP����]?�}�>B7��-�"?������Ͼ!=��c8���)⾈&���!��n��������$��҃�\׽��=��?�s?iGq?B�_?�� ���c�r2^�o���lV��1��2�8�E� E�W�C���n�M�<�������F=�IU�@MG�¹?f(?I��TT?����F�/�Tt��iB>�ԣ�����>�G�Ŏ�<�ވ>�?��E���,����?{6�>C��>7QE?>�=��7���H<�ed��o�==��>+-�>��>S| ����F���{þ�W�B��� �w>X�c?D�K?V�l?>8����0������(#��Q��:Ҫ��T>��>=J�>˒A��� �ұ&��E>���q�E����������=:�-?���><�>臘?�� ?<���%�����,�E��</��>�-j?���>Ac�>��̽�]����>��l?-��>y�>�����Z!���{�V�ʽv#�>�ޭ>ɸ�>_�o>h�,��!\��j��#���y9�vr�=�h?2�����`�'�>mR?�Y�:K�G<5~�>`�v��!�����'�Q�>�|?7��=�;>�~žy$��{�%7��QD7?&/?����r-�+IT>qS�>�1p>}�>�ƌ?K�>vΘ��-N�
�	?-�a?��E?�V?�q�>���>$�=oh��|��"}�;��>w8>a��=�N&>�a��ʼ;"����y�=|�=�^����$�=I���˙���$>i��=�6пA�D���߾P=�"	�@|$�#p�J���\��[��>o��w�,�{�v��|^��ޯ�򆔾t>j�����z3n�fR�?��?�X]���|�,L��D���Q" ��S�>����ݤ����ܾ�O޽Ɛn������b��3��r)�Μw�%X��E�'?�����ǿ𰡿�:ܾ,! ?�A ?-�y?��(�"���8�*� >C�<w.����뾩����οJ�����^?���>��t/��m��>ϥ�>��X>�Hq>����螾21�<��?1�-?��>��r�(�ɿe������<���?.�@�sA??�(�B��-`V=k��>��	?�1@>R^1��<����Q@�>3�?6��?[�M=!�W����ve?7�<[�F��߻���=A�=a�=��UfJ>�`�>\c��'A�Vܽ1�4>�˅>�c"�{���j^�6߽<�T]>��ս�Ҕ�5Մ?,{\��f���/��T��U>��T?�*�>T:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=y6�����{���&V�}��=[��>c�>,������O��I��T��=����׃Ŀ��R�!�E�s�=�齑d>�e��L��(D�=�Go���o��c!��z��m;x�>f�6>�t=�L�>�\5?�vG?D�>(�;6��b��?7��'�,/�0�Q>�h�=���;�哾����ۅ;`N��������
�2� �/�K>��P�DS��-�>�y�}��J��?�@>�~���;���u>��/�@K=�`�׏��&KP��a��}�?�Lx?Jˏ� P����1��>⭜��yY?vJ���S(����5}H��]=�w>�w�>��">_׿�Ejp�o	��9<?�v0?� ����?":>�������sH<?�7?��=w�>���>-`߾����h�>��>R�D>��?uE�>V>��3G���$?�QY?!��:ݝ�+�>�>۾�P���5>C�[>�`��?�
��=�U�=e|	���=�!j���ǽ�V?Ɯ�>��)����K&��@��t�G=Xax?1�?�B�>0�j?��B?O̡<�Y���S�1��ey=8"X?Z�i?�+>�4���Ͼ�y��K<5?+�d?�jO>��e�i%�@./�p���?sn?;?RŘ��"}�]��ZK�\t6?��v?s^�ws�����>�V�m=�>�[�>���>��9��k�>�>?�#��G������zY4�$Þ?��@���?��;< �J��=�;?k\�> �O��>ƾ�z������=�q=�"�>���}ev����R,�d�8?۠�?���>������<h>ح�����?䏆?�.�����?�b����8��B���V>� �7�8<��BK4��|���-���վ�5E���>�3@z�~��b�>0��	��l�Ͽ\A��bߴ�8��4�I?Ξ�>=�ž5O�=��T�K��G�'�� �[�R���>�{>�K��A蒾��{�@,;�p"���'�>6	����>UT�ґ��K%��|7<[Ւ>]��>���>$ڵ�B/�����?����t
ο����&��mY?\�?���?9?�3<1�w��6}�����F?��s?nHZ? ,�t	]��77�S�j?�f���S`�Ћ4��AE�$U>�'3?sG�>	�-� �|=j>���>�_>!/��Ŀ�ٶ��������?k��?l����>v�?Ro+?�j�8��e_��#�*�zA"��;A?w2>����X�!��.=�ϒ�x�
?�w0?;��b)�]�_?*�a�M�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?ֵ�� #�f6%?�>d����8Ǿ��<���>�(�>*N>aH_���u>����:�i	>���?�~�?Qj?���� ����U>
�}?	0�>y�? l�=�Y�>l��=����`�>��=��G�7�?��M?�0�>D��=�:�P/��6F���Q�E%�mC�mĈ>^^a?!K?�[f>#����V���!���н��0�����D#=�a����ݽ�7>��>>D>�#D�yҾ��?Up�0�ؿ�i���o'��54?g��>!�?��̴t�����;_?Kz�>�6��+���%���B�^��?�G�?8�?��׾yR̼�>"�>�I�>}�Խ����L����7>-�B?J��D��]�o���>���?�@�ծ?_i��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?oQo���i�B>��?"������L��f?�
@u@a�^?*�/ֿ0��P�׾�^���5t=��<A�q>҂ �}/�=�_� �нǬ4������gG>i��=�Ҁ=�
^>Ba >��=s��%Q��錄ժy�8E����=�����t���x˾r9�������iԣ�qz���н�(^����$Ǵ���=s�W?q=T?WOg?��>ߗ��P8>���^;]��RG�� >��>;�;?��R?�!?��=))���8_��y� f���np���>q�>ڧ�>��>���>J�w��?>9+>bS>c>���=@���?�=2�N>���>��>�V�>�þ>�)�>�I��p�Ͽ�	��e���Gɾ怣?�*�SW�J
��hH�����:��=�eK?��>�
��mͿ�jĿA�I?	������h u����=7?�0?�#�>1A)��">�Re�c�hP���=�+�=�L�=E�a��=�=��#?Ēl>��v>��4�0n:���Q�^���r>��6?Ԋ��N�8�3w���E�w~پ��M>���>diE��O ��j������i���t=Q�:?Fs?����1:���x�^����.J>��\>;8=?��=H> T��ҽ��I��n7=��=��]>��?f6>1��=�C�>�*�� iW��<�>R�5>8>&�??7$?�%P�k֘�Gfs����!*}>N[�>�d�>X�>��E���=���>�k^>j!�)�������A�S�H>^Z���P��P�s�{=����wl�=]��=���w�I��\�<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�3�>5���Y��B����u��#=2��>�#H?�Z���iN��=�o
?&?���Z���}�ȿ{v����>
�?��?�m�y5���	@�qj�>y��?�[Y?��i>�A۾ wZ��k�>z�@?p�Q?O�>i�:�'���?RԶ?a��?��L>Pݐ?�s?���>č���=1��㳿{O���f =���Я�>��
>�κ�l�>�q'���}��c�i������V>Q�=C��>y��+5�����=n�t����6#��2l�>�s>��C>��>3�?� �>3�>_Y&=�?h���x�������\?a9�??�1�_S��f}��_)=�1Ǿ@&?��?ړy�j*0��p�>�#`?�d?��h?��>H�D�_ݩ�/������b���x>��?�G�>�{�>ּM+;>S���b>%D�>�">"����8�_�O�/�:>ڏ?���>�q=�� ? �#?��j>�4�>�`E�d9��|�E����>ip�>�4?&�~?[�?�ܹ�1I3����j硿u�[�N>O�x?'T?J��>V���;���YE��4J��E��?��?"pg?l.彩?'2�?{�??��A?sf>@��R�׾�T���Ҁ>1"?�<�x�A���&��0��?�q?���>1�����ս+ �p�������?̈́\?�L&?�����`�dq¾N��<�e0��S;<�E��>�>`F���=�j>؟�=��k��78�)�a<&��=��>�g�=Y�7��3��0=,?Q�G�yۃ���=��r�;xD���>�IL>����^?`l=��{�����x��
	U�� �?���?Yk�?P��?�h��$=?�?U	?p"�>�J���}޾@���Pw�~x��w�R�>���>;�l���G���֙���F����Ž\�5����>`��>��?<��>�`A>�s�>,2��pX&�1Qݾ�j ��R^��:��;��/�r��������:��Nb;=����*t���>�o���^�>S?�|o>{�>�z�>LH|�^Zz>r�>>��>�K�>k�>j�3>lY�=�nw<UiӽS�H?#TݾB�"�~`ܾ����7E?�.w?5	?�T�������!���'%?3��?�͖?B�x>*Ko�z��\?A�?�qc�}?O�l=Π��w7�`�̾�Kz���̽��W<���>��ǽ�3�-�R���j�8j?�>?j�e�'vǾ~ȋ��{��o�=�R�?��$?!�)�JQ���i��=X��R�b��kS�H朾��#��qu�����X�������(�L\�=�)?$.�?�{����)ί�H�h���;���p>2��>hq�>a�>��@>����|'�!�S�$�-�W��B��>��}?
��>.�>?�FJ?��P?��7?hV>��>s1���?E��>L۟>ɝk=j �>O�3?-�>?8�	?��:?h0�>G�½�B�Uw���w�>�N?T�@?���>��>0�b��\��JՍ=X��=����
����" ����=>��=9���a=6�?%el�3a2��۾�v�>�<A?��? ��>�;5��!þ+SO����>3V�>�u>j��[��И����?���?���9<[;�B%>��i=6���oU�G�==�t�=p^�b*=<�JP=��C=o��=B�T=?��;BU�?酽[,%=�t�>9�?I��>�H�>5���� ����c[�=6Y>7S>{>�Aپ�}��.$����g�p[y>�x�?�z�?%�f=��=y��=&}���Q��������� �<ͣ?�H#?;TT?쓒?�=?�l#?}�>+�iN���\�����`�?_7?�>�x��`������+�"V>�?��b������ �@����Ƚ0�l>�2��TF�YF8N���m��l������?M�?�v�'$��������0����zF?�?X�!>zâ>���s�A]?��ӥ>�`?vt9?_��>P�b?Q��?�,?&8>]���S~�X����n�
�$*Z?I
�?,�?b�?,��>d�½�������E(ʾ����<�齁��*	�<���>ε!?.�'>9�E>ᚼ�]�g� ��~;>��<>�;?i��>�>�>���>և�=v�G? ��>ｾ!H�Aꢾ�f���C�e�t?�F�?��+?t=����nE�����3��>	��?^ͫ?�J*?Z}O���=��м ���
�r�(;�>�W�>Gə>�S�=6�J=B)>���>�`�>%�����68���I���?u�F?`.�=��Կ�񒿆�k� �I�_����*{=+����'���>1��4TS�᝾�&�l�%�������Y��;s�E=���>	>S2*=m=��9�L
�^��;b��=���=��B=Ѕ=>�˺=qy�=�R�;�e>/ۜ=z�?=�N-�``˾D|}?�?I?`�+?M�C?&y>,>X4�V��>�,��PF?��U>�MP�o]��{5;��h��C���֣ؾ�q׾L�c�"��� �>�EK�%s>�=3>XI�=a#�<TQ�=	{q=}�=�)2�C=���=�~�=p�=Zv�=݊>V>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��7>VG>��R���1���\���b���Z���!?�/;�-̾�%�>!��=߾C{ƾ�9/=�6>Hb=�?�O=\�m�=�z���;=T�k=щ>7�C>�z�=���&�='�I=��=��O>1��Ѣ7��+��3=A��=��b>�%>T~�>��?ߴ5?M?8��>ֆ�y2���? �`�>Ħ�=��>3��=]�K>fE�>��@?I #?�R?xz�>��\=�w�>�v�>{v+�F�P��ƾ	��������Wv?�U�?���>�L޽ �@�\����m��M �>��(?��?oƺ>t�����8�*���(��'�� �Xn=�1m�W���f0j�$/��f��$�=���>�s�>3Ǥ>��x>\�5>�JY>4��>9�
>r�A<{�==�s;��@=��]�r�=k�/�:�<{�/�Z�<��#k�X��D/�� �<	�!��<w� �NC�=�g�>%�>���>ˋ�=3����e.>����ѽL�?I�=�e��qB�.)d�u�}��.��`6�piA>��V>�ᅽ)���Y?b[>��?>ݴ�?VXu?�P!>D5�<�վk=���,f�2�T��!�=_>�z<�f�:�AA`���M�cҾv��>��S>Q��>�`W>�fF����s���N�~A��Y�>�U[�L��B{k���&�0s��}����Bi�\�$���>�`��B�,����?]�N?�N�?�
?��3>ۑ��te>z���qx��w�l���'��-Y�b?l�#?�
�>i������ݾ[1��>P�S��O�ԓ�X�$�!Kü������>9����n;"0��t���`��M�G�D���#j�>�tY?���?��G�	�t�t�J����������>�.j?oV�>3�>�4�>���@��(�0���3>��^?s �?\��?8 �=q�C>�w�mN�>[�#?�A�?�?,�?�����?(y罀hL=5e�=LU<�Ͻpi�񚀾G�[?ROh?3�"?mｴ����	�о,��E9�?�=J"�>�т>�l	>i�%��D=A>�g>�F�=�˽Z�=�ݰ>Iy�>[���8��X$0?e�=���> 2?,�h>!>�|⽜�z<�F��vq��?c"�E>���Ž>�=�sN��F;�S��;�>�Eſڔ?-^i>a�վ�>?�+ʾe�F;!� >�H>�	��V"�>��>>���>���>l�>*��>�"7>5Uؾp7>U���� �~�B�R�l�̾��n>�a��H���'�+}��6K�lJ����o,i�fՁ�1B=�~=8��?�n��i��4)�{���?���>F�6?t����-��<Z>C��>o�>[���)��[7��G���`�?��?cDc>�4�>	�W?��?1�1�}3�lZ��u��A���d���`��׍�����<r
�$@��/�_?�x?�wA?4�<�&z>���?��%�Í���S�>�/�9;�Y==�e�>x���a���ӾI�þ�9��%F>��o?Z#�?�^?�OV�ȼ'�=>e�??r�K?��l?�'?M)?�R.�n�?;j?>c�?���>H}%?�$?��?M�o>ٙm>Nc����ݺI��:�U�Y�'��zM� ���X7�=p�=������l���C��2e=�>�=t*=.����M<L�e��P�:��<q�J=h��>L�K?�L	?
��>2t<?����6A;�x4?Ƈs>��ս��վc�Ҿ5ҟ�Qce>H�e?i�?cQI?0=S>��7�+X���=x��>Ŕv>f2.>c��>�D��_���q<�q>�lI>�N$=�8 ������в��Nx��ۋ�=Q0�>3~o>Z��g->�f��k$a���V>y"$�^w��O�D���C�\�8�Rrv�˂�> K?�?�tf=�/�o����d��F?HX>?":O?�ׁ?��=�DƾF�8�[�N������>��-<<��)���9���	(��*D<u]>�៾PꞾ��b>h$
���۾\nn��{H�B��~�X=aC��>=���)־��x�9�=o�>�\ƾ�O"��疿�����I?q�{=����&U�b���D�>�v�>b�>�G��䈽��>�5W�����=^��>��=>��S� ���H������>M�A?��Z?�2�?����^i���@��Y�5���U��E�?��>"	?׶>>���=PlѾ%��}�f��>��P�>[T�>f���kE�ߵ���7 �"�]!o>c�>R��=�?Z�H?��>>kQ?M.?3�?]�w>*��޾�M&?;��?/�=��ٽT�Ҽ8�J�E�T��>@)?��C����>��?�?��&?Q�Q?0�?i�
>�$��@��6�>_��>��W�b��
b>k�J?o�>@�X?�Ѓ?�?>?6������7��Ì�=kU>�3?mN#?��?�ݷ>I��>O �=����=��b?6"�?�ܐ?5@���H�>x�>��#?��>u�?��F?F�P?fi?��Q?�-?.Y?�= �d�`�|z��\p���"��Ҳ���78>����5J��K�<�0���Y'�����/�6<�A=U�=햨�G7�>�s>���ӌ1>�iž����B.?>Jؗ��-��ͅ����9��X�=�E�>~�?�.�>x(���=�/�>h�>tP�a>(?I?]�?�;�b��۾�L��կ>��@?�f�=&�l����=�u��l=��m?*F]?�Z�mk���[?�@]?J���2�c7Ҿ�Pk����/?���>\3Ծt#�>�l6?yvZ?��>��m��
j����@����jʾ�>!��>V
-�k���A�?j�?�>�G�=��&>�����6��������>|P~?}N�?D�? <>O����������O���d�U?�M�>Y����?;�Ѽ�2ܾ�衾�$������e���戬��g��6�����Խ�[�D��t:>9?�x?��f?'�^??
�p�r��d�4�o��R���|��JE���S�PjX���t���:�ξF[w����=
�z���H�`�?��-?��a��g?�C¾����@辔�	>K	��7Ғ�c��<���8��<>I=�nA�e袽���Q�?��>��>��/?�`�ƕ:���(���4�U���J>�r�>�@�>��>5N�<H�g?���Ⱦfx�����4w�>!N?�U7?Y&w?םG�����l�=@�ξ��7>�5>�>I3(�~s��S���M�D�]���ľ�n��>I+��D>:w�>=s%=��?��?��>�4[�,�F��t�k� ������u?���?�Η>w�>h�������>�ل?���>�A�>ߨ��t:�����M>�[R?*%=9?�e�>7=	>eY�����c�����a�L�=L�V?Wlv�5Pþ�
{>�n?`Ȝ=���=x�>�9{�0)��Ҿ�$���Y�<X�>�G>&�>*�����꾨uT��J���A)??*?�撾-}*��>�0"?n��>ݟ�>��?��>ZKþ�{����?V_?tcJ?�_A?�&�>��=�5��Z\Ƚ�&��o0=�އ>1�Z>>�l=>�=���\�
����C=���=AҼɹ����<�����T<�6�<�g4>g�ٿжF��Ӿ�D�+k�V
��,W��(��aJ���پ�ܭ�.ώ�ң(��ڻGy������W�yg�j��?a�?:z����c�/o��Ȏ���	����>��W����<���ծܽ�vоV����޾{�$�ܺ/��BO�wS�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >bC�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾u1�<��?7�-?��>Ŏr�1�ɿc���y¤<���?0�@�yA?7�(����V=ź�>K�	?
�?>�41��F�����Q�>�9�?���?�zM=��W���
��te?Y�<<�F�X(߻��=�2�=�=D��#�J>�V�>z��yA��Pܽ�4>�˅>��"����cf^�e!�<�q]>�ս�B��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=u6�����{���&V�}��=[��>c�>,������O��I��U��=���;�ĿA�"�����=X�):��s�9��>ܽ`�������ly�8񽞕h=A\�=?�g>@��>��b>�h>A6[?g�n?�>]� >�
��u��Nؾ��;�ʃ�z��&D���J&� 3��|��h�꾰�����j�����"=�%=�=�#R�_���n� ��b��F�/�.?^$>��ʾn�M��[+<TQʾ���� Ƅ�ݦ��T̾��1��n��ȟ?$�A?����w�V�%�����?���s�W?�I����Ѭ��w�=�2��x�=�B�>䁣=���K:3���S��C0?^�?����[����'>�a��E=�,?�D?.�<��>o�%?�l*�*���eY>�E0>�V�>�5�>W~
>����G۽=?�S?���U���>^�>�����I|��\=�>��6��Q���v[>��<����`V��F��<!H?�f�>fD�]D:���ľ1G��ZA����?��?��?3~b?�7�??禽H�*�t2e�O��%T>��V?��q?V�>h�[ľ��Ҿ��?2�7?uU>v���6����a�����)�>��]?kl)?0�L��q����|׾¡?@�d?$�F��Z���%�샬����<�D�>m=*?����?�E?��=D/��DԾ�.'C��d�?��?2��?X��=�ѓ�
�=-� ?�?ƥ�O�������wؾP0�Q�>U�վ�z~�y�.���e�|�,?��?["?*�J�Id����=����u��?�Ƅ?�c־�|�=� ��*\�`���!���,�=35������6߾ۉ5���徒���b��OZ���>f�@alt�O.�>�A���ῠ����Vu��找����*?2¯>y5,��6��g�y���y��E���I��ܖ���>R��=��ҍ�%{�d�I�,`��?�3Z�Oգ>*�b�Ѩ��b�����ǽ$�>b�>-ĩ>w�ļ9曾��?b�=v˿����	�Q?���?��?��)?��>&�-��07<o[8?��\?�E?p%�t�0�A&�y�i?�����b�r�6��E���@>�/0?�q�>_*��۪=ŧ >���>�Q>81��ĿW �����u¦?���?��F��>Y��?�U+?ʕ�`]�������)������v=?�*2>m¾��!��f;��Б�
�?ܛ0?�H���]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?v�>K��?���='��>,C�=�﮾'�M��%>��=��I��?S�L?ϓ�>i��=	v8�"�0��F��.R�,���AC���>%�`?��J?c�^>����d�&�����q޽��2���n~C���>�6�ݽi8>m�8>>��H��SҾ�?F���ؿ�����8��g%?Yrx>��?������6��}R<<�e? 5n>�F�H���r��jͽ_�?���?�O?�BѾ����>��>�as>����o��g���=�>í@?x�����ci����>�<�?l	@Nr�?�?g��?1[��g����ey�� ��n��w�Z=Y�N?G���{�>YA�>ּ:>sQ��"��� �u�fu�>Z3�?�K�?r.�>}gN?�KX�s����O.>�I>X?vF�>�E
�a��7d>L�>�x$�ȱ��!��r^?ɬ@��@��X?������ѿ:���Yz�������>6��=e�9>�!�eO�=�%�=��<^�-����=CG�>>�>K�r>��H>��">�O,>����Y�(�憎�n��xB0�z�����J�����T>U��
��滾ٹ־�]��?�����c��t.��U"�A%0���Y>-�D?BcW?:�?��1?�u@>�/?7AO�}~8��nr���㾙"��"�>�!@?�#?s�>Fh���j��Y��x����Ҿ���>B�>��>��>e�>����U%o�KVH=��x>�#>�-c=��ݽ�O���+>�C>)�>b�?:n<>��>ȴ��7����h�m�v�r̽���?C����J��2��C`��������=l.?.�>���_Aп? ��> H?�ؔ��%��,��d>	�0?�fW?ro>�ⰾE�S���>���j�j�ט>�
 ���k��r)�"CQ>5S?�wi>!fz>N�2���6��sN�n����7�>��4?�մ���;�zv�яH��3ݾX&Q>p��>�.�VD��Ԗ�f6���rj�~o=�L;?H?.�������>�q��9���S>�_>i�=��=+�L>�dg��
ǽ�L��(D=�^�=@�`>�#?;Z*>��=���>�"��k[T��I�>|�J>�+>��@?�$?�� ���c����1�5xn>d�>Y��>��>~"J��z�=��>�F`>��g���w�!<@�dR>9A����[�T���4c=�$���P�=���=\���(=���=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾUh�>^x��Z�������u��#=(��>9H?dV��)�O�>�w
?�?_�ީ����ȿ|v����>P�?���?M�m��A���@�|��>%��?�gY?`oi>�g۾`Z����>Ż@?�R?�>�9���'�o�?�޶?ǯ�?��O>��?�o?	d�>���;B0����\Ї���=S�4���>�>޵�[�F�rl��0y���7l�[0��>i>np)=3Թ>������Tt�=H��턣���a�3�>�d>��B>S[�>�S?I��>�[�>i��<�!��9�{������E?ȗ?�M"�h
���*�>���=F:��@�W>R��>����/!@�v�4;��(?�u?V�o?�|�>��1��X��x�ۿ�ќ�xF����L>�?b��>�Pk���>^���/����j~>���=˲|=������&�<�q�>dL+?��?ѭ�=8T?.�E?�5z>Vܠ>��V�����-c����>H�;?/�>!�?N��>L�ܾ�n-��k�������wW�X�Z>I�X?<
?ٟ?���%㋿ӂ�>�_�G(���ҁ?�$w?>���9��>n.�?4o~?���>ޠ >�q���s!�pʾ���>��!?���D�A�
c&���<i?4;?6��>ʤ��h>׽Q�ݼ�������?�-\?&?���iJa�T�þ&u�<MW�s.S���;5y:���>}�>%"��Z´=�B>�=��m���6�޷i< ��=��>��=�6�oގ�$?dW��B��w?�=O.���P�5�=�r1>Y�%{?�;g�P��շ��3���*���S�?�~�?Te�?Iٽ�c��a?�4�?>=?���>V�<ꪹ�I���]�Y��E��}��<��>�4>�ͭ��������� B�gdI���w��>qe�>��?��>`�d>w��>�Ö��+����#���5d�}�g|6�^�,��������R�
�Ɏ���҆�S�>�[|�m��>��?��E>͸j>4�>l���>��(>�w>w?�>x\>�8>�=�=TZ<����O?7��bC"���ྰǴ��J@?�4^?�1�>�G��5���=�&0?�.�?�^�?!p>��n�$�.�R ?�z�>8nw�s
? �=1�>�K�?<cH��~e������RQ�S܂>�TǽD�9�l�O�/7o��Y
?ƒ?��6F־| �f���*=;��?�f0?g�U�:8���h���D�"5���<crνt�(5�x:Y�����V��;	f���2˼�\.?
��?������3Ͼ�T���P���>��
?A��>A?Զ�>�1� ���A��>�7�I��[1�>)#s?׾�>�*J?�U:?Q?C�L?Ӣ�> �>����;X�>��;���>�>6?�`.?�1?�"?�H'?,�M>?���@��`eپ��??�"?<i?���>�g���Ž�W#�
ʣ���p�Q��Hq=��;t>콗I���+=�M_>��?>���m(���0>�j2?]^�>��>�	��6����=Yc�>ؖ?r8�>C��������o6�>�k�?��$���/=x%>���=ޗ��'�����=�r������6n�q�;�'=���<DxJ=��C<���;]y��6�����Qp�>?Y*>c�R>6ڞ���D��Y�>Q�Q>8q�>�4>G�w��
��$ ��� _�'�>73�?ֹ�?H>�E>��=�ꩾwx�E� �������=�?Fm.?�'g?��?loT?��(?%@>>���=������d����?k!,?���>G����ʾP�o�3��?�Z?<a�����;)�R�¾��Խ�> [/��.~����XD�.G�����������?�?�A���6��x�ȿ���[��b�C?,!�>�W�>��>#�)�b�g��%�h2;>��>[R?c!�>'�O?�5{?�[?T-T>�8��(��ƙ��B5�q�!>�@?���?�?�y?h�>�F>+�)��%ྊ1��$2���*؂�l>V=��Y>���>�.�>��>$��=�$ȽEP���?���=Z�b>���>6��>���>;5w>'$�<��G?K��>@��/��[-��Hq���
>�e�u?���?�+?�`=V��(F�=���A��>h;�?��? S*?)hR��K�=��ռ�����\q��Ƿ>kj�>ꠘ>K�=e1F=��>q�>�*�>;{�j0��Z8���I�I�?��E?-h�=�ſf r��a�d_��zM<妎���j�i~�� b��h�=uÙ�5n!�#����\�8Ơ�&���Գ��i��**{��K�>��~=	��=��=�Q�<�������<�4==X@�<�=?�x�p<1>���o�p���>�s�Ԑ\<�K=:(>��ɾ��|?J?0,?��D?w,~>f>AP]���>�o���?
T>r1M����T�8��⧾�x��B�ھ�xپ��d��:��X>�H��*>�j5>"��=2<�<3&�=}�N=��=�5G�}M=���=���=�Ϊ=�n�=�>:>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>K�8>o1>�kS�%>2�rV^�Fmf��Z���"?�o:�&�Ⱦ��>�J�=/ྮ�Ǿ� =}�4>�Nl=���U�Z�r�=}y��4=��m=���>��A>��=���C�=�_@=���=QwM>�Z���,5���/��<=�G�=;c>*$>9��>D�?�a0?�Xd?�6�>�n��Ͼ�?���H�>��=zE�>�߅=YrB>'��>>�7?q�D?�K?��>��=	�>��>p�,���m�m�̧���<���?lΆ?�Ѹ>-�Q<%�A����~g>��/Ž&w?�R1?�k?��>������9?��AD��FS>�:�=�}�/U��c�P���}�jv%>�*��`{2>��>>� �>@�>��=;J>��>4�:>�M�=�=~=���8Ro�k�.=8��=oV�=
�*p����>��<��>>8ö<����:w�<�c2<�ʸ=��>�͏>M�>$�����=÷���M��A>�j��3�3�d�d�mqz��/��3?�ƽa>K�>]`;�I��+��>�>C"h>��?[�?�S�=�꽾�¾i袿�-�����]�+>��m> 	)��[N���y���T�6㹾/��>���>�ͣ>[�m>x0,�ٙ>� �p=V
ᾟc5���>����% �\��3�p�m�������i��	��_D?5����F�=��}?�PI?:��?�Z�>�F���ؾT�->EP���=�_�=Ur�v���� ?��&?_��>E����D�uྦ��Z>D��H�5ڝ��3��C=^ܾz��>rs޾��þ�MR�^���T�|�K�rc��QM�>�	Z?��?M��9����p@��:�t���8��>���?˰�>��]?P8 ?Uq>�����n���A.?J��?���?��=o�=?A����>[%?F�?l��?AĈ?&韾���>>H߽{d$>���@�m>�n�>�>>!uA>T��>	G�>m�>����[S�P�����;�S�h��=�>%vB>�3�>ng�>�(�=%�>C��>1�>W�>��{>_k�>�z?:!�>�������CT?�I>��>Ӓ0?gf><�D=�D��R�;�r��I���nf��[���#�#|�Y��<$Q#>X���2�>�ÿ��?.�k>��ʾ�9?����2n�=�RF=�!�r�1>}�F>Z��>D�>"��>��=a�>�F�=TFӾ�>����d!�-C�+�R���Ѿ�}z>Z���h	&�����x��KBI�_n���g��j�9.��<=�,̽<H�?����k��)�%����?\�>�6?Lڌ�y��İ>���>�Ǎ>yJ��_���Uȍ�h�j�?��? 'Z>��>-W`?�v?m]>�y��i�\���q���D�iec��_�al���Ā�N�	�Nʽ�Z?F$v?V�C?Eq<� t>�Vy?ߴ$��Ջ�l��>�[(��x<�[
=2I�>���>ie��fپ�¾�G�TbF>�l?a��?/?��a�+�0��?>�8?�8?q�x?�8?��F?4�?�X�?�$>���>� ? w0?��/?6�?��Q>]��=D(,�KC>=�l����� ���2����Y���Q=���=�ɧ<�
f<�=��g=z��#S<)J�<e�#��uv�@4�=&c�=�>���>7�]?�K�>ۜ�>��7?Z�� u8��Ǯ�+/?��9=�������~ɢ�����>L�j?���?�`Z?vSd>��A��C��$>]�>�n&>�\>�b�>���q�E�)��=zG>R>ѥ=�gM�Nҁ���	�ᅑ�ó�<T->P:�>���>0����+>M͟�ܽw��}h>-&U�����&T�Z�H��|2�Qpv���>j�L?X`?�=-��l��W�e��i'?�u=?�]N?\�}?���=�e۾��:�ŜI�����K�>��<������z���;�p��;:m>iH��Hߠ��Zb>����q޾�n��
J�z��$M=t~�%EV=:��վ3�I��=�
>����9� �����Ԫ��/J?��j=�t��DWU��m��u�>پ�>��>�:���v���@�����?�=A��>"�:>�������|G�X5����>XC>?|�X?��?�JP�1fT�'�:�F2�j�����Ƚo�?��>��?8cT>�z�=c������_�6�5��;�>�W�>��j)C������.�\�%����>o�?BR(>W�?`�\?�C?~�c?ܘ0?��?��>�:�����]3&?iX�?뛃=�ս��R��O8�GF��^�>-)?	�C��ڗ>u+?�>?9'?��Q?a�?y>�� ��?��>�ߊ>��W��+��:�_>��I?�²>��X?���?��>>�5��q�������)�=.c >k�2?�Z#?��?$�>�5�>�r��1C=W#�>�e?��?��b?�:�=�/?�u>,��>�� >���>B��>�?�P?7�o?�mC?��>I�<���������X���:/�
���;Cm=G��q�	��N�o�<袼3�5��r���/ڼ����(;�R;�\�>��s>
���0>��ľ@#��O�@>�N��DO����di:�%��=���>�?[˕>�#��ƒ=ύ�>)M�>����"(?��?�?[`&;7�b��۾�K�l=�>�B?��="�l�π��m�u�J	i=��m?ҍ^?|HW���j__?j�q?fn�\�6���i�w���w9�f�f?h^�>�*Ҿ~�>9�?xZv?�-?4�r��+��A~���N��c�5=���>�S!�Ǣ�����>(�5?�p ?֋!��FF>�FŽ�[��v%��a?0?h��?�i�?�>�S��,�� ���?����]?]y�>\�� �"?\��b�Ͼx*��F��:(�!"���!���J��͡���%��烾��ֽR��=E�?"�r?�Hq?��_?�� �1�c��^�^���hV�`��(���E��
E��C�K�n�^[������|G=�H�T8d��<�?OH6?�x��;W?�}�rH��bA��~1u>�����=�Ψ��4�>�+R>«��P_=�,����0?� ?��d>p?e?v����3k�`�q���'��ZCa>���>�st>|>v�i=�\9�"6B<��ؾѣ�<�
���v>d/c?�vK?�n?� ���/�5@��%� ��D�n䩾b�A>��>��>�HX�����&�O�>���r�ī�Tԏ�}s	�+�{=D2?���>.��>�З?We?&	�6ر�mCy�0�p�p<nh�>��h?Ǡ�>��>c̽%�����>]�l?��?���>��ݾ&�,�P������>�8?՚�>^�!?��	=Z�<��w��9��l����D�r��=�Q?S|�\�@�Lm�>+4?p��=�h�>���>۳��l��^5�u����鬽��?��K>E=�<+�����3P����/(?2z?�����w��s�>��#?���>�Mq>�Uv?;6�>ȑ��b>HR,?dm?�`Z?�I?���>D/<�w6���׽JȽ�1���>t��>���<�q=�"�'%��ù;�"�=lu~=^��Xg��NA=Y��<2�S=X=�!�=@�ܿ66��cžZh0�̚����B����KA�YJ�����.b��������]�>��v=�O6��l8��j���	����?
n�?�l�#
��o��e䉿 ��h��>�ʞ=�}��j.������i��i�َ�GE.�ٜS��e[������'?湑���ǿ߰��<ܾ�  ?SA ?��y?���"�[�8�ʭ >;9�<v.��z�뾲�����ο��� �^?���>��(/��F��>���>u�X>�Iq>n��V螾�1�<��?�-?
��>�r�:�ɿ`���
��<���?	�@��@?�%�V���_=9��>:�
?:�C>�3<��/�Cb��<��>���?F�?�\=�T�V0���b?$Ɣ�3�I�J,����=�v�=��=ӆ
��KI>{��>��$�ثF���ؽ�p7>B��>f`�T��)�b�v��<�Q>Q�ٽ��m�5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=A��ƿ�W �N "�x�=Sʍ<��?d.��\��*�/�e���uF�� V�M�=N/>*4L>�&�>]P[>ߦD>o�`?QW{?u־>�� >I'K�{L��"{ݾ�W�<j�s�@�U�!����78�"1��̃��*��?������0�$��!=�e�=�6R������� �2�b���F�d�.?�$>^�ʾA�M�K�-<ruʾ����_.��j好2+̾�1��n��̟?��A?�����V�7 ��e�a|��v�W?2>���笾��=���Xw=��>�w�=����3��xS��p0?8M?50��W����+> � ��s=��+?��?E\f<���>̣%?�(��E⽾9\>�4>Ř�>��>�	>�����=ٽ�=?);T??^ �漜�?Z�>1ٽ�V�z�ձd=љ>�5�<張�Z>�:�<8�����Q����<�<�Q?!��>�'�X��>G��u��}w� �?�
#?D9�>~�u?ޅ6?OY����WS�(��n�3=��V?Z�Y?���=���</鯾�P����2?~X?�B;>�?�kȾ��&�&���?oDe?k�>���\�s�n���6���WD?&zT?SI�\C��|��5Z��9#>��^?��?���Rx>z:I?(	 �����ƿ�F�'x�?���?���?��x<�~)��S>)K?_��>m$V�v�-�y�>8/�܆T���>a4 ��?����׾���E?uM?� .?!�0�" �ʹ�=W͖����?���?������i<?���j�����j(�<iS�=��/�Z�)���)W6���þr�	�����ȼ$��>�N@�����>'�:����ο����XϾ�Im�8c?R��>x�н�Ǣ���k�fu�$uF���G�pq����>�w�=U`?������|����C�\#)�T��>ZR�=Z-�>�,�Dђ���ྮ?@�"�#>���>8N�>�]��B���]�?p��C̿P^��n��Q?�;�?r��?�?d��V���������5�>?��J?�tw?7��8u����#�j?�_��|U`��4�uHE��U>�"3?�B�>N�-�p�|=�>���>�f>�#/�y�Ŀ�ٶ�2���Z��?��?�o���>q��?rs+?�i�8���[����*���+��<A?�2>���A�!�E0=�HҒ�¼
?V~0?{�e.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?츸>ˊ�?���=b`�>�>���@<��=WT�=�����?JK?#�>�C�=)&��)�:UD� W������A���>�%b?�:J?�zg>����j��B#�1 �yj/�#'��0��� ��X���>�>>�^�=L�g!����?�y���ؿ�k��'�'��4?lÃ>�?���[t�8��PH_?�+�>�5��3�������f��?Y<�?b�?��׾0�̼I�>D�>�R�>@�ӽ�H��蘇�FN7>:�B?���.��Z�o�V�>���?��@�Ю?��h�6&?]�&���<��&S	�,"n�GL>e�D?�н��>2?�0>ށ�e���%��P��>�=�?̹�?5��>;�a?!_���6�N�e<���>�f?O ? _=U����}=�[?FN�$�s�j��/�c?�b@�@�]?.✿ɀ7������gؾ���=;�=bq�>�*.��,=�2=&h�=ێ����)=(?�>b!�>�B�>�Kn>�1�=z��=ޤ���#�P����N���i:�Ō���"�!�G�����[��l��ݽþ$ӾAɽ�k�Y�`�^'U��nI�lZ���L>�`>?5�1?�<a?_�>?�/�>K>ι?��6�u*�B�<�&�>�3?-�?i	?�i�=o��I9��Iu�VI��W��m��>��(>�kq>G*�>eTT>�>4��=�"<y��G��=�(>� �����4׃=G+G>���>�2?�C<>��>Fϴ��1��j�h��
w�n̽1�?����S�J��1���9��Ӧ���h�=Hb.?|>���?пf����2H?%���z)��+���>}�0?�cW?�>!��r�T�3:>:����j�4`>�+ �|l���)��%Q>vl?��f>Z<u>��3�W8��P��^��Ĉ|>86?�����a9��u�T�H��TݾAYM>Ǿ>Q�C��g�G���E!�$i��X{=�x:?k�?�ݲ�)հ���u�PU��
�Q>;%\>B�=x��=�^M>�d�yǽ��G��C-=�u�=��^>h?=.>�Y�=m7�>�����S�:��>��F>�2>~�@?T�%?�0��:���v��'{/�9�u>"��>�a�>��>S�I�³�=2<�>/�a>Q���H���ǰ��G>�V>�����U`���j�N~=B���*�=���=`��f�A��/8=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�b�>���U[��/����u��L#=��>C7H?�@��}UO���=��w
?�?]�r�����ȿ�sv�/��>b�?��?��m�(@���@�/��>��?�iY?`�i>
f۾�kZ�i��>Ӿ@?>R?��>>�%g'��?{ܶ?̬�?�L>5��?��r?���>Υ�� �)�x4�������H!=�$���H�>��=붾GD�Qg�������l����@r>��/=M'�>�b�Nݶ�o��=���NW���F6�_�>SR>�nG>�I�>���>���>���>�"�<p���r�v�%z��r@??���?���ұs����>v�>I��=M�}=s�>��޽�(���>^??Pl�? �g?�G>p~ �����Vz޿�I������Sm>q;?[��>��=��>Iw��F����/>	��>�W��e�9�������'o�>�8?�F3>"Ā��F ?*+?6|>ys�>�3�1����5�u[?E~>�d�>�Oh?m��>Pf��ҩ��!���0���>m�w3>d�~?�5?Ѡ�>���\���Wg�=Yy����=��?�/f?�!5��*?&��?�$?wVP?+�>����۾"����->��!?� ��@�i#�|���
?�?�Q�>Ǫ���o ��R��k����?�\?`�$?�g��1c�fԾ`��<6E���5;1�p<�Pc��%>��>fw��㸂=y>���=��e�ݦ5�|ʳ���=�\�>���=k!<��-����?b8��'�jtK>�_h���9�^�
?;�J=Xk��m*w?&�Ǿ-}� P��~≿��V�EY�?+�?�g�?]:=�!k�!�?]w�?۸?��?������'���a\�
�b��jV�̏�=㲩>��>��m������������zG6=�:?�]��>�>�'?���>^]->��>Hs����(��߾�Y��c�=���*��.����C뢾F�C�^=J���3����E�>�2`����>�(?��>�ז>h��>T[ŽU��>s�>;W�>�3u>�m>���={>o��<�=��5R?�ɿ��'��d�����%B?�Ad?���>��j�,x��.����?
��?���?/#x>h��C+���?���>���<S
?R!7=�� �uߏ<�+�����*)��� 
�a,�>�ֽ��9�M�e�`�
?�x?�م��̾�C۽n"��{|q=���?G�(?Y=*�M�Q���o��vW��?R�Q���<h��_���$�Xp�\���|t�����@](�R�4=�P*?���?�N��쾔߫���j��}>�FCf>�P�>kؕ>���>��H>�p	�Z�1�u^��J'�����[��>n�z?WB�>�I?�:?ێO?�SM?�c�>0D�>3������>�r�;|,�>���>4�9?�-.?��0?1?j�*?�]>�] ��i��?4׾�i?,/?Q?�?e�?Y���^%ƽ8U��L�H���w�j"}��Ov=mJ�<bqӽW
z��nR=@U>�?����5��9��<i> �7?=N�>xo�>����p�����<���>��?j܎>�����s��H� �>���?4����=�$>�B�=�E�D���4��=壖��ˍ=? ѼJ�7�`PE<�}�=�l�=��9��=���N:+�
<`е<Wy?�?�=`>�
�>V_߾i "�ӄ�~�>j��>M �>ޮ�>����wu��w���hM�I�>���?�8�?�^��[�=8�>c[����ݜ��`�뾦��`�?}I?2
K?$Ԗ?��U?�?�]	�I�)��
���x��b�Ծ�?�,?��>�����ʾxۨ�q3���?�/?b:a�y���)��r¾�Խ޳>M/��~�J����"D�������Ƚ��ב�?��?�?���6�Uv�廘�ۀ��߂C?��>�U�>��>��)�_�g�n�+�:>�a�>:R?OQ�>�L?�u?j�W?�6e>��/�8��(���ͧ��u>��=?�ڃ?�R�?Nx?c;�>=�&>�$����	�������������R@=��S>�<�>��>��>���=�s��ԡ�6��w~=�Tn>��>�>���>��>,=??���>���$��	�ľ2�����{?�h�?��8?���=��P_�(+��kCH>@-�?��?O�6?���>O�Z���������u�>ᨷ>K�>��3>�-<j��<��>]�>yp�����5�n��=�M�>B/D?��}=����/tb�*�v���U��7f�؀��B(���н�H �z��=r����V:��W������s�ؾB��󻾁G���� ��>><�T��=�Z>�_>��[��}�<V,+=��y<=�=���`�*p��ڛ�a�Q�Yc�;�0�=h�=���������t?$*G?�.?��H?�@�>S�>՝ٽ��A>e���o?_܁>���<'����K��N������' �ʮؾ��e������>�JF�7C>�4>CR�=*؏=�L�=R��<�4�<S�w���$=���=A��=��8={��=4�F>3>w?�{������v�P�'��[[:?��>�R�=J�ƾ9@?:�>>�1��L������8�~?���?�z�?^'?��h���>0����z��ꊓ=5D��z	1>}��=�G4�3�>��L>��O���a���C�?�h@l??���_�Ͽ2�0>�8>W�>��R��H1�$[�0da��xY��!?�T;�]u̾f�>�=x�޾>�ž�O2=�6>�b=س���\���=yU{��j==?Jm=�>��C>M��=@������=o�H=c
�=��O>G���{<�>`-� �4=��=� b>K�&>Ͱ�>��	?�B)?��^?�f�>?4B��\Ҿ/̶�oPz>7+�=��>��=�sv>3��>�;?�&E?�fE?��>�O�=�D�>ƞ�>!9�j���ھq�ɾ�C�H+�?ш?2��>�d�=Պ ����6�+��誽
�?��4?�p	?@��>&(�$
�#��f?��!���=���=ʌ�����V�<�ѽE���=cq�>���>j�>M�>Ƿ�=6�>���>��>��<x>�=�I����<=%2�j��<�oѽ���;𘟽�U4��秼���<�^�<V����^Ղ=sv�;飞=b��>l�>x�>e{�=���	�g>M鹾�H�;�h>��EO��Pi��U����Jl��S�>�s>f9�<˔�v1�>H�>�=v��?~�t?�y�-e���m�����f���y�Z\>�>9J�sZR�w�v�̒U���پ�>�k�>�p�>��h>�p2��%E��-=!ྋ1!���>�o���5S�/�"�yn�jV������DBf�E]��:L?箂��=�2r?'CS?�R�?���>��|��kʾ���=pj�%E뼭=�<�=�*��Ҡ?z ?���>���6B�X�վ��#����=�LL>s�M�V?��;)#�=W����ܼA	?���B��M9S�>��Y��IX��G��(�>��C?�K�?�8���q��x�G��!1�*�_��q�>I&j?=\�>V�5??*>Z�T�"�$�v�=F�m?�?�[�?2y=N�>�[�����>��?�ۖ?@�?��X?E�U���j> �;��=l��=�G�>��>>:�>�S�=>��>���>�:?��Ґ���i�������|�}-���.y����>� �>�0�>�^o>��\>�C>:�>��>;ʴ>
l�>��>��>�����)��Z?*��<�/�>��A?~�}=.�c=��=�7�=F���X�־�e�N5�|�F;�6=�h�=�@>�M�;�<�>t¿��?�a*>�D0���<?�]"��H%>
��>z%>��G=%%�>�^�>�v�=hb�>j�>o7>,;�>�&7<�����H>���3��K_���W�f]���!>e��#�2���ᾀ�콍ޅ��8��Z���m���u�  +��)>́�?�J����Q�+��bv5��%�>�W�>�� ?�h �qf�_�<iW�>��>�n	��ߢ�N���3���c�w?*t�?R�p>���>4c?�A-?w���ҹ8�|xU�4�a�P1�6J��	]�Ɣ���}�Py��F9���b?FGp?��I?X�K;�Z�>��?m�E��>��W�g>�M�Z%����=6H�>'����Aa���ھt�ӾP��\dO=x�R?2�?�?��Y��G�=Yx>a�
?��?�؄?�P>?,��>]1D�K^?�Ɋ;�;�>��6?dDN?v"D?�d&?g��>G>5�}��p�=�����%S�b|�e$ƽO�h=ŝ=��<���<�Ȣ=a�&>2��<�XO��Ӂ�
��<'K#�#=��=i>T-S=o¦>�]?U?�>���>'�7?h��ps8��ˮ��$/?Z�9=����m��.������O>�j?���?+XZ?8>d>��A���B�c>�Y�>?&>P
\>�Z�>Y�ｻ�E�6 �=�V>4Y>�Х=��M�́��	�ҋ��`��<�*>P��>��>�3��}�*>g>��z�g�C�n>Dh�'5ľ��]��0A�v�-��tp�mA�>�QK?��?㢉=������d��&?1S=?K�K?�~?���=N2޾*�;���L����5�>��<�/�?���Ő����6�컼<�f>���ݠ��Xb>���r޾v�n�J�s�羖LM=~��EV=����վ82����= 
>&���� �����ժ�71J?ˤj=�y��3bU�0n��U�>���>v�>�:�$�v�C�@�����x2�=���>R ;>�e��� �*~G��8�:݈>�GE?�R_?�;�?����"pn��mC�W5�������*�T�?���>�	?�~=>�=��������d�D�C��>Fq�>(h��&G��'�������#��|�>];?��>S?�hS?T ?Aa?��*?�(?F�>:J��ƻ� B&?6��?��=��Խ��T� 9�FF����>w�)?+�B�ӹ�>M�?�?�&?�Q?�?Z�>�� ��C@����>�Y�>��W��b��J�_>��J?ؚ�>h=Y?�ԃ?��=>_�5��颾�֩��U�=�>��2?6#?D�?㯸>�+�>�ܛ�����2Xp>c�?��?X6c?K`G�w�?iQ>�"�>v�{>V�?g�? ?�s?Y�?�s�>���>�";/��Q5�܂"�����oz��T>��b<�X��-=�]�=M%>�ο���}��`�;�Ô���B=-=��0q�>n�s>/����0>�ž�����@>�����N��	u��}�9�ȷ=aF�>��?�)�>��#��=�μ>H^�>,��b(?d�??��
;%�b���ھB@L�1<�>B?i"�=��l� ���u���j=zn?f�^?�V��@����i?��o?��8S�b���)���t�E�k?�{>�y�7=�>c�_?��n?r?ic��ۈp�u����AX�务�2�v=�N�>��/�����J$?�2?�p�>"!	<1�k>�z^��J���|���?~��?�ݳ?�Ҕ?l5�=�]��oI�k��KM��Z8^?�6�> B��K#?<��^�Ͼ�`��^Ԏ����m���#���Y���1���i$�o�����ս�X�=�?�	s?_q?&�_?9� �v�c�-^�I���FV�y]����i�E�"#E��sC��sn�Y����������F=4J~���A��ѵ?�L'?}0��e�>������G;�IC>�U��!Q��R�=b���?=��X=<�f�z,�P��_�?�a�>���> z<?�[�K-=�l^1�r7�����+x0>���>�	�>���>�2�:b,�j����Ⱦ"䄾�׽h�v>�tc?s�K?��n?���+{0��k���^!��F5�����aB>�	>D6�>�qW�3��~n&�e>>���r�r���T����	��-}=�2?dv�>F\�>�?K?֧	����� w��W1�J��<�{�>��h?���>�:�>HbϽ�� ��!�>�jh?M�?�t�>� �M8��̈́c��/���d?�ߨ>�'?7��=":̼�pV�֓���儿:.�y|�=��|?ڼ��X����>��M?�W˽���>��W>6�Ž����+E���ȾN�q�X�'?�'T>�g<��!���ܖ���#���(?��?�����*�b�>j�"?^��>���>w�?y�>þ�I|;l?FH_?��I?KxB?(��>�=�,��
3Ƚ��$��,#=Q��>�!X>�_=Y7�={��61Z�Y��ӧF=���=C	ļ�.��F6<P!���><��=�z3>��Ϳ
v@����� ��F	�����*�j�"���S�5%̽R���A���S3p�z�����<���uP,�1�z�l���o�?���?�죾�����.������s�#��}�>9�	�?��� ;R�	l�O྾^#�F@��	5�W�!�����'?g�����ǿ|����Aܾ� ?Z< ?�y?-�=�"��8�� >��<�g��E��Z�����ο|�����^?���>C	�m;�����>A��>��X>�;q>����~�<��?�-?l��>זr�J�ɿ����Bܣ<���?P�@w|A?
�(�4�� V=���>=�	?��?>�W1��H����)O�>�;�??��?^�M=��W�T�	��|e?�<��F�Э޻f�=�\�=I�=2���J>�W�>��X_A��(ܽ�4>kׅ>Vn"����
y^�!i�<��]>��ս�;��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=2� �q�Ŀ�$����V�<'�;*`мQ��{�����YW��%K`��p����W=���=x�Q>�>�J>�4a>�\?n�t?�l�>I�>��&�>\���vѾ9�޻�r�g/�Ú~�+A1��ϴ�����پ2p����`[�8"��� =�w�=.7R������ ���b���F�7�.?�w$>��ʾH�M�e�-<�qʾn���� ⥽�,̾��1�Kn��͟?��A?������V�����w�󓹽��W?�N����U笾C��=�ޱ�֘=�>�~�=����3�d|S�b�0?�y?fܿ����@�>oG	����<4,?}?��=IS�>�(?|�0�{ � �U>D�3>��>π�>��>İ��~�׽��?T?� �:����l�>�Ⱦ��}��̏=�c�=�0��t���_>!e�;��������|����=�gH?�֛>b#:�Q���ƾ4W����>Ǆ?��?�E�>a|�?�:?�J���#���~�k$�Г����\?�wt?uJ>����L���c����?�)U?ƞ�>9�$[��
+�C�����?m�n?���>p.���}���a����� ??�s?*V�T֕��>����o#Q>��>e��>Q"�	2�>�8?���ו�uĽ�U�0���?I5@���?r�=aK��)�)=Qx?���>��=��h�����ӝҾ���=��>�`�"�Z����A�����Z?)�?~�?�!�K���D��=�Օ��Z�?;�?����P�g<2��.l��q����< ҫ=�3��("�/���7���ƾܼ
�ݫ��Ƭ��D��>6Y@�g�(�>�98��5��RϿ����\оiXq���?��>ΨȽX�����j�Ou��G�"�H������N�>��>����M�����{��p;�1Y����>`+�4�>ݸS��'������I�5<�>\��>)��>})���佾�ę?5`��*@οJ�����&�X?.g�?�n�?Op?��9<��v�#�{�Y���.G?Չs?�Z?��%��:]���7��ha?�y�� ~`�\.�T�_n���?�+?M}-�H[>�~�>�!�>�q���a��ٿ�Ƕ��?���?L=�?����>�ݓ?��#?�������?�2���F�9�>|z?���=*Hƾ��.����ݳ��44?��c?ljQ=bY*�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?I6�>H�?@�=�c�>�T�=g�;�"�&�">�=�2@��j?��M?q�>)�=��8�3�.��BF��jR�>e�p�C����>Db?A�L?�a>F����80��@!�6oϽ��0��⼮@��+��۽�`5>SR=>�>>BD�z�Ҿ��?>���տRz��`)O�,�?Cd{>�?��(4��:8_=�]?��w>��ke��z���%��?���?M�?$�޾ʛ�;��>nq�>��h>�l=�KS���M��ߓr>��=?Y{�-���\�a�~�>V�?@��?��e�b�?���;�����m��?�Z����`>:t<?L־��>�}	?֙�=|�y��ˣ��i}�GW�>�.�?���?��>BY?]�f�a��K�=��~>D�c?���>£ֽ�e���	p>=��>m��
�����C9�?\�@�@]�q?�����ϿB_��.������b�=���=	=1>�[����=��=��%t���=}�>(�i>b[}>��J>�R<>(�<>�G���*�8���P���0TH��B�?������Ż�	�=��J��	���
˾n���n���u��J�*���Rˊ�qL5>i'W?,zW?�Q�?}�N?��>��>�^��_������d���>�};? *�?h�?'��<�˾���]�������䶾��>�m�>7G>�>R
�>�3��O��=��>��>�=��z��o�>���4<�Ӹ<M�K>i:�>y��>�C<>�>Dϴ��1��K�h��
w��̽+�?����X�J��1���9�������i�=Wb.?�{>���?пk����2H?����l)�6�+��>��0?�cW?��>���z�T��9>i��Ŧj�>`>�+ �l���)��$Q>Il?��f>�u>��3��d8���P�u|���k|>�26?�趾�F9���u���H��`ݾMM>lľ>��C��k�������exi�φ{=(y:?��?�6��ⰾy�u��F��JR>�;\>�c=Ui�=�XM>�<c���ƽH��f.=���=ڮ^>E�?R�(>8a�=��>+�����V��Ѩ>z�D>8:0>͎B?��#?u�����z膾J�,� �u>�`�>O��>e<>��M���=���>�jc>���o��z�d7E��W>7�~�m�d�k��"l=��!2>�}�=�3��~\5�f'(=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ��>�[�����������x��7���>�Z?���ev��#����	?��>��������uο,0|��G�>2��?�:�?�Ng��7���:��K�>q\�? �\?�)�>��㾍zt���>�>?��N?1�>}B�?�G�w�?�X�?Ss?KGR>�?�?.3u?��>B��� ��������Y�<Du0�>���=���O1E�h哿]׋�cVh�h���u>��9=��>3�
�>���S��=�첽�:���m��8�>��N>�W>�`�>o4�>���>0��>
��<{hƽ��u�e��ˑK?�?x�+�����rŬ>�`�=l7r�9m�>cd?֌J�n ��7�>��O?wo�?�&M?��>�E ��>��+�ӿúؾ+��䍜>��0?�>��\����>f��+��ގ�>��g>J�>�i���!��HK�ed�>�E?K`w>�6=V�?�#?..>Co�>"�J��1}���L���?nF6>ؗ�>5�|?���>�����\ ����"쫿��m���:>{�y?m�'?ό>+}��{ޓ�iv#>H��a߼aE�?
0?�.[?k��?X�?�}@?�$�>+*J����;��ڄ�=h�!?��ͺA��M&����~?�P?���>
4��>�ս�Nּ���}��3 ?�(\?�A&?ܛ��+a�N�¾�3�<��"�(V�U��;�uD�u�>��>���$��=
>:ٰ=fNm�aF6���f<j�=��>��=�-7��w��ܰ#?V�Ͻ�#g;���=2x��'K��3>��Q>�~�W,�?�J־BU8��Q��o��������+}? j�?87�?3/?<�o�.e�>yJ�?��>�X?FG�� ��x5پnĵ�� Ǿe��k���О>��[=U��������n��	u�J��0����>���>*V?�a�>���>hđ>��z�&� ���>��b�'c��1�I�%�u���ʘ����� �Kq���Z���]�>%施�`�>�.?A?>ɳq>���>1{q���>�p >�2y>L�>��S>�+>���=�E0�q���KR?v���!�'�$������2B?)qd?�1�>ni�M������#�?���?,s�?�<v>h�I-+��m?�=�>#��Bq
?�R:=�O��N�<]U����D5��0�R��>�G׽� :�sM��lf�jj
?�/?��y�̾iA׽�_�s=���?ȣ(?2*�rUQ��o��V�@�R���"�#re�B���z$��p�cԏ��W��0烿�.(��`6=F�*?�?���xH��A�k�1I?�_�j>��>ت�>���>�
J>�$
��$1��6^��W'��/��9G�>��z?�.�>�I?'�:?�dQ?��M?���>���>h�����>;R��>\v�>S�8?��/?/?�?S�(?8�N>�i
�������ھs�?�?��?�t?�
?�y����Ͻ1t��P#�c2}��Æ�"�=���<,�`\v�I�q=��Q>�S?5%���8����ji>P�6?n�>��>���R������<�D�>�z
?L��>� �,�r�����|�>��?y��q3 =3E*>.<�=����R?	�d��=�M����=*u�h9���!<�5�=��=l^X�m8�9�A;�zo;���<�-?q�#?��>�?W>��m�Li)�H�s����>?S� >���>ޢ�_!��5Y����"��K�>Pr?RI�?��=�'>j�y>�]����о�Z��Hv>�?�g{?��u?�v�?b�?�<S?:x�=.}��9��0+��
q\�l9�>2!,?���>�����ʾ����3�қ?:a?�<a����3)��¾� ս�>Nb/��2~����:D��������▙�c��?���?PA���6��k�^���|Y��`�C?�!�>uT�>g�>�)���g�Z��A;>S��>~R?��>'�O?�@{? �[?=�T>�8��!��i֙�q�6���!>�@?ê�?��?1y?�r�>�>:�)�^0�-W�����*�؂��'W=6�Y>4��>�0�>���>0�=~6Ƚ����??����=gb>�v�>���>G��>Ʉw>�V�<��G?r��>�&���a��$���L���PB�ܗu?Ţ�?��+?�c=����!F�̼����>�[�?��?�s*?�RS��k�=��Ӽ�����q����>wǹ>J�>�S�=r�K=.>w��>�"�>�8��w�'8�w�M�_�?F?���=/ſ��r���e�^���;<E����g������I\����=Đ���D�W$��4�\����.$��hq���E��r�|�i��>�$�=��=
�=L;�<����1ǰ<f�E=��<���<�@i��N <6�1���ڻ�G���.;IS�<�6C=�1*�d����w?�M?��=?�L?U̓>RT>yV½�K�>mܽU�>�">o]}�����Ò��s���A��Vo�ܾ7e�#��t��= i�&�(>��/>6��=�%>��k�=�lK=��;=ؔ�;�.)=��=���=��<��=d�>�N�=�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>ڳ7>�$>X�R�p�1���\�|�b�}Z���!?5J;�PO̾�?�>��=n+߾N�ƾ��-=�e6>b=S\��N\����={{�|�;=��k=	؉>��C>���=3#���޶=�I=��=��O>< ����7��,�$�3=_��=ޫb>N&>l|�>��?�b0?�hd?I�>�m�Z�ξ�d����>x��=���>3τ=B>Y��>{�7?�D?o�K?�3�>:T�=0�>�ݦ>_�,�ԝm��f�_Ƨ��@�<���?�ʆ?��>OV<�SA����i>��Ľb�?�]1?S�?��>>�
�rgܿ��5���,�g< �%��=۝�>��:C�����;AM���z>`2�>�$�=3�>m��=�>�=_\=C�=Z��>�W?>���=K�#>���<QA��\<�X�<���ʳ�<$�̻�פ���<vA��(=�伾s<���{a�=H��=1�>��>b(�>�=���m��=3H��6�H�Vh>����39�oi�b�}��C ��)��p>�؍>Vks�Ɇ��xK�>���>�_	>@u�?C�?V*�<8M�d&޾�Y�������I���>�U>��b��}=��g���V���a�>Q��>p�>$�l>]U,��O?�m�w=�
�B�4���>P싾���P��:q��(���П��[h��D�9��D?�%��ש�=\X~?��I?<��?5��>�����ؾ�D0>hま�=a��b|q��疽�?�,'?��>����D���ʾ�۾���>�GJ��`P����{�/�n��e���ɲ>Ӑ��mnо�f3�<���4L��̛B�k�p�+��>��O?��?�>a�'���:N�� ��j����?�;f?!��>�?7�?���z���:�=��n?�r�?�A�?!�>���=z�)��9�>� ?ˑ?:��?D�?�ா-�>_�=���=NE����">��`>�>�M�=>�?��>�]�>T鸽�P��	�Q���4��<j��3�=餞>{ڞ>ܸ�>��R>T�!>��"=��>�>5��>�q�>���>���>�&��p��@H?0Ϣ=րg>}�0?7|>O�=/�뽑.�=�ol�t�s���]�����̽,�:��=�u>�O5��[�>�¿��?��7>�ݾ�0?%u�F���>0>N��=Z _��>~�f>�9�>�j�>aZ�>�
�=��J>n��= �Ǿ��/>�s���$=S��k��Ծ���>	M`��;�&��@?�����5���x���X���i����r�O>��?��9;�7j�a���� ���>��>�^?�ԍ��^�<y�E>��>k�6>���O���Е�zz��l�?��?~�h>�k�=�ˇ?CU?[��%:�;v{�{w-���L�g�s��cQ��_������ع%�r
M= �?_��?=�U?�� �>�?2N�3��;��=�y^�ұ7��u=W��>xPؾ@=4���
�G����R�&�>m�q?S'W?�k?�Y�+���>�>&?�	1?iɀ?��D?3AJ?A�Z��?� )>xN�>0b�>��(?z�-?�	?�5�>%4H>����UV=�P���떾�����k���<��=�.d<7vl=о=����� ��� ��$λ^,�<e���J�<��G=4�=tU>f��>̤]?:J�>���>��7?m��Kw8�/®��0/?+�9=���\���ʢ����>��j?Q��?�dZ?+]d>�A�c	C�>Y�>C^&>�\>pk�>���ϖE����=�D>Z>�ϥ=cYM�;с�?�	�͊��0��<�+>���>*0|>e��`�'>x{��a0z�̤d>��Q��̺���S���G�1�1�΄v��Y�>��K?[�?���=�^�M1��JIf��.)?.^<?�NM?M�?��=�۾|�9���J��>���>tA�<������v#����:�?:�:�s>�2��xޠ�=Xb>����s޾ޛn�J�B�羚>M=���TV=��t�վ^4�ɣ�=�$
>?���K� �#���֪�Q1J?�j=ax���bU�6q����>�>�߮>��:���v���@�R���Y6�=ӵ�>��:>�_�� �~G�>8���>�<??i^?�x�?�����T�р1����$���=��?.��>��?�0A>�P�<�3�v� ��h�����>���>*�E��'G�
S��V3�4�N�P8I>]?��=��&?�k?;�>�b[?�~^?�%!?q�=_����R�B&?*��?�=K�Խ�T� 9��F����>�)?C�B�<��>�?Ͻ?��&?хQ?k�?j�>�� ��C@����>Z�>��W�yb���_>��J?���>S=Y?�ԃ?��=>��5�v颾֩� U�=�>W�2?�5#?�?﮸>��>k*�����=�<�>�`?�~�?�H�?�M/=���>w<>" ?�A>?�>P?J�?��K?PMh?�z<?��>4�=�O��]���$C��E�<ᩞ=�ޱ=���<U����(���ݽ$g�<U'��^�i$=.�=��=!��T�=g�>\�s>�Ӗ�N�.>@Kľ��"<>:����J���ዾ<�<��n�=8�}>��?�ߔ>�� ��I�=�ռ>�>�v���(?��?*�?�k�9 �c��ھ�H��7�>�lB?�6�=,Wm��ᔿ��v��%]=�|m?��^?ߢP�������e?)�b?��ܾe�<��^���e��r�Z�B?��|>䯾�{�>�r�?�\?�{
?=�=��\�~l����n�rE��(|=��>�-�<�����>7�"?tq�>3E=�Z:>�&۾�.v�􆙾�?�
�?�R�?��?��<��k��*���������@?~��>"���}�?�⭽�����p���D��>���
橾��n�"敾���H?^��گ�;>� ??�Mj?L[X?6
�
�q��yc���w��KM�Ý �bQ�;�W���V��;N��Sp����j���i"6�4c^=��N��G��b�?�)?ό���a,?�?оn�����F4v>�2��!k����w=#�Q�g�>޴�=�'�kw��(���?#&�>;MU>��2?����/@��l�E�򺍾��C>@��>�ץ>���>U�=V�H������a�\�j��jv>�qc?��K?H�n?B7�9�0��[���o!�9�2��y��
KB>�
>���>sW����]&��e>�4�r�Х�b��5�	�7�}=��2?��>��>�,�?z�?r	�󕯾x��X1��I�<C%�>�"i?g%�>�ˆ>>н�� ��?�v�?�?
�>���$6���L��M?J5�>��?ѝ7?�<t>	>F�7��衿�����N���Q�F~z?m;�O�l��"�>D�*?S�*=��?>�?����T�d�:�Ͼ{�Ǿ��� �?�,>���<�T��3�j�X�$V=�K)?�@?:Β�\�*�{~>�"?{��>M �>�%�?��>þ����Ө?��^?71J?\8A?6�>�q=}��mȽ��&���,=�>�[> n=ϔ�=S��Ö\�����D=��=_�м�L��-<Sk�� ~Q<Gq�<:4>��ؿ�1G����P���辵{�}�����1���$(��ػ�xߤ�bz�n��&����;��aO�������E��S�?<��?)·��|�t������J��ٰ>�,q�ч��﮾3uE�L᯾��� ��5��d�>���T���]�P�'?�����ǿ򰡿�:ܾ5! ?�A ?7�y?��7�"���8�� >aC�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾}1�<��?7�-?��>Ŏr�1�ɿc����¤<���?0�@RpA?�{(�r���3X=���>��	?�,B>w�1�P����� �>�!�?Ê?GCL=?�W��'�'=e?�G<5�F�R$ٻ�1�=�k�=m=L[��YJ>��>��@�W�۽<5>+��>��"����v^����<�-^>N�ӽ����5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=0q�����8�2�?[!�'��=U�<
��|���ތ�3眽Yw��H�i����C�>��>Oah>6S�>	�2>͂�>�iX?͜�?���>"��=G9i�=�����%� ������������tk���о�߾#X�!��a� �
k�6wy�� =��=�6R������ �4�b��F���.?�t$>��ʾ*�M�<-<�pʾ����ބ�:ۥ��+̾��1��n�W͟? �A?�����V�`���������W?'N�l��cꬾ@��=�����w="�>���=��⾽3��}S�n0?,?KD�������+>i����S<=7�*?M�?�Hs<q�>-�%?1A)��K⽊�V>P->a�>�>B8>����,Y���?ZT?Px��Q�����>&X��#�z�3�f=�>��8��~ټ�l`>��<����� �uф����<��V?��>�B(��	�#��t�?��=�x?۔?�Z�>��l?�	B?��<�����RT�O�
�ߧj=��V?�6h?��	>�H`�E�;�g���6?�c?��H>��[�;��~�.����?3�m?�?r���D~�Jؓ��	�e06?�mb?��;�� ��d����]�>=��>�P	?�jf�h�>�v??f�=>O���dӿ�X�aà?�+�?���?���j�|��=*?��>v���kۉ�06�ێ��ཷΡ>�����t�&�о��=�M�>�1�?�Pz>�=��������=(�j�?�$�?p�ľ:`e=�W��It�#��d�=ρ�=l(��=��4ؾ�,�ˀ������I�����s�ڬ�>��@�mN����>�nh����`CĿ�v�o����Q���!?|/�>�鮽�}���St�U�o���8��	C��]��J��>v5>u\��!����z�L�?��ԝ�H9�>4���E�>N�_�e@��4Ъ�1{����>���>b��>�f~�Rx����?���+�˿�E����|�Z?�"�?�ʅ?�?�<�j�N�Z�o܋���??h7q?mW?*-̼?�O���?�!�j?y_��]U`�ގ4�rHE��U>�"3?�B�>b�-�E�|=�>j��>Fg>�#/�z�Ŀ�ٶ�H���M��?��?�o� ��>i��?ks+?�i�8���[����*�4�+��<A?�2>����M�!�50=�8Ғ���
?M~0?2{�i.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>gH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?��>(�?���=&��>���=Z,��Ae��Z�">uz�=�s?���?j�M?���>#�=�Z9�\:/��E��R��3��PC�3�>�Fa?6�L?
�c>?��'7��� ��ͽq20��	�ֹA���*�;�ٽ�%8> �?>@Z>�HB��+Ҿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Oz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>B�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji�w?0% �$���@l]�t}��������=8@?�_���>Qq�>�9�=�ӄ�Y�����]�:�>Bp�?	C�?"��>R]q?�&q�0�7� �;0��>W�w?��?�ba=�*���:>�"?)̾|h���}���V?r�@r3
@��[?-��f׿�ꟿ���ͅӾ\�q>�'�=��>.i�|�Q>��~������=�5>$�>��>`��>�XQ>r�>y��=���&�5 ��u����
��f"�����⽹��(��A��W=����Ͼc4���<sQ*=U���e�*�j�\�ŊD>�6T?9�E?% o?I�0?x��=�>f'�m�S�,�ξ�|��ac>�?�+Z?<�8?-[<�H�Lw��Ꮏ쥛����Lv�>L�>�ԩ>��?���>GtI�8�=�w~>�T2>_z��˭H=@M��$C��8�<��>t� ?v��>�C<>��>Eϴ��1��i�h��
w�s̽0�?����S�J��1���9��Ѧ���h�=Ib.?|>���?пg����2H?$���y)���+���>}�0?�cW?�>��s�T�,:>>����j�7`>�+ �yl���)��%Q>tl?��f>�u>&�3�De8���P�|{���j|>�26?�趾�G9���u��H��aݾ�KM>Pƾ>�D�sl�����
��vi���{=6x:?)�?O2��|᰾a�u�4D��sQR>Z:\>uP=
e�=!WM>u_c�6�ƽ�H�@p.=*��=�^>X�?o�.>���=�>�镾�J���>�m>>�=0>w�>?��&?�WԼ��9�����3��h>;��>NW}>�$>��I�݊�=���>onf>q����Jf�K��A���R>��l��#]�����Y��=p|��M>#n�=o�轧�/�}/=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>xx��Z�������u�u�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>:��?�gY?soi>�g۾=`Z����>һ@?�R?�>�9�~�'���?�޶?կ�?�7Q>j_�?wu?
��>1v���T+�����SH��7��<waƻ"�>���=���޽B����������.k�#0��7�>{�-=ȭ>+����g��da�=
�⠵�8�D�{m�>�W>��W>E��>���>b��>P�>c*=��iҀ�磢�> C?w��?gU�`�}���>���=n��&�>��?�ҥ�/��Wt�>�U?=z�?��u?��S>Nl=�m���oۿE鵾�����>%)?�'?dث�)ٲ>��¾.Tn<A�>��>����
վ�':�3J��x��>�8?�tp>��Y=QN?�3,?I��>��g>�yR�=��&O����>��?��#?��?�M�>Xt��T�!����
��:�L��xH>b|`?*�?�`�>�U}��B��`��=#B-�kS<�W��?q{Z?�*����>�?�?n�> 05>�Y���*��_d��M�>��!?�����A��;&�����x?%l?	��>�I�սxNԼ���`����?M\?8#&?ݘ��%a�*
þ���<K1'�atW�}<}zA�*�>.^>�����}�=�&>Ű=ym��)6�o5k<f��=���>ǔ�=l�6�[��R�"?׶K�������>@ƃ�kBK�n�V>5f�=��
���?���x���>=��Iߗ��6�����?L��?l��?���Vwb�o6	?g��?gW3?�Q?�d������� �3�ɾ��[�|��V� ?�Ւ>��V����?
��������=�_ɽx �>��?|?į?S�>�g�>�ɽ���9����3��_d�;y;����%��1 �3Ež�K��z��=�G�����d�>8y;��>�V?A#>�d�>#$�>�N���f�>�#b>J�c>/��>��>r7>�g=k͐=���GR?*�����'���鐰��/B?�~d? �>�*i�<�����dv?��?)k�?fv>c�h�F#+��_?~4�>���V
?�:=uk�K�<�3��~�}y���j���>�J׽�:��M��f�`
?n8?_k���U̾׽Y����o=�N�?�(?04*�(sQ���o�1�W���R�9��Og�����F�$�lp�����~0���܃��;(�i�%=y*?�9�?`(����X��myk�%�>�vnh>��>zf�>�2�>�+I>��	��s1��J^��4'�u�����>\{??�>��B?t2?oZS?AP?�\�>�]�>>������>P<|��>B.�>��2?I/?��+?x?��%?��Y>	s��z��9�㾼�?�?�"?��?���>񙙾9��Q'��>��Ǝ�fh���>^��=S1	���ؼo�=w�x>Ё?o`��|7�������m>26?N
�>���>�ۋ�}}��=�I�>�	?M�>)� ���r�/.�)��>	�?����x�<$D%>��=��&���Y;j��=Iɼ�J�=I�5�|�3�r�U;���=f\�=�<ο�;gL1<1�D<Xڼ<'�>�?O��>��r>a��
O ����(�=%�>)!�> �>�f�
v��B���aLg��Xa>��?VC�?N�<ǐ>��>>����� ܾĵN��7:� ?�M7?2,S?�ؖ?z5??�M?Ft4=�?�(�����,����Q"?j!,?��>��*�ʾW���3���?S[?�<a����s;)��¾��Խα>M\/��/~����^D�Y������������?x��?�A�0�6�8w辄����]����C?k�>iW�>��>��)���g��%�r0;>���>{R?M$�>��O?�;{?�[?imT><�8�`-��vә���3��!>@?B��?i�?�y?ts�>��>$�)�v��R������₾3W=�Z>	��>�%�>��>��=��ǽ�K��q�>��U�=��b>9��>���>q�>��w>>=�<�Z>?1{�>c�ܾR�о�۷����*G����?@�x?yD?��I��'Ѿ�n�S.2����>��?�ű?��L?c
� �P>�RԽr�����W��>ԝ?�֛>�l�=}����=��?Ht�>u���JM���C���<3�?v�8?�v'=�ƿ��q�C}q�/��c�m<����X9e�?���GZ��U�=}ט��]�Xz���B[��\���A��Yĵ�M�����{����>�Ԇ=���=v��=���<��ȼ�e�<�BK=Z�<��=�.o�!�i<�;:��ѻ����;�$���[<NpI=x��/����x?v�<?� (?��??2�q>�3�>�Rp���>����?I�z>`mT��*��#=\����������վ]Ӿ�U�>���=��*�m>�)>޾=D�=��=��=Ğ�=��n��\7=�-�=}�==�=�7
>�m>`>o6w?����s����3Q�g�s�:?9�>]{�=�ƾ�@?$�>>�2�����fc��+?���?�T�?��?�ti�}c�>i��r؎�^��=s����92>���=�2�X��>]�J>Ƀ�K��Հ��64�?R�@��??fዿݢϿd/>�7>��>�R�`�1���\�ZLb�+�Y�&�!?�E;��̾�Y�>+M�=�i߾��ƾ�,=R�6>�e=�k�!=\��=�2{�N�<=7�j=J��>*D>N��=2尽�Q�=@lH=��=.8O>�A��Ģ5��-���5=Ro�=��b>Ȏ%>!��>Q?rZ2?��Z?ρ>�7�>���?cܾ�3�>��>��>�f�V�E>��>R6!?(m-?�1A?g��>��<���>�`�>pkI��yn�Hg߾�)㾺��<x��?o��?�8�>{�@>r��n��3�Xd�U��>	u&?*?�Q�>��r�ۿ�����w����>K�=�0�Rnk���>����m�о�)C>���>j#�>�?���>[��>p�t=��>æ�>t#>k��=�Ul=�J��e1=3�����'ro��>̧�<��z�BBE=�y=t�ս�^ؽ@;��3�!<�̦=��=Va�>.�> �?�=V���%��=N�˾�O�X�d>��#V���U��=d�Ȋ.�F�"�z>-;;>���<�8���`�>f��>�� =;_�?ǯ}?��=�oս��ž�@��˳p�M�4��>~�d>����a��@��e`��и�)��>�>�%�>�ہ>�+��x7� ٫=G}ȾJ�=����>�|��w1��v���j�����͢��Hj�3�� ,P?�;�����=nt?UPB?�=�?Ob�>9㰽~�;��>�9��(X�<\��dB���
m���?�9?�(�>^��&�@��о��Jh�={��t2�s����/9������苾d�>�c�70�m_`�a���pDm��X��o�'<G
?6�K?���?�L�T8V�*�ʾI��]�q�1?c��?t�>?�U?���>x34>�\*���5���4>�6?BR�?���?�.m=�H>��=�Q�>fA?���?z��?"��?�q۾��>����V>��g��D>��V>C@=y���0�>ޤ>ҷ�>����'	��>b����Y
���н���<���>b�>Y
�>#8>�b>��f�r)[>��C>�a>G(?Mv?�ak>�Õ�nJ�,�E?U>lH�>]�D?%�>�0$<��!�ܟ=:�꽶貾��ǜ��ʥ�u(=�=j5�=}��<$�><u��"�?u{�=hQ	��d;?>���;���>Ĳ>�g<���>>�E>jy�>��>�v�=�M�>�4i=�EӾ��>B��Pd!��,C���R�i�ѾL{z>ě���&����x��HAI��m��ug�[j� .���;=�Ž<�G�?����n�k��)�Y����?d[�>h6?p،����$�>=��>�ƍ>!K��l���5ȍ�bg�i�?���?�P>+��>8�Q?��?#�=��>��t]��v��<��?a�/�^������5����½G�\?ev?Z�??�N�<���>.��?S�&�5.���(w>�N9� �4����=��>����!L���۾��ѾH�<�S� >��h?$��?�#?�V�tk�<)�=
? B?Ck?@	-?�$\?��5�8"?LOb>5r?�;#?ܚ3?�I<?�?ց >?�> +=��[=ͭ��V���8�p�,���i�;?��=n�>=�\�<�ތ=��=�L�<�{���T½C�,��0�=*��=�xH=Y5�=ؾ�>ؤ]?�L�>���>��7?)���w8�LƮ�V+/?��9=���K��'ʢ�����>��j?� �?�dZ?�bd>r�A�
C�>X�>r&>�\>�d�>�{�G�E��=�L>�X>ƥ=�bM�Fρ��	�v������<r&>���>DI}>����=*>B�� �w���e>�kT���qU�[�G�� 2���u�M��>i�K?�N?��=ނ����$f���(?��<?oWM?��?)Q�==g۾q\:���J�l��(�>*&�<�F�哢�^%��K;�L�"�t>�5��γ����b>N���A޾�n�?�I���羈�N=��)FT=� �-�վ�~�7�=|�	>t���8� �j���ª��)J?�k=wƥ�A�U��>���6>g��>z̮>r�:��w���@��l��{��=��>�;>� ��-ﾗtG�m?�x*�>@�E?8x_?*(�?�+��8M[�1�;��Kƾ������n(?t��>��?TT>jk=9nؾv3�vOY�*E4�]\�>_�>��7���F�<gZ�����Y�*�y>ޱ�>���=��>��[?Y��>21V?QB(?�>�^!>�2н�;UB&?��?e�=��Խ%�T���8��F���>G�)?}�B����>�?�?��&?�Q?�?N�>� �UB@�Ɣ�>*Z�>J�W�`b���`>b�J?��>�;Y?Nԃ?�=>q�5��⢾�ϩ��a�=�>j�2?�2#?^�?���>�y�>�����=���>�b?L�?��o?=
�=@�?�1>f�>���=S��>�<�>�?fQO?�s?q�J?H�>�ӌ<����[�����r���W��M�;cMN<�w=��ów�``����<S�;g����q�����IE��L��(�;�]�>{�s>c㕾s(1>��ľ'���
A>�祿NF���芾�:�R�=�u�>��?��>s#���=���>�C�>���<@(?��?�?v�;Q�b���ھL�K�.�>�	B?���=j�l�2����u�ʐg=��m?|^?�sW����TDc?{Xg?�����J����J������K�S?6�>,��O�>�$�?K�?�X?;&��p��䢿e4S��̊� ʵ=�i�>$�1�p��[{?�?=~�>���=�&>��-&s�OY[��L?�Ρ?酸?�Z�?A!>N~����Ͽ����t���CT\?���>m����-!?�Q��"о����j�����w��~<��
8���ʥ�WF%��O���ؽ�+�=R�?|s?�dp?�_?]/ �$�d��O_�O~�U�e�����E���D�V�E�R�o�o���x��`噾#C=a�D�	#H����?�+4?�U�.$9?Tc��H���3Ҿl��;�2���@��Jh�<,s��n�b>�*1>���^6=j!��D[ ?f�>D��>��B?ޠ����6��W;%Q���Z�]S�=vVU>u�>	 t>�>l=�=:;�=�޾<��}>�=Dw>�bc?j�K?��n?p���c0��T���� ��l/�p˧��!D>�	>�>��W����6p&��	>�3Tr��%�_o����	��=)2?���>���>�ܗ?�#?B
�X���'x��1�*�<���>��h?#;�>t�>,ӽ�� �bI?�Fk?}"?�>3x��! ���%G�@[>�?��>��"?���=�~�=��5����Tjh��%�h49>��O?I�i�eΆ�ථ>��*?�t��~�>93>i�<:6o�9@�l�P� �A��8?�E;=�}*>]��〓��f��彔P)?WU?	Ԓ� �*��<~>"?�x�>�#�>�5�?�;�>�Kþ��)��?��^?1J?�LA?�$�>��=�O��DȽ��&�vZ-=���>��Z>a�l=��=���/�\�Tv��bD=�G�=��μ�V���
<􅵼ȫJ<d��<4>׿C�YAھ�����վ�������[�ٽ0���9�#Ƭ�jޛ�����tI�JK�4�[���F�鮌��ZT����?-3�?_Ʌ���v��;���Ԅ����/i�>��Z��{�6�����`g��Ql� �۾f�'��Q�~�h�cZ�M�'?�����ǿﰡ��:ܾ(! ?�A ?7�y?��,�"���8�&� >C�<1.����뾯����οA�����^?���>��/��`��>Υ�>+�X>�Hq>����螾t1�<��?<�-?��>��r�,�ɿa����¤<���?.�@{A?�(�ۑ쾢�V=N��>�	?�?>�1��I�����[�>�1�?@��?Z,M=�W���
�Wqe?�<�F���ܻ��=�ʤ=��=&��cJ>)N�>�y�~dA�"�ܽ/�4>��>�5#���Jt^��A�<�M]>��սO|��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?5ۿ��ؚ>��ܾ��M?^D6?���>�d&��t���=�6�ֈ��x���&V�w��=W��>_�>Â,�ދ���O��I��[��=����'����$����7�=�]�<a����tP������)�aU�Z�w��b��=Ke(>�[C>Et>
B>�>WO?�9r?S�>ڲK>�r��W�����=�r��D$v��ϟ��TW��R߾�+�=�;�9ھpa;e�׾C ��=���=�4R�a���� ���b�ٚF���.?�k$>h�ʾB�M�{v-<�pʾLƪ��������,֖̾1��n�/̟?X�A?���!�V�j��-��ە��7�W?�H�!���ꬾd��=d����Y=��>�u�=0��� 3�a{S�~�1?�M%?�Y��Д�b��=��@��#�<^?/?mZ ?g��=���>mZ"?�04��7��#>�`8>�#�>:C�>�+>����ԃ���<?��T?��>�Ni�>��̾g�����0=&�=�<�BD����?>Bv��'��F�ܼ�ֽ��:=yV?�	�>/$�������ٲ��ؓM<p�}?
�?���>�v?�<?��[<y�_�P����T�=BZ?�Eb?+�>tL��x��*��TL-?E�X?x�M>C�p�w�ξ~A"�oy�.?� g?(Y?�02�y�"5��͌��4?�p?�F�K���a�Ҿ�ԝ��_>0�?4��>t�(�E�>hkL?Z�Y�7���Ѥ����:�05�?�@C��?L��=~yC��_]=��(?��?�c���ľ�*�=�龔�3���>���Nl���@��2@���N?�k�?Jn=?ⅴ�����7Z�=u|���Z�?��?ۛ��'�p<%���k�9~���G�<���=;��$Y����x�7�PCǾԹ
�Z����P��>TB@������>��7�
3��+Ͽr���JOоp�q���?��>�ʽ����2�j�� u���G���H�$���P�>��>އ���둾'�{�2l;���b�>[���>��S�m/�����5<6�>���>㹆>l��潾�?�Z��{?ο̪��I����X?Zc�?�n�?kp?��9<d�v�ā{�uA��,G?��s?�Z?��%�8]���7��j?M]��V`���4�*HE�3U>�3?�L�>9�-�]�|=�>���>�N>=$/���Ŀ�ն�	���t��?��?�h꾰��>~�?�r+?h��4���N����*�pp!�O;A?(2>�����!�.=�pɒ��
?�0?vT��0�Z�_?+�a�D�p���-���ƽ�ۡ>��0�f\�KN��&���Xe����@y����?M^�?h�?���� #�d6%?!�>X����8Ǿ?�<���>�(�>*N>�H_���u>����:�i	>���?�~�?Rj?���������U>�}?���>P�?�+�=��>"�=�հ��x4�0�$>S��=��9�.�?rGM?0J�>�&�=m�9���.��=F�ѲQ�����[C�Ȯ>F�a?yOL?9[a>��/1�O� �XҽW3���F�?�.�3�� 4>.=>Nx>J�E�JgҾ�?R��ƿ�q��߇��"@?��=D�,?;�����$ؽ[�q?�B=��u�������<����?ń�?wQ ??����N��	>mم>�(�>����c^��h��O=>=Je?s�9��h�4WK�c�r>�x�??�?���?>���d?2-���.����u����?/5�eC>C?_��é>�?�� >\	s��ۣ���~��>�ԣ?w��?��>�&V?��X�&.��h�=�.z>��N?3?n]^�����vy>�<?ij��ሿS���-wh?@m	@f�@H�f?�˘�qjп�L��g�a]ؾ��=�)H<�6;��O�M�>ɯ=���¨=�9>�c�>�@�>b	E>�n>�)�=x�=���&�*��y��Ɩ��qn����v,���f�������o���𥾢���%-�P(ν�#��@���6#���:�*>tb?a�6?�%e?��L?נͼnV�>T{1�Hӽݶ��0���cq^>�O?1Ig?Q�6?�l>+ܜ��̈�r����������|�? 4�>ğ>x)�>�Y�>,
:�x�b=PM&>��k>����6=	����b���>�I>��>�?�C<>��>Eϴ��1��c�h��
w�i̽0�?����T�J��1���9��Ǧ��i�=Kb.?|>���?пe����2H?���w)���+���>}�0?�cW?�>��\�T�':>C����j�:`>�+ �kl���)�}%Q>nl?�f>�u>̛3�ne8�Q�P�w|��Bj|>�36?s鶾QD9���u���H�`cݾtHM>�ľ>=D��k������-vi���{=fx:?�?7���ⰾ`�u��C��PR>y:\>U=i�=�XM>�bc�<�ƽUH��f.=Լ�=�^>�_
?��t>��=_�>�U���M��:�>�t�>iT�>O�P?�.6?H���T���<��Z�]�|n>�p�>M��>`?>cB6�֛�= ��>��>�mQ�M8��"gӽ�n��?	>���;��#��KDB=ä��re�=B�V=��l�*|�=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ\O�>ښ��葒���~��cr��Y��1�>�^N?VS����=�����?���>�b�֕���qҿ>�f����>���?���?�qc�^����C�K�>,��?�`!?�>p��*�i���>R�]?%�?�j?Ȯ��o�>9��?��m?�K>�.�?��t?�:�>�P��C�+�Fm�����ɻm=�ה��_�>�E�=����E�c^��1ʉ��i���L�d>#I'=+�>��������=b�������;f��:�>��d>KF>1D�>}��>c��>�U�>
=)������@+���QM?=W�? ���'m�n??�2�=�E�U�k>`%�>8���^A���>�:�?Ց?G?8�>?e�w���ӨԿoڴ���ǼG�>�?P�?"U��%�>��"���	����>^�>�9/�Ǭ¾Z���0�c��O�>J'?�4>�'!�'N"?p&?Р�>bL�>�=�������?��@�>���>��>mdu?W�?[~��A2.� �������9�\�!71>��l?�\?�(�>g���Nz��ێj=K��'t�Qvt?nX?�� ����>;��?��/?=�=?G6�>}a�}&����g�=>��!?�/�A�O&���}?4P?Q��>Y7���ս�jּ���X{��2?V)\?�@&?���r,a�� þ=7�<��"�jU���;�?D���>�>���ޕ�=>а=PRm��F6���f<@m�=#��>�=�57�,���%?n���)5��2>�>�9i�S#�{ ?uc�=�(���W?	�ž-K`��紿.���	���~�?x��?!*�?�IA��_�W��>ﭞ?�?�>�?E�w�z���"˾�״�4��j|.��b��&?��3=��U�����$����&d�n�[����(o�>��?�D?���>+ޝ>u��>��q���/�]������k�=���L4��T � G�)�@�ﹽ���k4ƾ�����ɇ>x�=�>�=?�[$>7�>��>ĸ�9��>w>��m>)��>!�`>�p>=D�=s��=̝��LR?��� �'���辀���'B?Sgd?�7�>L�i�i������B�?���?7x�?f�v>�vh�35+��T?��>����v
?�K:=��-;�<�9��º�a|���6�;��>��׽ :�M��8f��p
?9?Oь���̾�ؽ�¾�7�=�_?7?ʔ�ck�8ю���I��?�F�k�ځ:������-��2���r��Uq��()��ɚ=XR0?���?��쾴���_þcu�Js����>ғ?���>�q�>�M>��۾1�I�=�}�Ə#�4����t�>��y?���>��I?��;?�wP?��L?��>�>������>r��;*��>�i�>�9?�.?�0?(?+?��`>���N���̀ؾ�]?��?y�?�#?
s?fu��o�ƽV���e��gz�>=��jD�=�<%`ٽ`�u�$�P=!�T>�X?`��Z�8�������j>��7?Dv�>���>���0���f�<��>��
?EA�>t �O�r��a�}R�>��?����=y�)>���=������ֺxT�=J���;Ԑ=�����};���<�Z�=E�=��t�x������:��;�<�#?;�?Z��>M�>�/ξ.������:�>�
?��>��>�	%��ꁿ�!s��<��G�>a��?|ҳ?��	���>&�>����/�dw��{���&n�.�O?&�^?�r?���?#�z?H�1?T�=+X*�Z��v���=���p?v!,?��>�����ʾ��Չ3�ݝ?e[?�<a����;)�ސ¾��Խ۱>�[/�f/~����@D�s���[��6��?�?SA�U�6��x�ڿ���[��y�C?"�>Y�>��>U�)�}�g�r%��1;>���>mR?-/�>�O?�O{?��[?�T>!h8��&��<����}6��!>�@?��?���?'�x??@�>)>��)���������,��V==�Y>�t�>��>nߩ>#�=�]ɽEm���>�;��=�[b>�w�>�z�>��>D+w>+v�<b�G?��>L̾��
�b����ȃ��3;��Vu?y��?��+?�=��h
F�1 ��5
�>qg�?sܫ?�q*?0�S��>�=?�̼�J���s�	��>*��>�M�>�I�=��K=��>���>���>����+��8�-�Q�h�?��E?P�=�Cƿ5�s�3�{����r��<c���tX�Q�����]�j[�=�\��<��I����HP��2���~���������gr���>gՖ=e��=���=�l�<�?�k�< 1=�wW<�"J=�2���<qOU�`�ڻ�]��
<���<��>=~�;��Cʾ�e}?��I?r�+?e�B?.f|>�b>7{'����>a����g?�CT>\HA��`���<����Oꔾ�;ؾu־��c��o��Bs>�}N�`X>y3>���=$��<��=?+^=�Ǎ=b���=��=p��=`%�=���=*�>h�>�5w?N�������h.Q��m�/�:?�B�>1v�=^�ƾ�@?W�>>1������c�+?���?VV�?#�?ni�N`�>��򫎽N��=�����A2>��=�2���>��J>>��6K��o~���2�?i�@{�??�ߋ��Ͽ�Z/>/�7>t>I�R��1�0�\�o�b�n|Z���!?�H;�yF̾:8�>��=�-߾�ƾjd.=
�6>�_b=za��S\�s�=��z���;=Pl=�Չ>��C>��=�7��J�=�I=���=1�O>�8��F�7��,���3=i��=!�b>�&>5#�>,�?�e2?8h?�I�>!^�B	þǾ�d�>�)�=�e�>�O=?h0>>�>��8?I�G?O�K?e�>/��=��>b�>M�.��;j��������<��?l�?�N�>I%�<�TE�Bi�_�=�ܫ�b?#�.?��?ǈ�>aP �xο�:��$/��u�<P�Y>��F=0i�G���a3�.E�=/G�=q=���>�]�>3[=�#Ǽa�
�|R>��>�H>ۛ��a�<���=� b= �>��<�K��>��=j�ㅽ������Ƚ2�˼�(=�5C=OI>��=A��>݃n>\��>;�^=$i��e�>Y����OS�z�=􆹾�G��X�J{��m$��u��>�@s>ƀ���ҏ����>�Wn>�#�=�?x�|?Hq=���|Ǿ�蜿��9�.���8>�>jB��=���b���>�R����>�>G�>��l>m,��?���w=-��^5�p�>�t��k��E�^7q�?��3����i��"Ѻ��D?�D�����=� ~?`�I?��?i��>� ���|ؾ�0>�W��N�=��gq�>]����?j'?ӗ�>1쾦�D��pʾä��E�>%�J�7�O����j�0�?���޷�N�>����ξ�H3�~x���\���sB��Rs��Ժ>v
P?z�?��b��逿�VN����ڃ���?S�f?�U�>��?��?�������!��m�=�|o?�(�?ю�?g�>�)�=��Z��>[�?�֒?;ؕ?&d?��(����>yb��w>˒
�`��=o�=���=��>?�?��?�>�>�x���7	�/��,i꾏hh���n=cL�=��>�4�>�?>rQ�=�G=��O=��r>�p�>���>�S>�{�>ޞ�>(��R�^>?J�>E�>>J?vi7>�Й=� ��%;#�̽be���M�����0�� ^�=�J�=��=z���-��>-���L��?��->��H�?���B<Z��Xx>л�=�$f�W�>� '>���>ۢ�>R�>���=��>:�>�!Ӿf�7>����V	��P*��~���۾�?f>��e��E������f���CV���[�+��$h��{t�Rj=�/2>�+�?0h�:�`�� �G���_E�>���>)�F?�ǀ���=���9?���>#¾�h��l���`�ξ݇�?��?O��>C<h>_n?��E?ˑľ���<S�.��c�d$Z�I�d�P����%�������=�|?#�q?��Z?��;5�>nr�?�o6��h?���=�S��t"�=��=1�>��	� �����/b�nV��[:���T?�M\?O�?Q%E���l�tJ'>��:?�1?�4t?T2?Ct;?d?���$?8"3>+L?:]?C\5?��.?��
?�1>���=n�����(=�3��G抾 �ѽh�ʽR��	�3=�%{=(4!���<r0=ܡ�<)��wۼ��;�*����<2S9=t|�=���=t��>(]?�E�>G��>�p7?����8��ꭾ�.?;=���7㋾!F��x���>��j? �?aZ?�"c>~!B��tC���>K�>��&>�>]>�Ͱ>���f�D�kσ=Ң>�H>)g�=A�J��]��Ӳ	�����<�Q>���>��{>E)��II(>c}����y�Ңd>��Q����͂S�2�G�t�1��nv���>��K?��?7k�=龻f���Df�@)?(b<?�M?��?z�=+Kܾɼ9��J�t��.�>���<|��(������T�:�m�-:��s>�_���}��.ll>�b���Hq�x�S�ܞ��tǖ=��H�=����l���=��=�]+>�kƾdd*�0��j���q1L?B^�=�����S�������>��>�N�>д(<�R{�$TK�����'�=���>��>���� �ﾝTB����Cf>~�.?d^W?��e?X�m��{?�ѿC�?�Ő��3�����>��>��(?|��>:>\И�0��9S�4�8��z�>�y?�� ��d]��T�� ���#���=�f�>�9�=s�>5#S?�*?@D8?"W�>s��>o?�=��c�K$���r,?2f�?:�k=������X(�B�Q�b��> ?>G\�,e�>�k?�(?p),?�,D?�?�=�=`��y7��S�>z�>s�S��I��mp>�r??C��>nX?�z?�;.>1-��Y���}���"�=�)�=��1?�/?D�?2��>���>Oϡ����=���>�c?�? �o?
,�=}�?MS0>��>�s�=���>���>z)?;~N?txs?��J?�t�>�T�<V����K��&Ym�FbW�$�8;�x$<�4q=0��o�o�i�}��<o��;�<���y{��S�|GF�Qݞ���;*V�>v�s>��s?>���Ɇ���C>��|�r{�������-��U�=8�{>S�?8Е>�
&��̔=�Z�>�P�>����%?�?Q?�ب���_���Ծ9�W�f'�>�#E?y��=Ij����Z�v�*UJ=PSm?M�[?��J�y��U�b?0�]?o_�7=���þ��b�����O?(�
?~�G�o��>��~?j�q?;��>0�e��/n����Db�v�j��=t�>�X���d�2�>"�7?�F�><�b>;(�=�p۾ߺw�Vw��G?���?���?3��?9?*>Q�n��-����L��"^?4��>g3��3�"?����l�ϾhJ��q����
��{���-���S��Ǖ$�Ń���ֽ���=*�?�s?�Mq?��_?G� ���c�<^�M��>KV�v��'���E�E��C�-�n�V��@��v4��G={�����D�Z�?��4?~�����>�H����ܾ1꺾L��>��0�R'�?�>%!M=I�T>�i�=N~�������
?�@�>Vŋ>�?��'���/���Q��fR�����I9>E>�ڧ>.��>6x�<����.h�1K�Y-�� ��t<v>�sc?4{K?{n? � ���0��r����!�Vz1�)e��.>C>6�>��>}5W�4p��&��6>���r�'������ �	��2�=��2?�<�>�I�>�J�?�'?�	�񄯾i�w��N1�M�<cZ�> i?}�>}ӆ>"�ͽ^� ����>��l?s��>��>����dZ!���{��ʽ1&�>�>���>��o>C�,��#\��j��M����9��u�=�h?���\�`�c�>�R?)"�:��G<�|�>I�v���!������'�h�>^|?O��=#�;>�ž�$�u�{��7����3?��?����'�T��>�I)?iҢ> �n>1ux?��>�����9=�? Z?��1?Q<?��>.ǽ�qڽ�Ľ�	9�&r}=9Z�>��!>�2�m�>������ ����{k鼆��<��S�O��̚!<H��{��=i��<~�>Iڿ�N����Yd#�σ$��L%�|�A�~�\���A��^�$�����2���b�����%���g����oA����_{�?���?�ϲ�{�Y�o8���F�������>&Oo�
^�;��ľm<0�+Uža徤7}��B)��Gy��
���-i��'?:�����ǿ�����?ܾ ?�> ?'�y?���"�Ŕ8�^� >���<���X��-���%�ο���	�^?��>�
�6��� �>���>��X>~Tq>���F�~ �<��?@�-?���>V�r���ɿ5������<��?b�@��A?t4'���뾿Q=��>��	?ݷ;>a2�f~��װ���>�?%�?��S=�^W�ǖ����d?~�;�F���ջB�=?G�=&�=�����G>�p�>�����>��۽�0>²�>��$����2_���<�'b>��׽�M��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=n�@VֿZ�(�c@�`2�;%�=t|;=��ƽ�S�=؞`�����:��Х��ݤ�=)3)=�k�>"�>��>��>�q]?��o?✲>�]�=[O׾�����_��ՃP�EkξVA����>���ݣ�����澾ɞܾ��L��*��B��0�6��U�=�]�W��j�:�Gz���H�s�.?-I">g⣾+�K�N�ؽx���?������<`4�����/�4X��Π?��M?��~�<�D�s׾�Tj�r���6�M?6�o=� �g:����<���9">�(�>��R�����:�=�Z��]:?~�!?/�����^��~H>YU߽D���O� ?�`?yἷ��>"?���NV����7>V^6>��>�Р>
�=�ɱ�K�$��\&?��e?-U��rZ��b��>�{���������<2>�������$%>)�=�R�����C��=Kb=�bQ?��S>����ܾ�i��к��Zc>!��?|�	?��>�&C?f(?��d��O�o�"���7>�9p?��?ѭ�=������;ž��X?��U?�_>��>�վ�G��-�L��>\�I?�#?��<����Ũ���ľ]*??�v?�t^�Uk��.���SV���>�~�>��>��9�W�>Sd>?�@#��>��r���Bp4�駞?�@��?`H<�G��=�=h?��>nrO�� ƾ����l���r=[��>�����Sv�T���N,��8?[��?��>r��o�����=f�����?�+�?����-g���Ti�Z��>E=�=g��������e,�`U������Р��
�ׇ>{�@{�%8�>��&��ݿ��˿e����UԾ�g|��?�P�>!�s�eU����f�Hjq�ʹJ�f�H��0��RF�>�>>7��y㑾W�{���;�����9�>[e�� �>SIT�ZI��,ß��{1<F��>Yv�>~��>����آ��I��?�<���4οW���\�Q�X?�I�?�l�?�o?l1<�w� �{����]4G?��s?��Y?{E%�g�\�nZ8���j?a��)U`��4�7FE�nU>l#3?8F�>��-�j�|=�>���>bd>�$/���ĿYٶ�������?!��?�n����>G��?Gq+?�h�77���\����*�n�)��;A?2>����N�!��/=��В�-�
?~0?�x��-�\�_?*�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?h�?ص�� #�f6%?�>c����8Ǿ��<���>�(�>*N>cH_���u>����:�i	>���?�~�?Rj?���� ����U>	�}?�%�>�?5c�=A3�>3�=�ή���=��� >���=��>�b�?m�M?A��>�X�=m)8�G�.�)�E�WR�X���kC�z��>Y�a?��K?��b>o����?*�a� �6'ͽ|�/��ռ]s@��<��J߽�J5>M�=>Kk>��B��Ѿ7�?Rt���ؿc��74'��*4?̃>=?���޳t��/�;*_?�j�>�>�-��`&��������?xH�?�?/�׾�Uͼ:�>U�>?J�>.Gս����0s����7>S�B?�!�>����o���>p��?��@�Ю?v�h��	?���P���`~�k���7����=d�7?S/�l�z>���>@�=�nv�ݻ����s����>�B�?�{�?V��>��l?c�o�R�B���1=/M�>��k?7s?Qo����B>[�?��������K��f?��
@Ru@2�^?���Nֿ���kC����Ҿ�7A>�*>��P>�a���>d=�`��I㈽݁=W�>G�>�u>uY�>��>��y>
���r�$��$�������H�ԧ�8��Z�� �Ml�w� �9����ؾ���/���������2�}ƽt���V�=��b?>!I?��?d��>VJ>��<K(�$a-����1��=���>�C?��N?@ ?�>�<����u^�̻`����s�J�U��>06W=c��>݆?��>��><��=���={�>��u=�Ž
h�='�r=��/>���>�?�>T2�>J^V>L�w>�ý�ݭ�low���.���Ȣ?���c\#��ѩ�@��d��yY*>7�i?�D��9���й��r��\�9?^K{��W������=�
F?J�W?�>�0����M�)>�܀��)W�#�H�R�򈩾,[����>^�>�<f>nw>j�4���6�l~O�{���Ě}>��2?�弾_&L�AZu��,F���ྖ�9>d�>±��Z��Q���3Ԁ�=�l�B9a=6�=?�i?0����Ͱ��Ek�P��$�K>�fU>F�3=���=��T>I8V��hս��5���F=���=-OW>?�?&:>o�>>��>{���>;S�X��>`A%>W{w>�[?�f"?�X�λ��ԯ�������>���>�r�>�p> L����<?��>,4a>�ɽPҽ�M2��y���O>�y�2ـ�c����3�=��Q\;��=�K��2��>�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿph�>7y�PZ��*���u�?�#=w��>H9H?�U����O��>��v
?�?N_�������ȿW{v���>b�?e��?P�m��A��@����>��?�fY?Vpi>Dg۾�aZ�ي�>\�@?SR?O�>U9���'���?�޶?���?��H>�|�?5bs?<��>Ζt��.�5������r�{=��{;�Ə>8t>L�����E�Ws���)��u�j�z��h`>Y�%=n�>�>彆�Ρ�=�䁽V짾��l�z�>��o>�gJ>� �>n� ?���>���>�?=o���Pـ�0���?P?u�?m��B^i��xJ=$>�=�V����>�\0?�⾼�}��v�>�`?x~?�oN?�1�>�B�H���Dظ�ö����;��G>?/�>���>�ڽN�]>{��_�$�{i�>g�v>5OJ�5�Ծ������ޒ>�&?���>8*�=˙ ?�#?��j>|*�>~`E��9��1�E���>+��>!I?��~?%�?TԹ�[3�	��e桿�[�9@N>Y�x?`U?*ɕ>t���Ѓ����D��=I�����~��?�sg?�^彾?�1�?ƈ??��A?�)f>���ؾ������>�T#?����r@��T&���j�
?	� ?��>�a��E�޽[�_���X]�[	?��X?�{&?��� b�d,¾�7�<!�"�d���<�檼��>�->�zj����=�>��=��u���5�U46<F�=��>���=�@=��푽;,?�M�zc���I�=�r��xD���>�M>�j����^?ly=�c�{�qି�����GW�+��?q��?�w�?V����sh�ؿ<?�Ї?2�?�>"-���޾NV߾��w��\z���>oH�>��_�t��򧤿}U��'���x-Žm*�m�>Ѐ>���>^��>�H>�Z�>�~���lD�2�(���9�7��1"��U�T70����h��E�y�񻇾��̾`�����	?l�=:�>t��>�x�>|k�>֘�>ҡƻ��>�b�>���>�1�>�?>K�>�++>Z��<1����GR?���*�'�Ű�9���2B?�od?�*�>ji�����Y��Ł?Ņ�?�s�?�@v>%~h�;)+��n?�<�>H���n
?�`:=���(�<�T�����zE�����Ъ�>�@׽z:��M��rf��f
?s/?����̾vO׽�����n=�M�?��(?��)���Q���o�ѸW�	S����6h�	j���$�ԛp��쏿�^��%����(��q*=��*?s�?Ռ�q�!���&k��?��cf>�>'$�>�>�uI>i�	�>�1�e^�M'�`���=R�>X[{?]�>��A?nb7?�G?8�E?�X�>=.�>�x��U�>������>�� ?�U'?��%?f}?���>\?��>���'��"澻�?��/?�u?õ�>��?y���� �n�<�Tr=����(��01 <�y="�뙠�Q;�>�T�>�9?�.7��E7���ƌ>�`,?,��>��>a&_�t���$]μ�?�>V6 ?��\>�
���t��]⾽�?V��?8�laU<�w>��==�4��<ɁM=E�Ҽϸ�=����#.�}��87K�=��l=�|<,��:7��<�׍<��<@��>@D?7ҋ>�c�>钇�0K �GA���=��]>p\>5a>>�׾�뉿�D��S�h��}>H�?�U�?� �=�_�=f��=Aj��R\������x��<�=�}?	�"?�T?ŗ�?��;?�$?w�=�m��&���_��=���Wi?�5$?NV�>!wC�`�˾���B�����>%�>s�i��~��<��.��ǘ�;3R�P����?��聪��4��t3�v�	��4ֽh��?�E�?ϙ�=�ؾ�o��}��~�	��T�>�p�>�a'?��?�0W��ׇ��磾Sի>�>�>�J�>���>� Q?��b?�8?gѮ>����=����A�����bi�=�BD?0Ї?*�?��s?X�>�3
>dqz�����o辪�<R������Q½�">K��>�׫>o	�>���=ʵؽ��<�iF�|P�=}MO>�ڲ>�@�>eY�><<!>��<\F?̎�>_y����ʾ��¾C��˂�=ߜf?S(�?��H?-�:=ܣ�R3������?>/�?3ۨ?�6?�>��_�=M���fž�KN���>�V�>�˩>��:>1�<�:h=�đ>��>�� ��o
�l49��c轥Z?�/G?��
>��ſߺq�j�o�b��R�b<f쒾��d�|���S�Z��ǥ=jz�������@�[�qi���O�����A����{�ӱ�>��=���=PA�=?��<I�˼��<�bG=yے<1N=�q��0l<L)7���ʻ�7�����|R<OBG=����nʾ�}?.I?��(?*WC?��>(Y>� W����>��x�tL?b=W>m�;��긾Q9�\������پR�־�
d�oz���6>�M��>�4>Ϛ�=�(�<�u�=��n=���=�󲻏�<�$�='��=��=�P�=!a>g>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>%Q8>�>�R�?f1���[��*a���Z��!?:S;��;��>���=��޾m�ƾ��+=�P6>f�a=����\�6�=�T|�q�A=h�n=��>��B>�ֻ=�K��l�=y�H=���=9�O>G9��i�6�Dq/�^�8=��=h�a>7%>�S�>x�?޺4?Ěm?��>ET������b�����>F�\>9��>�>?��='C�>F�?n;?{D?��>��>���>�,�> ���]��e������>�4]?*�?�??���lr�����G^S��k��z&?��.?��?=��>�U����Y&���.�%����0.�W+=0mr��MU�����em���㽂�=lp�>w��>%�>KUy>��9>�N>s�>�>,9�<�p�=������<������=N���L�<�uż����.i&���+�򋦼��;L��;�]<���;�~�=h�>p�>��>��=p'��#�7>+����4L�o�={����A�w�c����g�/�<:��[C>[�Y>�����]��� ?��Z>�>>T�?xs?;q"> ����־o󞿄f���C�̾�=Ӗ>�(C���9��[���K�vվ,}�>Z�>�ו>�
g>g�,�� ;�R�~=�y���7����>;萾(�.�� ���s�j���ɟ��9h��E&��<?a���C�=��?[wI?�]�?���>�O���	߾��">͉�~�%=DA	���a�^ ��2�?p�)?���>a���G�n*̾�?��5ܷ>b�H���O�㽕��0�������ϙ�>&����о3��i����[�B���q�!�>��O?D�?�Ub��Y���WO���<���e?U�g?��>�-?�(?�i��>z��V�����=ʫn?&��?�9�? >��>g!�b��>]?4t�?�ky?v߁?}\\;)��>�d�g<�<���h�R=�v�<�Ƚ3{J�|�#?�$3?�n-?�Ƶ��M
�PV��s���нBXc=��ݻ�:�>�=�>��>��U=\U�;�*_=E�W>��>>8>���>��>��>Y���$��?.?�>��*>$��>gϷ>�"l>/`��?ؽ$��=��ؽ�EC�S�Y���3�PP^>�L�=G�w;�EK�̱f>�*��d��?N|�>��o��>�|�⩟=n�>�Y?��0=�@>�>Ԏ�>p��>S�>U��>�.�>�X?ECӾF�>��xb!��(C�2�R���Ѿ^dz>k���O�%����R���&I�Hf��4d��j�r-���;=�逽<"F�?���J�k��)����a�?�Y�>Y6?�݌������>{��>�э>�=������4Ǎ�[g�%�?Y��?�;c>��>8�W?:�?��1�r3��uZ��u�?(A��e�M�`�x፿ ����
�(	��
�_?�x?JyA?&Y�<�9z>9��?�%��ӏ�B*�>�/�';�B<=\+�>n*����`�z�Ӿ��þa7��HF>6�o?.%�?~Y?TV�� �� �E>�:?�t?ˢu?�=?O�-?�R����>�q�=�]?�o?��6?)�C?*�?�I�=Q��=j�$<;\=�����|��5�h���L��C:i�<�8�<e��jE=�%�=!�<��}p�����@	#��3�=��C=��=�yb=��>��V?���>��>a)?�'���%�����2?��=C�u�?e����G�����=�_o?�?�[?g�>��C��R�*Y>���>C�)>��C>�l�>�Ɩ��M��(.=���=��=%�=p\w�E���	��݂�<�7=��0>���>3|}>sz���$>^��z}v��c>3tO�#���[�X��tH��2��o}�I�>G\K?��?��=�(��0���e���'?��<?�XM?P�?�g�=�׾�;���K��V%�*��>�-=����:��|Ģ�5~7�8�<�Jl>�¤��P���v>��F�꾕v�A�����l=Ҕ��5.=�#�)߾������=K��=!��!���X�������J?��T=,����E��p����>�>嵱>6lo�fט�C�@�T����r=�.�>O67>�KǼZ���F��� ����>��J?z�K?,��?$�]�^>x�80󾺤��پn\>�8&?�y>�� ?%ͱ>#>F��6.3������_�|��>.F�>M��O=�v���k޽�g�/�Զ�=B��>y2>1?pZ?Bd�>�P?�-?ip�>n=D>�nн��,�a�+?�X�?�G�="�����u�8��\�㺮>e�?�6�����>�1?��-?;X'?��X?��>��=�Z��-����>��{>@.R��E��@��>�@1?�B=>�dI?�z?�.>A�3��sN��H��+��=�zu>k?'?5��>��>���>���>���z�����=68�?׉�?(L�?
E�>�j?Q��>uU�>�TE>>�9>3��>�3?
nu?[�\?j�]?$�4?�?�<�� ���%��ڌ��;�A/=!�>�N?=�]�º���,f���~�.5�|��{-Ͻ~�t�"� <�O=A��>`xw>z��Z�6>g�þJW��Z�B>����~����ۆ�ɥ5��s�=nڄ>�� ?q#�>�O$�/ؕ=���>{��>G����&?ڀ?4?$ܹ��c��Ҿ=H�W��>tfA?�#�=k��В�5Ks��;I=��l?�B`?[P�����Y�b?�]?`d�=���þ��b������O?��
?^�G�k�>~�~?Y�q?���>Z�e��6n�>��0Db�^�j�Զ=�n�>�X���d�tA�>��7?�L�>�b>f�=�p۾�w��l��@?y�?� �?E��?�*>��n��/࿊��z���k?�,�>˻�JC*?��ϼ�6����c�^l��?!��ԡ�ߩ��h�x������p��◾�Mým�=�2?t'|?=bR?_Bo?�~羡rV�̥M�Z���Ae����T��H��F�HU5�u1h�q\4�g�!���?�x<L�s�"AE���?��"?�I�t��>B_���Sɾ�����X'>� P�\k �T8�=��B�zrB<��=�v��K�����4r?��>:;�>�=D?F�V�x�3�Wa!���H����D>*��>�f>��>��=dP"���5��'���_���b�>��X?&K??0q^?�H��������8#�Tӓ��精{g�=��=��>����>����J+�EY�ݲd�s�羺���)���!>�=?��8>�t�>��?n6�>��
�򳾺���;���vz�>A�?��i?���>!+?K�q=l�A��> �l?���>}�>W����M!���{�8yʽ���>8^�>�M�>�o>�,�:\�+b������-9�,5�=Ȇh?󀄾��`�&�>�
R?T7�:%�Q<���>�u���!����a�'�+>ˇ?i��=��;>-Ož��}{�q6���U)?R?�G��hN+�@w>�K!?�,�>k٤>�m�?0��>��þ+f�:5?>�\?��I?�L@?4��>)=+���[���)�PL=},�>:X>g0k=׈�=�7���b���"�14=Q?�=%��<ȽHZ�;@ڼ�V<i��<*1>,ҿ�8���ﾌ�0�r��?���k���¼������]sо�`���h�������%==���r݀�\I�<�"����?{b�?���L�,��[����K�>�����=
���/��f�e�����
��U돾��ľ@/�PO�`�e�8���P�'?�����ǿ񰡿�:ܾ5! ?�A ?7�y?��7�"���8�� >C�<M-����뾬����οE�����^?���>��/��q��>᥂>�X>�Hq>����螾g1�<��?6�-?��>Ǝr�0�ɿa���_¤<���?/�@]nA?}|(��5�vJZ=�S�>=	?o@@>\1��P�Ĩ��&\�>5�?F؊?l\M=AsW����^e?[�<��F�����=%i�=��=���3�J>}��>_����A��ܽ�w4>�E�>@�!������^�Z��<��]>q<ս5�5Մ?,{\��f���/��T��U>��T?�*�>V:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�&���{���&V�}��=[��>b�>Â,������O��I��T��=7���ǿP�$�I�0��? =[Ҙ�mb����E'&�Z��_��
Hc��S�h��<@P>���>�6�>�ׂ>��>!_?o`}?�>�N�=V&:��D���>۾�s��;�����g����E����׾a�վ����Y����Ʋ�V>��u���[�]�f�,�4F=���?0�?՞���<A��S��W����o���7�"-b��!^�W}"�t�d���?&WF?���+�9��67��>�	�g�??���=�����ľ�>֓#����q�)>�ZL=����8:���8�V]=?w"%?w#����;�ߺ->�.p��2ϻd�?�Ql>��=P=�>&�=?�)�ַ!��>����>���>���<BP�����y?MBm?����[k��*?rT;�u���n����=�pоY�0��TS;z�V��:��+1>�P|��]�x(W?曍>��)����a�����S==�x?�?.�>�zk?��B?^Ԥ<Qg����S�z��ew=H�W?�)i?�>�����	о�����5?��e?��N>�ah�����.�<U��$?��n?�^?�y���v}�]��]���n6?��v?s^�xs�����I�V�g=�>�[�>���>��9��k�>�>?�#��G�� ���yY4�%Þ?��@���?��;<��T��=�;?l\�>�O��>ƾ�z������6�q=�"�>���ev����R,�e�8?ܠ�?���>�������g�=�z����?N_�?�����у=���;q�H
���ͽ��g>ĳ8���	��ɾN�s�ھ����v��U�<͘�>�A@����M�>K��޿�KǿL銿���p�ľ�a�>���>X㋾�����}�7���X?��X�:���?�>9�>{c��0����}�:�'m��^��>Uΰ�PF�>�U�u1��C-���R?<h��>���>d�>����վ���?֡���bο�,���]���X?ߑ�?�0�?��?�$&<@z�Нw���T��E?�r?^4Y?G��I`�6�%�j?�_��~U`��4�wHE��U>�"3?�B�>S�-��|=�>~��>�f>�#/�y�Ŀ�ٶ�7���Q��?܉�?�o���>s��?ws+?�i�8���[����*�A�+��<A?�2>����E�!�E0=�]Ғ���
?J~0?2{�g.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>eH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�L�>��?^7�=7R�>w��=�	���/�d\#>��=�m>�֐?D�M?�6�>���=�V8��/��9F�i6R�n ���C���>��a?��L?�a>���� .�� �#5ν��1���Y�@�t.��Bཟ�4>ѱ=>=z>�D�� Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?kQo���i�B>��?"������L��f?�
@u@a�^?*?+ٿ���T���ƾ>A5>:0�=Џ>Ui_�Ϲ����8֮<�A�/,=l��>=�$>?ne>�X0>�$h>�\>뒅���"����#9��D�e� �L���´��\m���b�2���{ҫ�ۉ.<Ɍ��z9�JF��^��d�3���=�^U?�>Q?;�q?�@�>?��};)>S���f��<���}�=ⶄ>e�0?$M?�=*?��o=���	fa�����A��T:��0��>��B>B"�>L�>�e�>��̻�I>��A>S��>`G>[�M=&�;��=�xK>&��>���>�`�>�i>��I>�i�������M|��Y1�?z�	v�?� �8�H��G���w��\6߾*(>=
� ?��=�W��*�˿㧿lC?�؝��|���ԽN�>N0+?5N?�t&>��Ѿ�vսcr>t���j�N�n=2V�o�w�=)�S�">��?'�>LG�>�Js���)��k�j�I�\@<�?� ��t���|���fE���)��<;��ц=.Fݽ/d�������􃿿�k�m�c��n]?��?�?>F�;�v�U�x�u�:��}b>�!]=ֹ�=S|>H�f�h�yQ����5:=��X=x�?�;4>��>	L�>�����j�抿>fD(>vE�=�|4?]�'?N�F�ʲ)�7�'4��d9>u1�>��>��m=ޑE���=4n�>L�[>�����+��тʽݠ��E�b>ZԷ�A�"��4���5�=�3�<�]>��M=�{ʽ�-ڽ�?=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>zx��Z�������u�w�#=P��>�8H?�V����O�i>��v
?�?�^�੤���ȿ5|v����>W�?���?h�m��A���@����>;��?�gY?woi>�g۾8`Z����>һ@?�R?�>�9�x�'���?�޶?֯�?��Z>s�?��\?mT�>�R���8��෿��~����=�l���z�=`��=�0񾔓k�7���뉿��?�4�h>��(=�^�> ����׾9>23Q=+�����;�&�>���>�9;p�>��?]�>��>)��=�U���R��/j���L?d�?P\�%�k�Q�=��R=��s��� ?O10?�;�˾��>
\?�+?��^?~C�> ��3��3Z��)��X�E<ʊ@>�+�>���>�8��af>�Fо�cT�f�>ō>I����$㾏
�����!�>�C?�!�>D�=l� ?��#?��j>�7�>@QE�":���F��t�>z�>�?��~?S�?����s3�^���꡿9�[�A]M>!�x?L?I�>%�������RFE��+J���V��?!�g?6.�x�?x�?�c??�`A?�af>�J��Kؾ�!����>."?G�	��$D��2'�����?��?�?�>E)s�ݽ5^�5]�����u?��Z?�D%?p���Ya��eþo��<;[�2���T<i�"���>�m>_J��@١=�#>A��=g�k��6�|><��=k]�>0�=^�8�+H��@,?�^F������= �r�_D�ѕ>�RL>� ����^?��=� �{�����{��XQU�@��?f��?SY�?���;�h�^=? �?.?�M�>|h����޾W��F�w��Vx�%p��(><��>]q�P#徘������[F��Oƽ=��;p��>��>�?�F�>��>�>=Ps�/J=�r��O���7j��Z�H�I���)��l#�О���P��I�y��¾,�~��,?���=��>&e�>��>$�4>��>iR>���>�S=�t�>��?��}>�m>d"N>�W�>�����KR?������'����4����2B?�qd?u0�>�i�܉�������?m��?s�?S>v>�~h�Y,+�nn?�=�>F���p
?zV:=�2�=�<AU�����0�������>nF׽� :��M�-of��i
?�/?����̾D;׽@H����=�h{?��-?w��$gS�Z�v��}\�;VO�����B�͹����.�ʙw��f���ǋ��[��<�7���7=��"?#��?��(	�Q~��o�q�j�N�;��>���>�=��
>BM$>���\�P�%�O��C�Mk��)[b>L�f?ߐ�>�FE?��??	�N?��5?w<>Q2?�z����>��>ԫ�>�?�T1?�UK?�m%?߲�>�<?:q�>���� �rN�3u?�w>�T?U^�>��>�o���x<�t�=��g�}��ԁ�䦶�4��o�j>w�����>)��>�N?N���8�����qk>,�7?'��>n�>>ҏ� �����<��>��
?n�>����{Rr�EO��m�>���?5���=�)>���=�1��C�Ӻ؊�=��r��=�낼.�;��3<i�=P�=)Ά��q*�G��:O��;!p�<zx�>��?	��>�v�>3���� ���Tl�=��X>xS>�>�_پ�z�������g�y>z�?�p�? �e=#��=ɶ�=So���8����������<�v?SP#?sfT?⑒?��=?�c#?E9>W�bH��V���ࢾȤ?<�.?y��>�s%��až�������3��>���>�`�f�W��2�X��a��/��YB�BBq�Z��W Y�N�򽒎��Fɽ�?�?�I�? �=ǡF�7���Ə��z��?�C?4h�>6��>ӡ�>L&�0�_�:���r�=x��>�/?Xs�>�Q?4
^?ύO?��Z>Y#T��Q��{���ʜ���>zs0?~?�Ȝ?�d?�W�>�!�=����签ݱ�d<}����o��C)�=__>�h	=!j�>*��>1(��.��B��u��qi�:6�K>w��>��c>$��>FQ�>�1�D�G?�W�>��ʾ� �x2��J{���P�Qet?�[�?E�(?S�<���H��$��7=�>�˦?�@�?p�%?�qV�p��=EM��6����}h���>2g�>�f�>ﮝ=�=0�>��>�>(���Z�a�6�i\�
�?�fB?��=Ѹʿ�y��p�����ɭ<����^Y��}Ͻ��a���=����^�#�����N�i����֕�ZQ���h���r�� �>���=4K�=��=[�<���r�<&�=C�=�7=�ʈ��;#;��C�ޣ&�Y���憒;��<s�^=�x���˾�u}?4/I?�+?��C?ҵy>��>�X.����>82��q ?U>�Q�G���J�;��Ψ��w����ؾ�׾d�2���C�>�D���>Z�2>b�=�2�<�m�=�rt=\�=�ŀ� �=���= ù=Nܫ=k��=�,>��>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?~�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��D����4�?��@��??�ዿТϿ6a/>t�:>�f>�FS��1��_�Z`���Z�M�!?@:���̾���>���=�cྫ�ǾM�*=��3>�Xi=���KH\�#��={����F=qS~=p]�>�zB>fz�=܃�� ��=|OD=�3�=�XM>�c���g>�c�5�~l-=j��=�pa>�g#>r�>�>?��0?�e?�>�샾f��9mʾ��>y6>�_�>UY�=a�v>S�>�65?��=?ËI?쏳>O[=�ݷ>An�>e(���c� ��rй�Gd =H]�?E��?���>���<#�(�m��	u5�'zԽ�?U
5?�v	?��>�M�%a����H�tA\���<�p>� �2@
=���(����"�U=,�>t��>�(�>��=v[�><��>6f�>�'>[	Ҽh�S=1mټ��X<��<Fld>��=�M;=�����@��(+=� /�jw�M�=4?>�#>'@>8��=?�>g�>�>�	�=c ��0>g���M��$�=����A�H�c�>M~���.�1�7��TD>r�U>=6���ᑿ/-?��\>�C>��?Ӧt?r">��\^־���g�d�4�W�x�=�>b�?���:�1�^���M�T�Ҿ���>g�>員>�k>n*�;�<��D=��޾�4�=��>o{���G�@�Wjr�kͤ��5���j�6JO�҅@?%p��N��=e�?�/H?W�?�K�>�����Ӿ�31>R|r��F=�_��)Z�t�f��?�'?���>Z���@��̾����׷>r-I���O�b���έ0����u᷾r��>���Ѿ�3��d������|B�G�r�iͺ>�|O?�ծ?�b��(���JO�t��tv��z?,�g?�P�>�I?�i?p!��E����I͸=��n?Ҝ�?2C�?��>��<�����>.��>6ͧ?�ԙ?��?S�T�.��>�>>@֑>�Xp> �G>��>���>)n�>D�?�<?VdI?p�ս�i!������{��ՖM>�F�=O�>,~>r�4==�=T�9�}@;�/>���>m�>�=
"X>+Ŋ>|$}�Xk��n=? ʃ=�F2>��?�i�=[��>�8ۼđn=��>ꐽ�y�����W��3K�>�7���<��C;�G�>�G���X�?�d>��P�?+����=e��>&*>���>�K?��>_�>U��>�	?�>�=��>��>DӾ�>���d!�w,C�˂R�пѾ3~z>j����	&�A��p����EI��p���h�<j�.��0==����<G�?����ҽk�G�)�-���]�?�]�>\6?،�3���>���>Yˍ>MF�������ƍ��f�4�?���?)Tc>��>m�W?_�?}1��)3�VZ�V�u�4,A���d���`��⍿{�����
��	����_?<�x?oA?7��<2"z>A��?��%�}���]�>�$/�;���9=;A�>鰾w�`�ۙӾקþ��w]F>�o?��?�c?MJV���n��>��<?i�/?�q?��1?]�8?k+�� %?w0>�
?G?��5?��-?ߪ?8�A>2��=�Ա��&>=����6�ǽ������`�R=G��=�n5��<NU�<;�<n��ۼg6�;%Q��D�<�<=�3�=���=\ҧ>]?��>2,�>�6?�����4��߭�P,?�<=㜀��R�����B�G�>�Kg?��?iY?��Z>;�A���?��E>:m�>i">�V>J��>�4���>���=12>�>k@�=����^~�FU	����Q��<� >��>�;>������>����wh��]>��H����FSa�P�G���2��J����>�)F?��?�/�=��M����c��!%?��=?��N?;�?�ف=�ܾ�z7���O�z����>4��<���y���0f����8�������f>������Yr>RZ��龇�v��\L��}�MR�=�T �#+B='���ξ1L���O�=��>����������p��hJ?=GN=�G��P�T��F����'>�c�>���>#�K�O�<�FK�����e�<g��>�~0>�"��M龗�Q�f$��R�>:�D?�^?���?����q�P?�i���!�����?>�>�?�TE>�ݳ=���E���eb��sF�l��>�|�>��YxH��ٟ��7��b&$�'�>#�?%�%>��?G�Q?��?��_?�'?�%?��>L���*���-B&?���?ẅ́=]�Խ��T���8�F�,��>�v)??�B��ė>C�?ڳ?��&?uQ?T�?/�>�� ��;@�̓�> Y�>��W�d[���_>�J?R��>�*Y?5ʃ?e!>>��5�Wɢ�����_p�=�%>	�2?;#?ա?є�>쬹>��¾���=���>�ky?r�u?��}?��z>z7?5�w>��>�D=�4�>�� ?g~%?=V?/�s?��O?ɖ?*=X<f#,���"���f ��;[#����-:>��5�ek��v����o��u��~��<�͞�${=y}���$=�=%��>[�s>�唾J�2>v�þ�#����A>Է��.b���Ҋ�H�9�/
�=ˁ>F?+k�>�Q�<�=��>���>�Q���'?��??���6kqb�vZھ�	F��?�>�@?���=Tlm����hv��ya=�^m?�]?z<V�N�����b?��]?�5���<��PþACb�/��%lO?��
?Y`G��:�>S$?��q?���>NHg���m��휿ޭa�j��7�=�u�>�\�ԑd��]�>Y�7?q��>�"b>v�=�۾�w�^B��q�?�Ռ? ��?�̊?��+>�xn�>�t����&����]?MM�>ტ��"?͈c�e�ľ[�n��f�ݾ����l+��ϐ��m�����ᆾ�dɽtr�= �?�#r?�Jo?�6\?S'���b�w�^�v�z���V��7�����EF�·F�Y�D��so��m��:������B=�@^��v3�9N�?��)?^�Ͻ�D�>�ih������?���m>>u�L��m���5S=��<�ș=�m>�]n��Z\��0��>?���>'c�>(�+?-S;��G���G��)����>h��>�^e>��>�|*�����������־-0e��m!��%w>rhc?w�J?݃m?����%E/������"�	�/��L���MC>>�!�>X�T����B&�|�=�^�q�6!�����u	�6�=�2?]�~>��>�S�?�?�&�������y�O�1���g<Ʒ�>Tri?S��>���>�%ӽ�U!���>˿k?w��>L�>R���2�+�{��n�A�>�:�>/�?���>@&��![�È��҉�t�6��>F]d?�s�N?K��f>B)J?m��<�#=��>�D��P� �o���j>���A>��?�:�=��]>�$��";����p�S4��0�%?i�?�ً��[%��̓>�e#?���>�<�>SO�?�7�>$L����� $?P`?�cJ?� C?�U�>� 5=	̪�����}�$���;=gq�>�J>��E=ח�=n�콫�b���*�F�3=p��=�+ �T�׽���;[
Z����;y!=��->SIο�=9�#��
��i��z7��X@`�w����2��f��b��!��l�o������-Mݽl�l��!��@�"����?9��?��Ѿμ�v0��dm���1+��l�>⯂��A��+Z�3
��ރ�ݕ便VF�2��[X��cn��7��P�'?�����ǿ񰡿�:ܾ1! ?�A ?6�y?��7�"���8�� >9C�<`-����뾬����οC�����^?���>��/��o��>ޥ�>�X>�Hq>����螾�1�<��?8�-?��>ǎr�1�ɿb����¤<���?0�@�A?)�&����P=���>�	?��;>�23���Cӯ����>���?�T�?M�@=�W����>(d?&8A<��E�9�Ż���=Ө�=B'=1���K>%b�>
;�p�B���ܽ'0>8ć>$?!�G��8�V�]��<�mc>�׽!���5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=k6����{���&V�{��=Z��>b�>,������O��I��U��={ ��Ŀhp'�[�,���><�%>=�H�����߸��ҽ�,��+�U�N\ؽx{=���=x�m>���>��>z{�>�d?!�~?�r�>!Z>�J,����w��u���?����<�m3�b���T��
�ξ7Z���%����J������M==>�3v�d펿��M�6x���K��=:?٭�>�[ԾqE+��NT=���씭�bf�=5�"=�'ž���<�h�᧤?�@?O���h�I��V.�/]�v o��]G?�?M�q���i��Ì=@�(A�<�-�>��;�ꪾ~oh��_��,2?��&?�{��!0��d,'>�--�� >��?��>�6��B��>�aK?R��O�o��V>>h=�M�>z��>-IŽ�艾i9���?)Dr?C���4���?�ǽ�ؔ��5w�ǻL=[���H��۝c>�&p>;�����=#픽>�(�W?��>!K)�L���󎾢���&=,�v?�,?x�>��k?�{C?�z�<�J��G�T���
�'�i=0�W?߼h?��	>�wz�?Ѿ ����5?�e?S>8Nj�s��QB-���U�?��m?��?�p�Q%|���������s4?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?o�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������[��=-������?�>�?&jO�7��WD�Q�N�����:�=%d�=߂� 5�!|���,����}��i���dT�7ي>#�
@>�}���>�X���Jҿ)�п�����t�^�YB�>m��>UxP�Baþ� |�����`�?�BS������>I�>����矒�UB|�Ȳ;�謁��>�m��׺�>cT�����Cr���-<�\�>���>�v�>~��d�����?���� ο񅞿R����X?��?jH�?\_?�O<m�z��|��X4���F?ISs?��Y?ʼ"�ri`�ϋ<�%�j?�_��wU`���4�tHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>q��?ts+?�i�8���[����*��+��<A?�2>���I�!�B0=�SҒ�¼
?W~0?{�f.�]�_?*�a�M�p���-���ƽ�ۡ>�0�f\�N�����Xe����@y����?N^�?i�?׵�� #�g6%?�>d����8Ǿ��<���>�(�>*N>bH_���u>����:�
i	>���?�~�?Qj?���� ����U>	�}?�2�>P�?eb�=j�>h�=�ܰ���*��T#>Ѽ�=:�?�#�?e�M?�%�>)�=��8��/��FF��,R��"�7�C�?�>;�a?J�L?-b>2���0�i� �C�ͽ�`1�����A@��i,��&߽qS5>G�=>U>I�D��Ӿ��?6p�,�ؿ�i��p'��54?��>�?��|�t�����;_?Fz�>�6�,���%���B�\��?�G�?;�?��׾3T̼�>C�>�I�>��Խ����e�����7>�B?���D��`�o���>���?�@�ծ?ji��	?���P��Ta~����7�M��=��7?�0��z>���>��=�nv�ݻ��Y�s����>�B�?�{�?��> �l?��o�P�B���1=9M�>Μk?�s?�Ro���l�B>��?������L��f?
�
@~u@_�^?*ɳ㿍��^�þ�N��;ļDd >*z>1:=�V�>'��;����
�=��`>}2�>�+�>{�>Nݟ>U�H>o��>)���� �w����͚��	J��b�������G&�1a��ھ&�)��۾F1�<�T���;��@�^����>��Q?:JQ?�ar?���>Һ@���I>�s�37F�x�*�'!�=Zp>�-?�O?�+,?W`T=)w��zAX���~��ܤ�t|����>��>OH�>���>c��>�<��>>�G^>��>�� >	��=�`�<!��<�D`>���>��>�$�>4k�>�zM>��ſh>�����J*y������F�?w�>���=����=�j�xI�;�EP?�m"�%��w�ѿ%��Z�)?����ܾ&����>"�?^� ?�`	=�Y/�ڤ�v�=@�t�����V�l����B����E�5EX����>�ކ>.8t>�)A��);��T������3>%�4?Ӿ��j��<h:�g���!`�=M�>2F���*�����j���c��d�=��B?�?j��
ž�F]����;�K>0�f>˯�=d�=|qA>�,o�90�oP���ڼ���=w&N>��?]#3>��>l��>fĜ�vp5�7i�>�LI>W�=D
 ?�6#?@����z,/��R����C>���>A��>� ]=�?B�)f�=�C�>ߤ>�K���!}�O$2���/>NA7=��"����L>�V�<��=;"�=�0�Lz�I=�~?���(䈿��e���lD?S+?\ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��J��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿrh�>�w�fZ��}��o�u���#=���>�8H?IV����O�N>��v
?�?_�멤���ȿ-|v����>A�?���?&�m��A���@����>"��?gY?�ni>�g۾u_Z�\��>�@?�R?��>�9�p�'���?�޶?���?bl:>�5�?��W?���>�V�=�_�쇲�������<�qN>e̺>M�>riX���	��Vu��JQ�K辨	�>�bq=��>��-�\ 
����=}T>�p�1~z�0�>�d�>�6�>�u�=�R?�x?3Y�>�Ȏ���Ľ�����Z�}�K?���?'���2n�[O�<���=3�^��&?�I4?�j[�o�Ͼ�ը>�\?f?�[?d�>9��F>��=迿*~��w��<k�K>24�>�H�>�$���FK>��Ծ�4D�6p�>�ϗ>����?ھ�,���O��IB�>�e!?���>7Ү=�� ?�$%?�_>���>:�4�Ao���P�:s�>��>$[�>�Q�?"�	?�r��^�6�~��x��%-^�d}h>A�v?�?���>�ŏ�$)���W���Tμi���dX?"�Y?5uB�v��>�p�?�S(?ʯ&?..>o�#����Iΐ��{w>�f!?����[@��n%�>���?o\?�k�>�G��ս |ۼ�r��"��>�?�[?Fj&?`�'a��Bþ�G�<Z�+�xn�W�<EsH��>��>�U��FѸ=��>�{�=�n�v�3�k
�<�o�=O�>���=�"7�Ϗ�0=,?5�G�yۃ��=��r�9xD���>�IL>����^?al=�	�{�����x��	U�� �?���?Xk�?���;�h��$=?�?V	?d"�>�J���}޾4���Pw�~x��w�N�>���>ۡl���I���֙���F��F�Ž�M��n�>L��>��?���>�:B>ʹ�>�I���L4�Z2���x㾐7�:�-����"��U�:�W���2�1����/��/N���?�>������>A�?\�>���>��>N�,=�V;>��>X��>���>�%�>�+�>j�=>�FP��]ڽ�JR?R���e�'����ޮ��Z4B?�od?],�>�i��������}?���?'s�?�>v>3~h��,+��m?�=�>���Dp
?iZ:=8��-�<fS��|���&������>jF׽�:��M��lf��j
?b0?Z&��,�̾�B׽cv��%�={.z?g�)?�T��\/R�<Aq��RC�\�K�]�B�*��q%���O��P�k3���Ձ��7x��A� �>�I"?�3�?\!�)��N%���N�ϜY��4Ǽ���>3ـ>�?�>��>���nA���o��9B�J���2�>
?�R�>��:?��C?��O?�| ?b��>:[
?��}��x�>Q��=ώ�>�U�>H>6?9s>?�3?W!�>�O?Cǚ>y��8\��ƾ�u�>���>Ի:?6�?1[�>Y�#����=�>%o��~��,=<�8��^=$o�;d�<]�>_'�>�?�S���6������0n>��5?���>ϑ�>����E}���=X��>'	?`��>�I�^�o�}7����>�-�?���x�=v&!>�S�=8�:�N�];��=kGм��=���$.`��_�<Tr�=Є�=cxY<���>5�<��`:��;�t�>�?�>�E�><��.� ���>t�=HY>��R>�,>�Jپ~z��"����g�@Ty>@q�?�w�?�f=u3�=$��=�����Z��\������j(�<��?NG#?�UT?#��?�=?c#?5�>.��K��[Z�����߮?�:/?Hё>:I��U��LI��}�\��>���>J"c����7�#���z엾|p��GG���N�@���<h�K��@	��r��}��?�9�?pT_=�;<��͌�f9�������q?�I"?0�l>���>�����#��������>8]=?��{?��>�*O?�He?`	$?Tt�>�yA��ϟ�����k�=�!�>=�5?��?�~�?$��?f�>���R���;�þ��^H�^��9�A�~��=X�0>��>��?���>��u>K���ҽ.��ڄ>zi�>��	?P�?�S�>�4>�\��r�G?��>Z�����r줾�Ã�w�<�+�u?���?�+?We=����E��B���H�>m�?P��?3*?��S���={�ּo඾��q�#�>�ڹ>	0�>ē=n^F=�e>A�>
��>G)�i_�]o8�3^M�k�?�F?o��=��ſ��q�>Zo�~���ug<E����wd�������Z�ť=K���(������0[�́������Ǣ����/|�k��>���=X��=�c�=���<�μM��<X�I=s�<�=fom�զd<:X5�6
������т�AY<w�I=2���Kž��{?$�G?��.?�t@?��{>b)>Ĩ�6?�>�R���?��S>DY��ǣ��F�/�k�������>�Ѿ.۾��`�{J��D�>{�4.>��->�-�=��-<���=��=ރ�=������4=�7�=b?�=@X�=�Q�=�u>��>�6w?X�������4Q��Z罥�:?�8�>f{�=��ƾq@?}�>>�2������xb��-?���?�T�?=�?Ati��d�>M���㎽�q�=K����=2>p��=v�2�U��>��J>���K��@����4�?��@��??�ዿТϿ4a/>�3@>1�>mkQ�C5.��]���^�h%X�h- ?ŋ;��ҾDs�>�F�=���ĳʾ��=C5.>.tL=��7i\�%��=�(u�e^P=�1�=5�>8M?>w��=�����=�wP=[��=!P>�����b[�Z9=`��=�^>�M >���>��
?�o-?��]?�R�>���9��o�����>���=B�>�P=`\�>l��>�C;?��L?�\:?��>F��=�2�>;D�>�Q!�*�L����Gþ���=2��?��m?��>݈��	~��l�'��@�����?�.?�?���>�������8)��=e��#�nl)�cR>Ҕ��>��>k��BQ�=Q��=⪖>5,�>���>3��>��>�V�>G�>�r>����{�=�����WS=Y�{���%<~��ਸ਼=���<8u��;읽&^!��Ռ���⼔�9<�=�L5=���=N��>Le>���>,��=Y���?/>{����L���=�B���B�T;d�wC~�i/��h6�'�B>�X>M����/����?�Z>�H?>ɀ�? Qu?c >����վSM��Sxe��CS��Ҹ=�	>�<��^;�'B`��M��}Ҿ��>�@l>$Ʋ>ی>��Έd��̔<l� � 	]�&�>���-G�;W����z�6!�����	�V��]��&�3?�~�}������?Fq+??l?5ɤ=�S����>����3+�q�Ͼ�ă�L�#>К?ɫ?��0?�'׾*B �4̾@پ��ٷ>>=I���O�������0�ha��·�"��>4٪���оq3�Wg��f ����B��gr����>S�O?*�?�(b�tV��}TO�}��q���ol?rig?�>L?)8?\���fx�er���[�=?�n?���?r9�?��
>xP�=�%�����>L
?��?�s�?��p?Gf�I��>� �=���=9�Ƚ�b>Cg>��z>*>�?�!?EV	?�8ҽCZ�u����Ⱦ��̼ڰ�;c�=�<�>���>}�>�n�l�S=��=���=ٳ�>�0�>��->���>]a�>难�C��1?Ԩ >h�>�.?2�>ʢ>=��ǽ�@=C
���k���i�u!��JM �c�=�<�Ҽ|U3�3��>񔿿�S�?�I>v���'?��޾:���J�>�u>��Ž`��>e>�O�>Pm�>W��>ė>	oh>5g�=��Ҿt�>
��!�Q�B�dxR��Ҿ�Nz>�����0&�jF������H��U��)���i�'��=���<i4�?ż���k�*������J?�N�>8w5?Er�������>���>�s�>I���p���=΍�9�T��?���?�;c>��>7�W?��?��1�23��tZ�n�u�(A�	e��`��፿}����
� ����_?��x?�xA?�J�<�:z>
��?1�%��ӏ�T(�>�/�<';��?<=8*�>�)���`��Ӿ0�þ�8��DF>?�o?�$�?�X?�RV� Ci�D#>q�:?�1?Тs?�1?��;?ct���#?�2>�I?�
?*64?��.?T?��5>� �=o���Q$=���|��CϽ@�ɽ�2���&=>�{=nx�;��<p�&=��<6y�t���m��;�n��؂�<"UA=*!�=�g�=X]�>c*]?U�>	
�>~�6?g��v<6�gᬾwy-?��=�D��)k���j��FQ�#�>}^i?���?eZ?�_>A�,�B�~k>�9�>�.$>�[>��>v�JGG�R7�=o�>'>�+�=ڄ=�܀��s	�WP�����<~�>���>��{>ߒw�o�0>9����>p�Nf>�bA��
���X�"CE��7���i�^T�>&sK?�?�Ӈ=-侕
���lb���(?
^;?kuJ?�/{?��=}�޾5�5��!K���$�i�>�S#<i����(�����:�&�-�+�m>���3��ȶ�>]U�M6�i���6@��:��=оs��<'������*����=��">����m"����C���q�K?��m=����[�\��B����1>D�>�B�>g�1��z�;a�P���Ͼ	�V=���>�0>�w���=E�I��L�T>��;?q�R?��}?��ú~�O�/�a��a����>��G�*?v�>(F$?�T�>�'>5��������D��YC���?��?����l��썾��ɾ:E��ǒ>-?�4�=�;?��J?��?�=E?�6
?�>;�(>�J�kL��;n+?���?��.=�_�?R���27��tG�반>E?�e���Ǽ>�)%?n�H?�H?��C?�*?�==p����'���>tr�>Ok[�Z�0�d>��V?��E>��
?�p?6d�>Y_0�$���i!D��U<c��=}�>1�?�-?߇�>�p�>�ܼ���=k�>�c?���?)w?�K9>��?��@>c�>Qr�=q5�>�$�>�(?:�R?�v?C�S?z�?V�<�G住����E���(�տ�<8/K�_�{=��`�ѽ5�y�l�<#ԃ��bѼ��N<�(���e�V�ڶZ<a�>�r>�,����;>�þ/ꈾ��G>&ᄼ27��9���G�:�sy�=�"z>���>�)�>�w+����=N��>ݾ>cK�ei%?��?g?��;�ya��z;s~F�'~�>��>?1��=�m��蒿��r�/=yo?^?�%S�~��<�b?�]?�g��=�4�þ)�b� ����O?��
?K�G���>��~?��q?��>J�e��9n�����Cb���j��Ҷ=r�>NX���d�9?�>��7?�M�>y�b>�&�=�t۾��w��q��&?1�?��?���?"+*>D�n��3��#���Z��C.b?ƛ�>Cc��l?K�;�p�Ⱦ/���A����Ͼ���︾	)x�牟��1*��|k��b�|�=�?��v?�f?̘_?i/�mPa��[��\����W��U� ��cA��D�~1I�'�_�+���+������j�<MN����R��?�*:?�7��vju>�a)��eξx�ؾP:}>Z���ܛ;9��=CB^>��)=s��=��������$�	?��>2�>�;?	j.���9���'���&��=�Jv>]�>>���=@%�-��=�D�4��1{��~�����n>5�_?��H?��d?"Ľ��#�8���"�[lT�66��R�,>��;>g��>�3��7��!�Ke7�Z1k����c嚾�D
����=��0?pt>P�>}�?(�?T��=��BZ��#��p"=6"�> �k?z��>DҞ>\|��Hz)���?��]?T��>S7^>j-]��:
��f�d�\�q�>�8?��{>��V>�����U��}��c�����8>C�Y?T�d�ֳ��|��>z$c?�IF�⨨���>J�9>j%��.�����<�>�4�><���U�=p谾/ٻ�(녿������,?�?�d���>-��7O>/ ?���>�f�>���?''�>A7־Q�i��n?1�X?��I?v8??���>��=8�Ľ�Oý(�/��=�T�>ys>�ݠ=u:�=8����x����'$=j��=%7��	��;~�K� #�<�Y�<Bd%>s�쿬BT���%,�՛ؾ���5cJ��o��kQ�S�i�7Ҿ�پX�D,K��V�<1�b�T���q$��������?�+@i����q�y���Ί�6\6��_3>�*��������^Խ������}�X�N�
bR��8O��b���)?%�z�J:Ŀ;5��s�ɾ��?�}?�]j?�
�z���/�o1>��<��ݾ����A�̿r@����Z?�Y�>�#�?�����>I�t>��b>ڥy>𘐾�����4=�
�>�%?���>Y~�%�ǿQM���5�<1s�?�9@��A?��'��s�[�F=���>�	?��;>�2��G��v���>�>Ş?U)�?��7=�:W�,��� d?��<؇F���	���=���=%�=�m��F>���>O@��D�u#ܽ.�1>��>S�.��(��*c����<y]>CQٽ�n���Մ?}v\��f�Y�/�-V��*]>�T?{-�>�\�=��,?2;H�XϿ�\�&a?&/�?���?~�(?.ۿ�ZӚ>��ܾ��M?�C6?���>
\&���t�]~�=n%἖⧻*��]"V�D�=��>�l>�,�����O�2������=��Aȿ�"���X=܄<:�4��ؽ����Jl�H���A9q�Z�r�s=`W�=(Z>]��>�RS>�h]>d	[?w�p?�l�>�>76���Ǌ���Ѿ��̼W��L$������ �M���b��۾�	������оa�*���F>��f�H#��w�>��{i�e�V�ێ?�E�>�*�D�!��2<��Ͼ����C�>nc�<*S˾e� ���B�K��?"�7?�ĉ��+��0�K=^;��4H?�;�=,5�`{�Ĳ{<�:��]'�=�V�>�U�=}���)��5���9?U�$?�z��`؝��G>͉ٽ|{���?���>g�>Q�>�r?�<����<�a>w��< 4�>���>�{>�����0��Q?�U?$'�]u���H�>�����.����G=1��=��U�M""��>9����黾2�7<��i��H/=��W?_�>^})����\����%&=~{r?��?�B�>'j?�A?C �<�v��P�����W=�MY?��g?�E>?%����ξ@ߢ��B2?WEd?$�Q>n/j���`�+��U���?3,g?��?�G������6�����g�6?U�v?vs^�Os������V��>�>�\�>���>`�9�l�>�>?C#��G��κ��+Y4�AÞ?��@x��?�#<<, �嚎=I;?'\�>�O�0?ƾKy�����^�q=�"�>����ev�����Q,�ׇ8?���?M��>������ �=`�����?� �?�䚾�*�W��b��[�}�<�d�=$*<U����x¾v%�6;Ҿo�	���������n�>)�@�B����>Ȉ<��;׿a�ſ>p����̾('��EN�>���>8 o�+�о
�c�־|��[i��66�,mL�t�>9�3>��x���yꄿ>5�`]���Z�>l�=\�K>�L�a��������P��>��>Z�c>����L��z��?q��Z�˿������Z?ڊ�?0Ԁ?<�?���=�L��HƟ�����lyA?�yW?DzV?�悽0�r��D��b�j?	���'�_�Pt4�:ID�1.U>Z02?�Q�>�f-�x�=��>���>�/>/��)Ŀ�Q�����Ӧ?�?/���q�>1�?�+?�.�����DR����(�
��h�??+>$���U"��1=�M哾Y�	?��0?�I���^�_?�a�U�p���-��ƽ�ۡ>�0��e\��K��"���Xe����@y����?I^�?g�?��� #�a6%?&�>_����8Ǿp�<���>�(�>*N>NH_���u>����:��h	>���?�~�?Gj?���������U>��}?(*�>��?�c�=�]�>�.�=�����-��o#>���=sj?�ߛ?=�M?(:�>��=e9�:/�WF�BKR�X)���C�C�>>�a?P�L?�<b>*���1�{!�w`ͽ-x1����8o@�M�,��8߽�5>��=>}>8�D��Ӿ��?Mp�9�ؿ j��p'��54?/��>�?����t�����;_?Oz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�>:�>�I�>A�Խ����\�����7>0�B?Y��D��u�o�w�>���?
�@�ծ?ii��	?���P��Sa~����7�x��=��7?�0�#�z>���>��=�nv�ݻ��U�s����>�B�?�{�?��>�l?��o�O�B�{�1=;M�>͜k?�s?Po���k�B>��?#������L��f?
�
@~u@`�^?(�hֿ����MN��F�����=���=ֆ2>�ٽ6_�=�7=R�8��<����=��>��d>$q>F(O>ya;>��)>���N�!�r��W���Q�C�������Z�E���Wv�Vz��3�������?���3ýy���Q�2&�R?`��w�=�RU?F�Q?��o?~ ?��s��) >�u����<
$���=��>ص2?�\L?�)?�m�=(ț��d�c0���+��3��4�>��I>A��>��>7X�>j�A;�H>N�?>d>oo>��-=���=�P>�R�>���>T�>���>D�b>П��8O��Z%��r�H�K����?TҒ�t�7�~��A��I�Ͼ�N=_,?�!;>:���]������^<?���=h������A>G�3?��N?	G >@�Ͼ�I���s+=U���`�@V=B����h���>�U�>y+�>�,s>��@���7�{IC��;���=#L0?��Ӿ�����{�ۇ+�8 ⾭����y`>%�"<42�P^������y���D�=�Y?�4?kV������S��c��BY�<��'>��>R�=R!E>�J���{���(��[<E�V�2X�=��?��I>�>g�?s(���Li�b[�>�J>�6�=��-?v�#?��,�}������S>�G?>o��=᠇�1��=�A�>�,8>_���|���m���L�[�K>5��=F�8���=FWG>r�N�N�5>T�'>feʼՐ�����=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿsh�>x�{Z�����y�u�5�#=&��>�8H?�V���O�G>��v
?�?�^�Ω����ȿ-|v���>H�?���?i�m�}A���@�J��>'��?�gY?doi>�g۾`Z�J��>��@?�R?��>�9�M�'���?�޶?ѯ�?,�=�D�?��^?[�>�Y>���`����D���n�<5�F=�G">	Ԝ=_ŉ��;�jA��t����~����z��>�ٻ��>$��Ⱥ
����=�N�=3�þ���)��>q�f>��)>��>��>?�d�>�)+>.�>�eI<�m��U"r�(�L?���?�����o��(=4��=��j����>�m1?�B<��ǾF��>�x]?�b~?�{Z?�Ð>��f���＿*İ��er<�c:>��>l*�>D
F�E�M>�8޾h}F���>�a�>������#̓��Ǩ��>�n?�	�>��=�� ?4�#?��j>.$�>�]E��8����E�,��>���>�K?��~?��?5Թ�?Y3�n���硿��[��BN>A�x?HU?�ƕ>���5���N�E��@I��������?lrg?�V�@?�0�?��??��A?^f>���(ؾN�����>�%?�?⽖4K���)���H��F?��>��>�����Ž�J���Q(��l��)\
?�Y?r�&?� ���\�(Aľ�O={K����0T;<�*<t�,>G$>��v�+�s=��$>D6j=�����5���D��2�=˟�>R��=X>�"����=,?j�G�k߃�2�=��r�vD�:�>VKL>� ��|�^?�s=��{�[���x���U� �?ҟ�?\j�?�����h��"=?�?�?�%�>�H���}޾p��GYw�s�x�?v�h�>d��>n(m��徯�����F���ƽ�����>f�>,� ?D�>�+�=�
�>�K�}�/������'p^�ej#��.�
*�J���f��2Z��r���y%��T��>�@�=)&�>0��>a��>�F>RR�>��C�t��>�N�=���>FG�>l)y>���>�p\>��Z=�6�	LR?������'�*�辙����2B?�pd?}/�>Ki�l������3�?��?�r�?�<v>Dh�Q,+�|n?�=�>{��fp
?�V:=��T2�<YU������0����Y��>�C׽� :��M��nf� j
?�.?�����̾�;׽�%��p��=e;�?�{:?���R��d�y�`�� T��;�6�V����z&��W�)����p���܊��3�ʡ =��?���?������|�&�h�R�,
:�￺���>���>��y>���=Nľ�l1��9f��60�����}�>�k�?�4>�;0?�:?ѿP?��;?,=~>o��>a����>�S�<���>��?��T?�%?.\.?��?�B?mZ�>,x5��h�a_�U�>��
?Sp�>0�>�
.?f2��@0%�М�=\���|�<�� �����b~>�r���:�<�ht>uՃ>i}?����8��1����q>A7?��>È�>�����h�9S�<���>U�?��>~���Itu����Ay�>.��?��5��<H�'>}�=F�Ѽt��)Y�=�X��Ū�=�?e�M�|��@
<qC�=�W=坼yO�� ><�;���<x�>��?>�A�>�;��� �L��'E�=Y>�/S>�>Eپ4}��6#��L�g��Ey>v�?yz�?��f=��=͂�=.z���O����������<��?�G#?>VT?���?a�=?�e#?ܫ>�+�xM���[�����^�?��+?>��>���ʾw~���^*��&�>� ?m<s������%�Ϥ�a��CH����I���Y������f��J=��3�������?�͗?;#ؽ�K�3���A���%��?D"?p� ?ag>�{�>�yӾ�q�}o��]>6�>��,?��>n[Q?K8s?t�>?Z�>��O���W}��M�����=[0?@��?�?��}?�f>��6>[�b�1�����8Խ�-���N�-B<M�L>Pٌ>x/ ?�� ?p�=���-���U+���]C>Iqx>&�>���>.�?�Z�>L1�\�H?�1�>�ž�U��4�����2�E���t?Y��?q�*?x�<��ǣE�p����>"v�?;1�?F�(?�U�V��=�����h���1p�� �>�d�>l#�>��=5�=��>P"�>���>l3�;��}8�4�c��e?��C?J#�=�ſ�s�!�`�2N��I H<v+���b�ϧ����S����=t!��zZ�	����C�rܨ�ԧ�����򦜾��s�0P�>�Sy=���=ƒ�=���<k��U��<�O5=��;ʧ0=�L��π�<@�l�ܫܻ�dp�mͻqB�<��^=LLu��o˾��}?/9I?��+?f�C?A�y>au>�}3�R��>W���NB?�U>�"Q�����s;�<��������ؾws׾,d�`����L>\I� �>[13>z}�=�<�5�=��s=?؎=;I�)�=�9�=kg�=ӭ�=�8�=��>�]>�6w?U�������4Q��Z罣�:?�8�>s{�=y�ƾm@?k�>>�2������xb��-?���?�T�?<�??ti��d�>J���㎽�q�=S����=2>���=s�2�Q��>��J>���K��K����4�?��@��??�ዿ΢Ͽ*a/><�8>��>��R�y�1�ME\��b�$/[�\b!?�-;��!̾T҅>���=��޾��ƾ�--=�<6>i�_=��P\����=��{�kE?=�m=�݉>lwC>ؕ�=����ɴ=��J=�8�=rO>8�����7��|/���.=�-�=�b>�%>J��>�A?�f0?,�c?���>��o�-UȾ�⽾5��>��=�D�>�"�=��F>+�>�8?n�D?��M?�ǵ>�R�=$з>~��>�,�4�n���a\��1(�<G<�?�G�?Tw�>�L,<d�B��h�`�=��MȽ�T?�<1?�e?a�>�U����-Y&���.����Ý5��+=�mr��QU�����@m������=�p�>���>��>JTy>#�9>��N>{�>��>�6�<�p�=㌻	��<� ��r��=ꞑ���<Ovż����Q~&�t�+�l���D�;���;d�]<r��;��=)�>�>6��>i��=�}��j�*>���Q�K��@�=����
�A�/�c�-h�HS.���6���?>��Q>"���q鑿�#?�ec>gA>9��?�s?;�>P����پ�M��D~]�x�F�0�=Vg>X�B�ε9�L�^��M��fӾK8�>���>���>�|�>'�*�"�6���5=?�s7��I�>O�������'j�j�����qm��CON�N!q�NO"?�����5=,ǃ?�Z?+�y?���>(�=�r����=>?��,7>���4E��q�<��?�1?�{�>lu̾C9�D̾��Nܷ>�AI��O�����ٯ0�	��i̷���>����о�$3�Zg�������B�Kr�!��>5�O?��?#:b�xV���QO����1��
q?�}g?��>hG?`??P$���y��r��Zy�=��n?��?S;�?��
>I�˽�X�����>Kp>��?p7�?3N�?T�>�B�>#	�>(]L>��� ҟ=�*�=��>��>i�[?`?,΁?w���"�N�����1���<> �=��>+��>X��=x��=Ib�<�e�kl:>Τ;>��N>���=G�>i��>hIþ=-�@�B?xa>+�/>L�>�o'>4�>�]�=I��o�>�57��1׽�9�>�u̾��Q=( �۴�D�2F>7��w��?�4>j���&(�>����B꽨ˣ>��>���)��>��v>%��>��>fd�>c)�>^�>��>� Ҿ�o>(��h_!�,@B�qR�]�Ѿ��v>,����#"���5����5I����O��&Nj�A+��RD<�+�<��?����Z�k��^)�$���}�?�X�>�%5?������>&��>��>��������&��+�G�?���?1<c>��>9�W?M�?�1�a3��uZ��u�l(A�e��`��፿�����
�����_?�x?yA?�P�<�9z>=��?��%��ҏ��)�>�/��&;�1><=q+�>�)��i�`�|�Ӿ;�þ�7��HF>��o?=%�?[Y?TV��m���">��:?1�2?/=t?Uj.?�p<?w�wG!?z6> �?l?�6?��.?D�?�5>��=��;�=�Í� ���۟ҽ#۲�>��v��<�rt=��%�8�];�}-=��<Z%��\��G�ӽ��Ƚ�<}�=�ۏ=$�=�q�>��]?:V�>���>J�7?z��u�6�q����c-?�f=�$������24���]�u>��g?��?{�Z?U.d> bB��E�yC>��>�Y#>�u]>�ӱ>z��~�E�	E�=�>�>B��=��[�x���r~�_U��=��#>��?�8�>�E��F��<�a;~�R�B��=DS����������h`�S�K��-��(�
>� 8?�?�f�<���7�+�ET]�%?�>�kP?/�5?��?�c�=��|(�W^{� ��>���>f�پו��'�����+��̎<uf�=���u�%��c�>�2L�!���B��2�V�=�����c�E�u�=�lT����"����7�!�)>L=ξ��_*��E-����G?��=\l����l��� �>���>��>��:�]��1�;�l��7�g�>�T�������0e��T��Q�>��E?ݵ[?Y��? ^�s�h��tE�����ҩ�ڪӼ�S?s��>�	?��[>R-�="¾n$��e��E�d��>���>�p
�p�B�i%��,��I��>c�>�i
?��6>U?fF?	g	?�e?�44?;?K=�>_L����@&?
��?U��=�bӽ�T�u�8��E���>�e)?�B��З>�?��?��&?qeQ?>�?a�>Ԙ ��<@�8h�>c=�>6�W�PU���`>�J?�ϳ>-&Y?�у?;>>��5��ע��Ԫ�!��=44>��2?t#?��?���>���>TS�=q>�6=\�@?��?��?�"�>}��>O�?��?��=��f>wB?H?Kok?�8}?I�?D`?�-7����M�:�r�"�1?=��>d��=w�>	|7='����r=�2��8�(Z�܁6���=)���8�=�q8>@*�>�<|>������@>X��-B��G�<>2o�� ����"��=�4��Ɣ=܇�>�`�>7��>��Sx=]��>��>�����#?[�?��?F}a�.{^�:�ؾV-8��>�,<?̮�=\�r�'����}���E=b}k?U?Ctm�����d?p_?�o�A�<���ž����6��Q�Q?2�?�h��V�>��z?
Ac?�,�>���K�l��⟿G5b��[^�h3�=��>���b���>�]>?���>�zH>Q�=��۾��w������?�Č?Cݮ?���?/�;>C�d�Ѫܿ3�߾چ�l,]?���>�瑾O?���(��φ���I���XӾ��ξ{�z����d�����2P������e0=��?�ih?�@i?��_?���3!U��^��q�+�U�&o�}��GP���F�CsR�Ȣi�R����Gþ��<ޙ;��P.�u%�?�0?�b����>����y���߾z:%>k�j���v�֛�=j�ʽ&#�=`T�=?��X '�n����?�q�>�κ>k�??�W���.���6���7��
��o�=���>��L>�@�>��f�k�U7��-	� ���&�Ū>3I]?��6?b�e?r$��}+���m�F �V��pȾ�3,>v��>_x>�]�Y��r+�'�*�w��q�^ԓ��%����h>7H7?ju >��=��?�4?����ԃN�xݯ���,��E#>]?]8g?*��>�,�>���z����>��n?k��>&�`>�����T��?��n������>��=�E�>զ�>50��Co�S��ފ���N��Z�<*"L?,ap�5�]���x>Q|P?R�_=Ҳ>6I�>r�2��$�����
M�^�>��?x"_>��>�̾69��H0e�X�����(?T?�>��F�*�->#"?	�>;̤>>��?*��>o���xй�?S�^?_�J?��A?�>��4=Y>��N�ǽɏ&�.`(=s?�>˩[>7m=
}�=Xp��oZ��8��F=u�=��ּ�@�����;����J<<jm�<$�4>��ʿ<�2���Ⱦ���d~���Z�
4��u�`��ܫ��&�4e�?��� ̾N\���X�<�Nc�+���u����^��?�<�?�}�A��D螿S5��1�<�KL>^���w�=<�)�c�G������X�,��A���:�ҳ\�;3��o�'?j���-�ǿ�����<ܾ�  ?�A ?i�y?�D�"�W�8�0� >�&�<�:����뾑�����ο+����^?B��>�S,�����>z��>y�X>Iq>+��^Ꞿ��<9�?��-?ϟ�>�r�,�ɿ�����ä<f��?��@�{A?�'�ka�]=�C�>��?$�=>?�0��N�z���/Y�>G�?ي?}�J=�=W�#��d?�T�;a�F��xݻ��=���=�%=*��P�H>D!�>����A�m{ؽ�O3>��>F��p�~D]��x�<�|_>� ׽𳘽4Մ?,{\��f���/��T��U>��T?�*�>U:�=��,?V7H�`}Ͽ�\��*a?�0�?���?%�(?3ۿ��ؚ>��ܾ��M?_D6?���>�d&��t���=D6�D���{���&V�Z��=W��>_�>˂,�����O�;J��Z��=O������YG(��l5�_��='@>ns=\}�:8�=�ɯ:�4����@�j�	<���=���>*,�>̈́�>}p�>�R?pcq?���>�k:>�������r�L�R�ҡC�n�6�#������V˾�����G��b߾�?��'�aí���Kk>�9[�z6��/x0��҉�J�Y�X��>~��>�.��O�5a<=$��DX����:>�	;���ݝ�yI���q�?��V?����D�;�B��yd�+�սV�?��=L��6�	����=�v�=7� =�j>����� ���F_�}:?�%?�ɣ�K_�4�=Ӓ(�����F?���>�ƽ%Uw>+�Q?+,������R>�7=O��>�>�lY=�X����ӽY�?==l?��C��?��[��>�,ž�iR�@�D>G#>8�+��ܼ=�>�>�w�=/�m�ws7>]���PΏ�:?W?�>��)���_���s�$�Z�3=ܺx?]c?�8�>�k?l�B?��<�S��F�S��0��m=�<W?�h?��>����Ͼ����P�5?5�e?��O>��h����O�.����!?�on?}?�I��XE}��Ւ�$��9�5?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?|�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>�������>˙r�r�?�j�?[�,�۠�������R���6���v�c�_>��=����U��FE
� 
�=���}���c�<��>,s@�Xs�?(�>�>p�ƿ�˿�e����#��������>���>3�>����ҟ��Mϑ���n�8O[��i��l��>�>+[��#i����{���<��ʿ����>�ּx��>M�V�刴��"��H<���>��>��>�곽�6��@^�?����Ϳ��ή��X?z�?u�?�{?��n<*�{�&�{�	�ٻl�F?��r?3�W?���ִ]�̻!�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�U�|=�>���>g>�#/�y�Ŀ�ٶ�?���Y��?��?�o���>r��?ts+?�i�8���[����*��+��<A?�2>���H�!�B0=�TҒ�¼
?W~0?{�f.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>eH_���u>����:�i	>���?�~�?Qj?���� ����U>
�}?���>���?~��=}�>ѽ�=�o��!���!>���=]�8���?EM?!��>Hd�=�:���.��?D�4�Q��\	��rC��8�>��a?s�L?~�c>6<��]q��� ���н�1�����B��V��Խ2�1>a>>$5>�+>�O�Ҿ��?Np�9�ؿ j��p'��54?0��>�?����t�A���;_?Oz�>�6��+���%���B�`��?�G�?>�?��׾�R̼�>8�>�I�>H�Խ����[�����7>/�B?\��D��t�o�y�>���?
�@�ծ?ii��	?���P��Va~����7�e��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?sQo���i�B>��?"������L��f?�
@u@a�^?*d~ֿr+���ھ�d���^>�Ϡ>E��>@x�<m1>l��=��=�8�<�A>ĕ>�D>�>�Nz>���>��u>j��m!������B���t,����K�6L(��m̾/��y1�����ZRսA�.i���Q��5�f��ח~><�W?(wV?{�?�R�>�Z���GT>����V^�����h>"��>(�>?:�j?��>v�伍_��s@�(��� ����c���>T>�%�>��>��?,ʽ��`>��.>i��>�=[C�<W�o=��<_8�>��H>z 
?�I�>�&W>�PB>���T����w�3���2 ͽ�}�?��o��JD�"�����n�ξP�=:�&?�-�=鎿�Uο�ͫ�F�C?{����/�n�׽�q�=F�2?�_X?�D">c�ξ0��=�8>�f�Qq���>X�/�ϵd��C$��%$>�9?���>���>�N���0��Cj�x�����p> ?���Κf�2؁�9�Q�P��+O>Ӟ>��B���������}�O�\��\<�@?"�?�Y�������U�^�J��=��=�H>���=P�>3���M4�X�� aB=&��=SC>�?.*'>p��=ި>�퐾��M�Su�>�,O>��>�;?h�$?�*�S�a���{�a ��Np>}�>�t�>���=VOC���=��>�k>�Z!��Hf�:����/���@>��|��jb�.����)=��Ὧ��=���=U!��<�}{=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�h�>cw�dZ�������u���#=_��>�8H?}V��g�O��>��v
?�?x_�ة����ȿo|v�G��>+�?���?2�m�pA���@��>;��?�gY?�ni>�g۾�`Z�%��>׻@?�R?g�>h9���'���?�޶?���?�5�>��?[T?�\�>UB�>8�����L��������l��Ș>��c>��νU� ��ʞ��Х�������.�EWO>s7"=P*�>��P�H�����=#�>g
����l�R�?,Q�>��>+oU=)�>C�>���>r$�=/ �L��2��~L??3��H�m��s�<��=�^�J�?�4?+�W�B�ϾW3�>}�\?ӿ�?��Z?���>�{�2��+ܿ�n����Ȗ<�tL>l��>]��>�Q��.L>��Ծ�\D�0̊>N}�>*]��:qپ( ���6���k�>T!?Y�>��=ֱ+?Q+*?�c>i�>.`G��0��2Cg�d��>�̾>c�>n�n??G�����Z��q��kИ���s�{*k=i�j?�b?՞>T����æ�	J=\��&�_|~?�2f?M����>K,�?t�	?��/?�g�>y�C���;C�d:�>��!?����A�EK&�B��L}?�Q?���>$,��`�սoּ����y��W�?k&\?GA&?@��*"a�_�¾�J�< #���T�r��;�ED�%�>c�>�x���y�=��>�װ=m^m��R6��f<�I�=x�>C��=�87��j��}<,?WH�Oփ�v�=G�r��vD���>eOL>����^?�d=���{�����w����T�) �?��?�j�?����h�u%=?y�?Z
?!"�>rL��=~޾���Yw��x��v�J�>���>�l��徵�������F���
ƽ�۽���>z��>�/?j�>�G>LJ�>�䱾8G4��`����a�R��h��3�(C�}��1��z�d�#5�	�˾���O��>��c��V�>��>�J>�#�>_[�>Cu=�/�>cg>�`�>���>ڀ�>k>�/#>�:(��Е��IR?���=�'�ª����/B?�md?�-�>�Ci�s�������z?���?rp�?�1v>�yh��++�p?�1�>����m
?�p:=���̈<;T�� �����G�4��>�g׽6&:�jM��f�6f
?�/?r����̾�J׽����&>|�z?�t=?��.�(E2���w�p�-��=\��݉�(�߽���ɾ־#Q���㜿��c�ߡ���5��-g���)?x;q?h�
�0���X�怿�su���}>ه�>��_=w��>f�?e�*���K�k�e���#�ܞ�Ҙ]>mN�?�	�>A�I?βO?ެ_?�i&?B|n>�/�>ξ�s�>���=\E�>�f�>~�$?�u9?��?B	?o�?hƆ>�}ҽ�4���V��_?���>�e ?�?�=?B��Qc8����=G��dW��E1�%o����|=�d<S;kN<>
l�>@W?���Ѩ8������k>��7?%��>���>����'��B(�<���>��
?�E�>���vxr��^�dZ�>?
��Mr=��)>���=�����Nʺ�i�=�m��.�=�����z;��<Pk�=֔=�u�p�~���:��;ެ�< u�>6�?���>�C�>�@��/� �c��f�=�Y>;S>{>�Eپ�}���$��v�g��]y>�w�?�z�?ɻf=��=��=}���U�����H������<�??J#?(XT?`��?{�=?_j#?ϵ>+�jM���^�������?&h3?7�>w�=��@r��캿�	�C��>�G�>�E��=޾��(����1A��M���e\�L�W�}o����Y�[���
�Kc5�C�?���?C�R>��j־.����!����>�� ?�-�>N�?:�����i�3$ھ��#>��>U�?�>/;Q?�i?qxP?��>�o
�_Ԝ������v��z�>iQ?2?D?���?̇?���>��һ�g��8�����3
��S���R���=s�=�1>�?��?��=�s�3.��	���O>j��=ڊ�>$��>�?�8�>������G?���>\��T��x夾㺃�p|<���u?옐?@�+?b=���E�U;���O�>�m�?��?�4*?ݙS���=J ׼�ܶ�2�q��%�>;�>#5�>,�=�uF=cM>�>���>{5�O`�&r8��yM�w�?�F?�û=ɪƿ(Es��&w��	����<�Ր�]�^��w��~�T�}�=�����c����[��I������F���,���zu�*��>��=�$�=�j�=��<����<`P=N'�<,'=sD��V�2<�J���������;#��<}Q=2G�Ё˾��}?�>I?U�+?:�C??�y>qT>��3���>2^��=A?d!V>Z�P�\�� {;�ģ�����g�ؾk׾kd�9ӟ��C>b�I���>�B3>�@�=U��<���=1@s=eێ=�R�.H=�=oX�=�b�=��=��>@b>�6w?X�������4Q��Z罥�:?�8�>f{�=��ƾq@?��>>�2������yb��-?���?�T�?>�??ti��d�>M���㎽�q�=J����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>è;>�>��Q�u}1��a]��e��`�d�!?w�:�"Vξ���>��=Q2�hɾ�v=S�2>:�A= +�AP[�Y��=vz�!8=�Mi=V�>&�I>�$�=F���"�=#�?=ք�=�vR>�+��QH%��&�/-=���=E�b>8�!>��>��?EA0?��c?�K�>4�l��˾Nֽ�+��>4��=���>��=/-]>͖�>��3?��@?�FG?G�>\�T=��>���>-z'�j-g����Y��b\�<���?엃?�ӵ>
��k�O�v���C� ý�?W�.?�?}H�>�I���ֿ�)�_i�%[�=!>���=} �=\�n>FE�=�N�/5��Q�=�2>�4�>� ?�g�>�|�>|α>�2�>��O>(�=ri>P� =��f=��9�c��޵'�"\��ۢ#�|���	=u_��fB�< 6*>	�V=�6��Λ����=�>�>�>�m�>�w�=�$��L$.>�d��t�L���=P*����A�]�d�z~���0��r5��[@>O�Q>�E��㑿v�?	�c>�/C>���?�At?��>����پ�蝿�,]��O�p�=�$
>
�>�#c:�^e_�Z�L�V)Ӿq��>�>@Z�>�{>E�.��9�'�d=�Wp8��c�>�ц��C-��"��o�A'��4u��f(f���ܼ�7?h���M�=`�?"G?5��?D��>#t��m�;�=>��q��f=�B���U�k>��?��!?;��>��<v@��B̾�����ڷ>�GI�i�O�ĕ���0�K:�����>������о�)3�h�������B�s\r���>��O?��?>b�%V���UO�6���X���g?�tg?{$�>�P???x	���{�n�����=��n?0��?,;�?��
>=��=�!�_��>�`�>��?��?�?�����>�>��O>VX�<�=~n>�FE>��1>^U"?o�!?��"?R�޽v��I���	���9�sQ�=��=y�>1�E>m�o>l��=�#�=���=�m>���>�>�>_ei>-��>#מ>��t����j4?kA8>��k>^m�>��D>�A!>�`߽�Y<���=G����b�Ι������t�YV>��ϽV��2/�>��ȿ���?!�=N���X6?s+Ͼ6CD>M�>���>-L��Xb�>��=��>�?��>��>���>3�>5�Ҿ9�>!��`!��YC���R�۰Ѿ
z>}A���!&����2�����I�����ib��j��'���I=�ź<�;�?I(����k�*�)����J�?�p�>�6?e3�����0#>���>�|�>�#��`���η���Q����?j��?�;c>��>4�W?/�?�1��3��uZ��u�o(A�2e��`�r፿����ݗ
�O����_?��x?�xA?�J�<�9z>��?~�%�Kӏ��)�>�/�';��D<=�+�>a)����`�h�Ӿb�þ�7�JF>C�o?8%�?DY?LSV��WǼ~q>pqD?`.? g?^N5?0�C?}���A?�>�?`�?[�5?��@?i)?Y�A>ߣ^>��=��=�[�������G$�x�S��
��"t=!���0�=�r��t =fFc��s*�;A=)��=�=����L�=?,�=�=LŦ>��]?Y�>)��>��7?����]8�笮�`/?c�9=�������zh�����>J�j?��?�_Z?�d>��A��C��9>�t�>�;&>�[>bU�>���#�E�_��=Z>��>�W�=@P�vҁ�ޯ	�G������<��>pd�>�>~>@�����)>�����By�\c>��R��f����W�ͱG��u2�|�w����>z�I?C#?I�=M������;e�[�'?4�<?��M?m�~?�ʘ=�۾�!9�	�K�^ �E��>B	�<�j�h�������9�	{�l�o>�����T��0a>��h޾vko��QJ�&��QMX=���x=K=f����վ	~�yz�=L{>I;��� !�4B���򪿓�J?�Fn=վ��G�T�U����>[�>W]�>�_@�N}�u�?��9����=�s�>�<>(���^K�{�G��'��ϝ>i8>?L�K?�*�?������E�o̠�1��������<C?E��>���>�>=��n=RE�����Yj�X{Y�=�?^��>�M��=�zP�<�$��s��I=_�>�A�>��\?��?ldl?v��?�%?s&?l�?��i���4�:?(/{?���L��kϾg�c�R�}�Δ?��F?�
�z-?dGd?�GI?\�?��`?�N'?&�>�YH��ڏ�RU\>��4>RL\�\N�����>��;?���>�".?�e?e�=�dE�/���ʇ5�w��<�Qz>�I?�?d�?o�>���>��u����=n�E>7�u?|�?�ߊ?/�>t�?���>�gq>�>�_�>_X?3�?�H?�Zp?  ?��h>=΢<=�I=h�	��򮽅�C�_��=�iA>i�=;�=�Rh�C&!;���;oȞ=��\<" �=�,=���=���=�V�=LI�>	]t>�+���0>�ľ�È��zA>�Q��Q~���i���H:�SA�=�1�>�o?Rc�>a%�֋�=�>���>j�T(?$?�?��9�]b��ھ/K�9&�>�9B?{��=�<k��6����u�se=��m?oe^?�2X�o��A?c?�]?N��k�7�԰˾�/��>�����N?d�
?ewM�`��>�"�?Fur?�D�>�kZ�'{h������Af�	����"�=+H�>����k�Ny�>D�7?�W�>$�v>��>����w��N����?^�?�x�?p��?+A>�np���߿أ߾{M��?�b?am?i���T:?�*�={%�.�������K����Ⱦ,T��1���?侦@S�����Jh4��}>19	?��u?�X?�Յ?j���]b���M��B����w�t�Ga0�dP���N�S�9���l���xR�$����"�=-�~�WA�bx�?�(?I�/���>I�f��L�̾w?>����ݡ��Y�=[�����==t�X=�6i��0�Mp��� ?嫹>��>j�<?��[��w>�n�1�B8�͇���x4>�0�>��>#��>M;�;�>-��轰Ⱦt��(sֽ]c>	�b?�S?9�?��׽���ׄj����֬��ؽ	��w>�A0�E�š
�8[�z�"���H�����׾`/u���턼=�??�hf>�c�=�_�?ܹf?�Q�ˢ�����^���A>Q�A>�ad?���>�a$>�й��!�Fd�>�m?���>��>\����>��x{��T��� �>R��>J� ?��`>��K�rv^���������G9����=�f?A��mc���~>uT?,�+��T�:�C�>T�$���=��3V#���>�O?��z=��B>�R¾��	�^Az��:���'?�?�P���o&��b�>��?���>9�>�?�j�>������5=�z?ka?n8N?��G?�\�>&Xj=��Ͻ�u½��!���=�>��a>[�=q�>$��yY�2�׶K=�q�=�uY��dX�Og�<8�:Nm9��-O=�R>θܿn�W�%�߾�o���Ң���l��� �+���D.���ؾh���r�t��Z��@�<l'���u�����_����?���?�����A��:���䌿��qQ?�d��S��{�Խ� ]��ʽ����i�'���t��+��7��Y�!?v-ľ�o׿"�����3�\�T?<<?�w?�bd�;> ��処����I�8���о�����ܿ�ǔ���u?LV?�W������=��?�>s��>tu�͐�!|>*�>�z�>'�?���=(a�-|ɿ�H�<��?�v@N}A?�(�����U=��>ߎ	?)�?>�N1��F�����U�>�<�?��?�M= �W�!�	��e?�a<��F���ݻu�=�:�=S?=G��6�J>V�>7���TA��-ܽ��4>7څ>��"�����^����<��]>��ս,��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=�n��Pο<�$���%��^\<_b=u�߻�D�������W�侚����)#���=��&>�:r>K��>�y>�R>_?9sv?kA�>~�>:��b���w�ؾ$��=��l�����4�F�\�"��ˊ�����u2۾���R�3��3�M~޾@�C��z<M�X�}݈��ZS��p�3�@�WA?�\M=$A��.�2��Ҽ�|���%;^�a=�ix�j龨0G�KC~��k�?��E?������7�B�(�ZH�����ub?"�?�>��|���>�}��짽���>
K �D'��4S�Z�Z��`>?��"?vy޾?�����=5���ݑ���*?g�?��<��>�V?Z9B���=��>�ʾ>+��>±>���t��R��yQ:?��x?Y����qu��>��ʾ���S�f>�Q�=+�t�:e_�6e�> �f=Fr��J��n�G���>d(W?���>��)��ja��� �fV==��x?�?.�>_{k?��B?�٤<�g��@�S���	dw=��W?�)i?��>T����о6�����5?��e?��N>Gch�f����.�U��$?��n?%_?�}���v}�a��0���n6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?s�;<��U��=�;?l\�> �O��>ƾ�z������3�q=�"�>���ev����R,�f�8?ݠ�?���>���������=�M���ܩ?���?	��2�==\��c~����%���`ټ�N�鹯����F�E���̾9(�" ����=��y>�J@�F�����>ڝ1�S'���Ϳp:��i���l���?�ɋ>s�e�%����|]���j��;���(����QO�>	�>����4���'�{�5t;�������>.����>"�S����<���(�5<��>@��>���>cB���뽾ę?_��?ο2���ҝ�w�X?�f�?�n�?(t?�9<��v�#y{�<��e.G?�s?Z?>=%�G]���7�<g?A��$���w=���&E�U�>�@?�Ev>�xM��ا>s>ɽ-1>.>����ҿӼ���$���?(�?Q(ھx�
?J��?� /?���9���|�]���y>�O?�������~5���k�ySk��vJ?�%7?@s�<j/=�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?  �>r�?�i�=I]�>�b�=�ﰾZ�,�pt#>�J�=��>���?��M?�G�>�H�=i�8�I/�AXF��CR�y ���C�F�>��a?SL?KAb>����2��	!�<@ͽ�a1�K��.F@�̦,���߽""5>-�=>�>:�D��	Ӿ/�?N��ؿZx����'��64?��>!�?0��bgt�Kr�_?j��>���1��6�������?I�?X�?r�׾b�ɼX�>S�>o�>&�Խ�����O���U8>�dB?E�f0��5�o���>s��?��@Lۮ?�h��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?pQo���i�B>��?"������L��f?�
@u@a�^?*C���A���Ӿ�6ž�?>�!C>�i>!.�Dc�=��'�B5G��f(=M�)>gn_>z$1>��s>�,">��r>S/a>H��T%��ɛ����.84����@W����' �O6;b�%��ؒ� �þ�3J��
����,�S���|�8?>�TS?ȓS?�Zr?�f?�B���.">c ��`�<#����5�=�3�>B�/?3�P?�-?���=Τ����a��k���⨾�Ӆ�c�>fmX>��>�=�>0�>Y:���,>XY8>P�x>��
>�)|=(����J)=bfD>�;�>���>o3�>7 �=Z��=����[����f��m���1��V�?7#پ�Ha��Fk����������M_:?q��=T�����ֿ_���]?�����1�:6B��>��d?v�:?��>�!�l���8�y>��i��m�=���&�,ON�ݟh>��N?!�f>�u>њ3�^d8�$�P�"|�� i|>n46?�涾�D9���u��H�Kcݾ4CM>�¾>)D�uk�������ti�_�{=$x:?ȃ?�<���ⰾ�u�C���UR><\>�m=Ow�=OZM>q[c��ƽ 
H�Pq.=9��=ެ^>��>k�?>佀=
0�>�\��J��1�>#`[>��]>0�B?$'&?�H�&���9���nJ�NQ>��>��>>�>�'9�*��=ٸ?�eI>�p�B�c�
��>T��=�>xM�� �.�l��l�T=𷮽��=�}�=��뽭D���=�~?���*䈿��e���lD?W+?^ �=��F<��"�B ���H��E�?q�@m�?��	��V�C�?�@�?��B��=}�>�֫>�ξ+�L��?��Ž.Ǣ�Ô	�D)#�hS�?��?R�/�]ʋ�7l��6>�^%?��Ӿ��>�g>��t������w��0�=��>�`C?aP�n�i������>���>��辢R��xLοY�k�>�
�?�?��j�Å��4�G�=�?���?�|g?{@>����p�;�E>x6?%W?7�>y:�.��?ϼ?�Մ?��>WJ�?��?�H�>|��=�Ͼ\���%��9��l�3��=;=EЩ���u��"D�{5���6j���O�ʻ��~�>�YM=,�>{������؝t=-m�<_b�������j�>�A�=J'�>ǎ�>��=�	.>�r�>��:�U8��l������(M?~-�?���ۅp�ƃ<�)+=z:��;?�Z9?gm!��!���¸>Ys_?�u{?vC[?$��>q��0:���R��Tծ��sm<�A>vs�>N0�>�1����Q>�ҾܨG����>s��>��i��ݾ�pd����آ>�?�\�>��=× ?��#?��j>�&�>|_E��8��o�E�״�>���>�I?��~?$�?�ӹ�{Z3�����桿�[��=N>_�x?zU?W˕>I���/�����E��GI�����1��?xg?�H�]?3�?��??�A?5&f>����ؾn�����>�!?���y�A�<>&�RW��?S]?s�>�ܑ���ս�ռa�����1?�$\?�F&?�T�ka�þ�e�<���(X�W�;F�&�>D�>r߈�c�=�H>ѭ�=�*m��36���h<�@�=ig�>S=�=�6�L!��)5,?C�I�0݃��T�=M�r���D��.>��K>����,�^?j>���{���������U��ʍ?`�?��?��/�h��A=?y �?�8?(I�>�Q���޾Eྣw��>y��^�K�>r�>�c�%u�F{��$����D��JPƽ��Y����>z�>BX�>�8�>��+>ڍ�>*-I;k�ٹ�`����k�1O��6@�C5.��+� Ͼ�Z�x�=N�U+��lq>Jk����>�y�>��>��>|c?��=�h�>�x�>
��>�ѣ>�\>�In>s�>��˽�@���KR?����/�'���辺���j3B?�qd?N1�>Hi�3������x�?���?Qs�?�<v>h��,+��n?�>�>>��Qq
?�T:=e;�j<�<,V��K��`3��x�B��>lE׽� :��M�nf�Xj
?�/?����̾�;׽����?��=\�?��2?Z�#��G��a��e�o�S�g���\
������c+�#o��$��S%���&��l�=��?pg�?ي�+��_�.Am���O�S>-��>�Ϝ>��>� +>Ǐ�z,3�P�M���!�;�]��K ?�m?�e�>C�*?�5?�d?�^S?H8n=
�>�-�����>�z�>�>��G?�o"?��^?"�I?p�A?�b5?]A�=z�\���c��i�)?78#?�&?�}�>�}�>�᤾��S�P]=D����*��AD=]�?�����ҏ�lPl=��^=��*>qW?���_�8������k>"�7?���>���>����%�����<U�>ٵ
?xF�>4����yr�c_��W�>*��?���Y�=g�)>X��=�����Һ\�= ��� 
�=�9��No;�,f<�|�=\��=�&s���t����:�Ї;�j�<	t�>R�?Z��>�ǈ>1����S �,@�)�=��Y>7�T>��>�Uپ�B��� ��i�g��w>8�?�S�?��l=#}�=>"�=<4���^��.���nS�<e?M}$?hpT?�Ȓ?�x>?/#?8>z�C撿����=��K~?�!,?���>7��,�ʾ���3�8�?'[?�<a����Y;)�O�¾��Խ�>:\/�0~����D�"u��m���~����?p��?�A���6��w辽����Z����C?F �>�X�>��>l�)��g��$�i3;>)��>R?vB�>�O?kI{?�\?�W>n}8�j�������l�?�s$>s�??�܁?D̎?Hy?8V�>�c>�[&���߾�7���d!��T�������^Y=l�Y>�ɑ>Nz�>ǩ>�v�=��Ƚ�ҳ�	�?���=�a>�^�>!ʤ>��>x>0�<� H?(�>���w�������n��7�E�+�u?|��?J�*?�==����D�����o��>�o�?<�?n�)?\�U�<j�=�k׼Q���{@r�2H�>G�>�G�>t��=G0D=�>���>{�>������*8�N(G��q?�_F?���=��ſ�q��p�q˗�J�d<����A�d��[����Z���=s�����ȩ��\�\ˠ�Ϛ���굾I���#�{�^��>
��=!e�=
��=��<�Fɼz��<�>J=!�<
�=��n��2r<
9�]xһ���Y���^<H I=gj��ej˾�~}?�1I?˜+?�C?4Ey>]�>_t/����>j���K?+kU>`T�9��Z�;�俨�dW��W�ؾ�.׾v�c�՟��		>�{K�Cg>�B3>��=�؊<+��={lp=�p�=8D7�[=���=א�=�j�=��=��>�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/> �>>�	>՞S�q�2�� ^�{Pj�p8d�^�!?q6�ǭ;���>L��=�׾�vþ��K=gMA>w��=6��_]�X̘=�h{���;=�$`=2~�>��?>3��=B���;��=�6="S�=��Q>�{+��J��k*��H=�`�=�k>Ћ0>��>�?�q1?Sg?�5�>��x�?�ɾ_?��@ǌ>dy�=P'�>�E�=.�M>�><H7?�gE?�aN?�ԯ>HHt=@8�>��>g`)��gn�&�꾺h���ܶ<!�?堇?���>��@<Y9V�"�)9�z
����?A.?)�?�Ø>������2}+���0��w��[��=��>�����T3���)��&۾8�ݽB�;=R��>� �>vB�>��>gۇ>nYg>	O�>l>�`{<g�ʓ̽���=$a�J� =^8$���<��xX��6����=��=,R=���<R��;�j��O�=���>�0�=&��>%�6��{߾��=Mp��AD�=�->�ϾiT�G[�",y��>��䕾"��<Pζ>��ѻ�����?ʈ&>��>0�?�^~?�^>�jb������v�	����L�=�*v>:�ɽFG4�JO��U�����$j�>S��>V*�>:�">[�4�"K�t��<�1�*��l?�֢�הǽ�3� y�h���T��ߚj�8��=v@? ŉ��W7>�K?�QT?�T�?��>o���;����#>���QY�<~t�~|������k"?�?��>����j�<�tp̾�e���J�>\RI�o�O�~���@0���g*��� �>������о�2�P����2�B���q�'=�>��O?ظ�?j�`���i.O�x����?>?�)g?*V�>��?)�?��#�ր�LI�=L�n?z��?.��?|>R��=�g��C��>d�?}��?���?% t?�"9��*�>q <3�>-���T{�=.�>)��=]�=�?�n
?�	?����n �V���P]�(�=r�=>ڑ>,�>j�u>��=��=�]�=)
[>J>�>�Ȑ>|h>=]�>Ŋ>0Ȩ��wݾ� ?�c</tp>�5?�ѓ>�߇=$ȉ>���=���=8Z7���-�6l.�'��^z���<���=�=@��>[ɿ���?uY�>V{��*?^��#a��o�(>z�����l�9�>��A>���> �>��>���=Pܼ=�@>� Ӿs�>�'��c!�0�C��ER���Ѿ{'|>oS��m�'�L�����uI�G������i��M����=����<�T�?�-����k���)�����A	?%�>^�5?f���	w��y[>�^�>U�>kF�� ����0���,⾲�?�(�?\qY>w�>\\?P?I.�!14���T�Ĉ}���C�:�b�#!c��ڍ�L킿�3���eR?Q�m?L=?Y��= �l>_P�?.�c���K�>�@/�B�G��{'=�>*;��^K��.Ҿ�;Ծ��%�xO>��g?WE�?vi?��O�Vs�=��=c�.?I# ?8#s?Q��>1?c��R?Z+?."�>="?5	Q?��^?��!?Э�>+��>'���X�8��%_��pp�2���Z�^�� *>��=\G�=)�=PN<Sӕ�s8��T� Cؼ@���$퉽gni�t�=ԝ=xǦ>Â]?�D�>���>��7?�P��P8� ���!+/?==$h��ڕ��7?���t�\x>��j?���?2Z?��c>��A���B��
>��>��%>t�[>	N�>k��.�D���=&E>��>�a�=OL�!�����	��������<�>'��>�0|>m
���'> |��1z�8�d>t�Q��˺���S�A�G���1���v�8Z�>��K?��?h��=+_龈+��If�d0)?4^<?�NM?��?�=��۾��9��J�	=���>hJ�<�������#��p�:���:��s>�1��`����[b>Z��5޾w�n�� J��~�1�N=?��t#T=��N־�T����=-�	>ȣ��� ��"��eت��!J?^qi=2M����T�쉺�{_>���>x�>�g9��Nu��m@�k��� J�=���>k�;>������qG��V����>�w%?��>?3�?*���b{�N��f,�G���R|Z?!�=�?�T�>�:I>�S^�*��w~�G
t���>�|�>>_/��SA�J���2�7�4�n�4	k>Im4?��>�-?�۝?�+4?��j?�$�?�?���>��[>����9?A��?��B�^�m�پ��u��@��՝G?���>����$c5?0fn?s?�O3?e/|?��B?���>{�þ�S�1��>䚲>�@=�=x��"��>��+?��>0(V?xo?�+>#f��p��DR�)f��h=w�9?a	?�-,?�,�>@<�>���2�C=�Q�>��l?�^�?�?���=�/�>���>�2�>����՝�>�-?��?�[,?]�h?�p ?��>!�=.񑽔\t�[�/���ż�n���gq�|ܛ=4>��B=�#q�
P#;�-�̌U�XĎ=�n�;:�s=JNd=Lh�=�`�>��s>�
���0>��ľ�P����@>i����K���֊���:�ܷ=ƀ�>G�?Ŧ�>%X#�	��=>#L�>����7(?��??�c";�b�e�ھd�K��>2B?���=E�l�����F�u�c h=y�m?�^?��W�'+��K�b?��]?5h��=��þy�b����b�O?#�
?j�G��>��~?V�q?I��>�e�$:n�'��Db��j�Ѷ=Er�>IX�G�d��?�>b�7?�N�>��b> %�=cu۾�w��q��n?��?�?���?+*>��n�\4��`ž���-Dl?��>p1�y�)?K�=��.r��r��d���ﾾ�ݖ�I����ι����M�{�ǫ.<��=�N?Wo?a�t?7ƍ?n��\(x����j���'h�Y/�BmF��O�1�%���:��mk��<��4���������=�{��C��?��&?5<4���>Y]���S�
�̾XfD>iS��N/��	�=Rh��/�.=��,=�f��Z �`���&�?���>��>%�??�G\��`<�C�-�p�:�i���(>:�>R��>���>;w���(��3�Ӆ̾���޽���>*c?^P=?䉂?m�@�^
��OG��&�c޾7}�%��>罧�$���������og7��~C��ɀ�y ��=��.I!�����3?�w�>�yB>���?tDd?����uE/�Z�t��>�o?�U�?b-?�>�▾ya]�E��>!�l?���>ચ>Mˌ�.����z�Q�Ͻ��>�´>O'�>~�e>��J�خ^�Jŏ�������6�~��=�]f?��~�w�k��Z�>uN?�F��:t�<�@�>F"���"�CC꾶����>�?S��= D>h:��wK�Q
t������,?��?�?��4�*��Y�>��?c��>�ٻ>֌�?<�>9w¾t�a=��?�T?F=M?c�K?��>�K�=�}��,ƽ&(��g=`�>�c>\v[=|�>x,1��G�	��7�<�j�=�jJ��H佟|�;�=ٻ�/�>��<5B>��ؿ��E�#Gھp(�����Cp�JH�d���U��%t��-���8��;ｿ�@�OQ�۴O�N����7P���?b��?+BѾ1���%���|(q�����68�>�@�1�,������,�q�x����\9�����)o��!n��]���? ��pԿ�颿q�4���O?O&
?:i?z�<xp�����ՃA>�)=��ǽ;��~���j�DI����?�z?�;��&9��u�>ֆ�>P!�>�-�>�G����#4<=�O�>�/?9S?���(ܿRw���R�;v��??�@�|A?��(�����$V=���>��	?��?>rU1��I������T�>f<�?���?d�M=��W���	��e?s�<U�F���ݻ:�=�C�=F=X����J>�U�>U���XA�/BܽK�4>{ׅ>�m"�	����^����<y�]><�ս�8��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=����Ŀ$!�4\(���g����	ս\��s<%3<u6��Lz��b�ܼ��=���=�KS>r(�>$�*>��d>�W?l@j?��>ƴ�=��5��&��v#ھ�<��.��2��y{���`���A����6���	�Ӄ�!����0�A��̈=6�^�����$(-���S���-��_=?Az�>�<龈iP�LK��S���x��x� ���p�.l>�18S���?99O?����l�Q��3�~A5=�A��SM?��n�i�+�G����r�=����c�>�"�1�P��D��g>��A?�
>?=�׾���8>�E�_�b>�>?�?�s�<��l>�8l?�ŝ�.;�HK�>G
?0ӣ>W�?k�|�	k��%G��)?71l? *�τ��_�>��%U;��o���<@>8��Ks��m��>2Û�w���?ܵ=�����ɼ�(W?���>4�)����]���:��F==�x?~�?�/�>Ywk?��B?6ݤ<Ih����S����qw=H�W?�$i?��>⑁��о����5?�e?��N><gh�����.�fV�%%?��n?�Y?�w��?q}�������m6?��v?�r^�is�������V�8=�>q[�>���>��9��k�>ב>?�#��G������Y4�Þ?s�@���?"�;<!"����=�;?�\�>˫O�6?ƾ�z������m�q=�"�>L����ev�����Q,���8?Ϡ�?_��>�������>r �����?�Փ?��ݾק���߾�	���������A*����"�j�O�*i��{A�r��'v �)V��]s�<G�>.�@ V�s�>-�h��D鿃�ÿ򽅿M���P���Y?V�o>���<��`�n���1�)%���Q���/�M�>��>��������{�wp;� 3����>,,���>ױS�5+��i���+F5<�>1��>���>~@��<齾iÙ?�b���<ο��������X?�f�?oo�?q?Iu:<��v���{��j�R.G?\�s?Z?A%�V<]�8��_n?�����`v�d�Z�E1X�5��>��z>��p>;ʾ:�=zHB�s�>X����@e�ȿ�������Jֻ?���?�쾝J?`+�?;c?��"�����IBվT�8��,>��L?��<������k���T�ܛ��r�4?�#N?�ƽjS�]�_?+�a�N�p���-���ƽ�ۡ>��0��e\�N�����Xe����@y����?N^�?i�?Ե�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>	�}?y$�>��?]o�=b�>)e�=��@�,�Nk#>�"�=��>��?��M?�K�>5X�=��8�;/��ZF��GR�v$�5�C���>��a?�L?�Kb>e��4!2��!�]vͽ�c1��L鼺W@���,�q�߽(5>C�=>%>��D��Ӿ�[,?h�$���Ɲ�NqA��UD?�s>��>�B��ۈ���w�f?o�>���=���}���l̾�6�?��@a?��Ѿ��;��>	��>I״=Ͼ�����X�=�>g)#?b�N��ō��ٗ�4�>u��?���?�?ՎS�'	?x�BM���a~�����6����=�7?��{>���>��=�mv������s�Z��>�=�?px�?|��>�l?p�o��B��2=�3�>�k?�t?#k����B>��?���6��H��f?B�
@�s@X�^?(좿��ݿ:����W���hݾR�=��=�);>j�b�V>q��=����Ͻ�۹=�3�>\Jj>1\>���=�;>�g">�@��t�!������!��6�R�?2�����s����o|���'���־�À�۝Խh2Ľ�N��sX˽�˓�4�=>?BT?^R?��o?�@?�L��&.>t��K��g�B�5�I>c��>uXI?�O?G~??��G>�u�z�h�)����V���BS��>/��<�C�>�>0*d>J9=�9W>W;>`�h> 8��#��<�ܐ�ɑ�c�>�y�>���> ��>�)>n�+>h���C��	�v��i�m�ݽۢ?Hx���FY����������h��9k;=��'?燿=�Y��pmп=@����S?k��Y �rD��(2=��@?�C?4u>��Mb�2w>ϥ���^��	)I=0k&�I����L�lEV><#?9�f>�u>!�3�d8�&�P�h|���k|>46?T붾�F9���u���H��cݾIHM>ľ>I
D��k�����=�7ui�u�{=Yx:?	�?�;���㰾��u��A���RR>=\>7Z=�k�=\M>�Qc�a�ƽ,
H��m.=s��=]�^>h%?z,>E�=j��>}ᙾs�O��K�>��C>��->�>@?��$?����\�����S.��_v>�2�>2��>]=>��I�Q��=SJ�>}b>�?	�N����@�D�>�6V>�ux���]�}�p�[a=�ܘ����=>p�=����I<��A"=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�h�>��۽������n~��P>���>5NB?�l�=�b���'�z�
?�f?&��Fܧ�N{п<E���4�> Y�?�q�?�u�K`��q 7���?��?D_?Q�>�ľa��GL�=�$J?\�a?cd�>��=�;cG��?��??�?�΂>p��?���?H�?��0=X��W,���4��!����A=�if>�����J�8NS����5���WE;���'�Y �>uO�<��S>�;�>Պ����m >��|��4ڽƔ�>���>��>�>�!Q>h��>5�p>˷��P����}��-����K?���?���1n��:�<d��=2�^�|(?�H4?ގ[���Ͼ+ڨ>��\?���?�[?�g�>S��=���翿�|��E��< �K>�1�>�J�>4���LK>}�Ծ�/D��q�>:ɗ>���?ھ�0��R�B�>d!?8��>�Ӯ=*P ?O�#?OQi>�v�>�D����$F�9��>ȏ�>�?�Y~?��?6ܺ���3�l���ۡ�$t[���N>�x?�+?[x�>o;���{����`�kG��2��&��?pg?ͶݽV�?�G�?�??�+A?$�e>�����־H	��룀>��!?aT�M�A�06&�8���?�_?���>�>��{ս8+ռ����F���	?3#\?	=&?��#a�4þ�2�<@G!�"`N�|E�;�`C�2)>h�>�H�����=��>�߰=7m�E�6�O b<G��=-Q�>�.�=�[7�I����8,?�'�Wh���~�=cxs�qD��Du>Y*E>*x��x�^?�E��^{����Jל��+Y�c,�?'+�?q�?Lg��4xi�:>?�?�?Ul�>/;���ݾ��޾"{�j�}�i�����=�Y�>ڱ0��������0��1X��Zuڽ�R��a
?���>.�>q
?>[��=Ϛ���^����Ek$�P|p���W��K���A��$��߮��#�����=`�Ⱦ
Lo��d\>���|�>��?��o>�;�>�O?�M>և�>C��>p�>-��>H��=$�=G�)>̖�������KR?����|�'��辸����3B?�qd?1�>�i�<��������?���?9s�?�:v>ch�/-+��n?�?�>����p
?�R:=�9��@�<�V�����43�������>EF׽� :�zM�of�<j
?�/?����̾:׽|t��KCp=�P�?�)?i�)���Q�$�o��W�a&S��@�h������$���p��U��H��e�(���*=�}*?+!�?����X謾<k�?�ff>j��>��>;��>ՀI>	�	�R�1�z�]��@'�X����=�>AN{?��>A�2?��4?�W?��c?�p��,��>�O��wR�>kt��>��#?�0?W�??v�S?�I$?��U?�]O>p�������о.(?�;	?�c?A�%?�>�����9�d��=��'����������k>�[5�k־�s�����^�:=@X?m��S�8������k>��7?ޅ�>���>����&��p�<N
�>��
?�K�>
����xr��\�$O�>c��?u ���=V�)>!��=?����̺�O�=�=¼��=3����;��d<���=��=~v�m*�����:��;�<��>��?��h> �d>�rf���������=�(�>I!M>ב�=�����t��9l�i>>���?�?E��=i��=({�=R���Ͼ��������=�W
?��$?��i?��?�vG?�1?n��=������p��Ҏ�@�?i!,?��>�����ʾ��ȉ3�Ν?t[?�<a����;)�	�¾��Խ��>�[/�Z/~����:D��򅻬�����/��?࿝?$A�P�6��x������[����C?""�>9Y�>��>7�)�J�g�S%��1;>��>?R?a5�>}�O?��y?	�[?o>��7��릿�����&J�c>�PC?`�?b�?�^x?�7�>&�>>�!��u�����y;8�L.�tRo�bU,<�F>��>	:�>ŕ�>���=ٻ�귽:]�Q�=f�M>�&�>���>��>��q>�|�=�jK?���>�l;�j��Y���5���A�� �?�?�9$?�,$=�:���>;�0�i�>鞪?d�?L�1?�|����=a�	�ԥ��u�B0�>�ٷ>���>��4=�~�=�A>ܞ�>+8�>)��^!�K�5�C괻a ?�M?I��=	2ȿ��r�Qqk��Y����(<�����i�|����8�a2�=�x��bG��L���V����I���0������%ix���>d�=S>*��=D�<�A�u\C=��='=�1= !u����M�E�n<UÆ������:"kP=�%T��}˾�}?DI?{�+?:�C?�y>�e>�\3����>3���@?n�U>-�P�dj���m;�ʩ�����	�ؾ��׾G�c��ß��R>.I���>�G3>���=縇<�?�=ccs=���=TL��^=�<�=��=^�=���=��>�'>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/> �:>n>��R��1�|3[�df�e�Z���"?R�9�4˾2z�>��=~�ݾ�=ƾ�!==}J<>VSg=O���\\����=i�}��&@==�h=k�>��C>��=sU��=�=��R=��=�P>,�j	H�^K.�)�==�)�=�od>I'>�D�>?41?�c?��>�r��;�oƾ]��>�=��>���=�Q>�n�>}�9?��F?x�L?�*�>��Z=�>�͢>DB)��m����&Z���v<H��?Fo�?��>>��9�L�N����;�Q�ٽ\?��0?�Y
?b�>o	��1¿�6Ѿ�<�����f�����)n���ފ>��>�o���X���x>���>n	�>�M�>�^e>� ����=~�>�,�>���=�>O.=r�<�=}� >2�=��$=�i=n8(=�V��t<pL�,���L�@=_,F��>�����=C�>TQ�=:'�>b�<�A˾�<E��d��+�b�<���`S��1��ɼ����5���n��t=�x�>$��<x�����?�=�1�>l8�?ad?r�>l��<��׾�t��R3]�V��Ыֺ��X>P�6�.I��KM��k����?��>��>e��>32>�S:���=�O u��w�����r�>����]��d�������.��f��*c���>aL?����L>�W~?L�P?�7�?g՗>��{��qƾ�;�=���
̂�5Y$��?��gN����(?��?&=�>�����%[���Ǿ|ap�D��>tWj�Y�B�q��uJ4�|��<(��Q��>�b���Ծ$_=��ሿɲ����D���v�(��>�yN?p�?�h���f�`iN��E���&�4?jyf?���>�?��?YQ��q��;Y����=h?�s�?�?��=���=�d�t��>�?�H�?�!�?�jw?��6���>���<>�㪽�4�=�)>�=���=�?��?3'?d{���������:�쾯n\��g�;�̇=�F�>3��>+�`>_��=��v=���=��f>���>�u�>o�^>�U�>V�>WP��J���W�?[��)�>�-?�T>Λ^>B
G=j�P>��{�*��gj�Ju��NှL1$���u=�̉>��=4��>>�ӿ�g�?{��>�����)?)������	��-�=�o/�TI�>�ó>�K>�v�>)�>>+)>�*�>c_����Ѿ��>b���b#�֠H���M�X�Ѿ�\�>%ɘ��*B���ҁ���L�O'����Xj����� @�˲�<'Ր?.�潬�j��)�q[���?ԫ�>x�1?)���S����,>k��>��>3=��k��v������,"�?���?c#s>n�>yod?��9?Eh�}����`@�hՈ�4o��zf�=�t�b���:y�p�)�@�m�]T?(.e?lH?���=X�O>���?��ոԾl0�>�0��Q��K>56�>���9��������������=Οh?SOs?��?��7��җ=׶��n�R?�;?3�?"�T?��G?�=�����>�"?W�?�\w>��? �X?�x?��>�k�>	��������sY����&�K|��ʃ��>�)�;ʽ�����Ȃ=�"<א�;N��<������di^=�e�y�=��6>��>)�]?���>gO�>��7?���,8�l歾��.?F9=������G���I��v�>m%k?�ͫ?khZ?Hc>��A��B�b�>���>)'>
/\>�}�>�y��qD�wu�=��>>��=oN�������	�ȩ��@��<�Z>Z��>p0|>K��@�'>�x��.z�O�d>��Q��ʺ���S�B�G���1���v��Z�>�K?*�?)��=/^�+2���Hf�r/)? ^<?�NM?��?��=��۾�9�>�J��<�)�>xM�<�������#���:��?�:~�s>4���T��0a>��h޾vko��QJ�&��QMX=���x=K=f����վ	~�yz�=L{>I;��� !�4B���򪿓�J?�Fn=վ��G�T�U����>[�>W]�>�_@�N}�u�?��9����=�s�>�<>(���^K�{�G��'��ϝ>i8>?L�K?�*�?������E�o̠�1��������<C?E��>���>�>=��n=RE�����Yj�X{Y�=�?^��>�M��=�zP�<�$��s��I=_�>�A�>��\?��?ldl?v��?�%?s&?l�?��i���4�:?(/{?���L��kϾg�c�R�}�Δ?��F?�
�z-?dGd?�GI?\�?��`?�N'?&�>�YH��ڏ�RU\>��4>RL\�\N�����>��;?���>�".?�e?e�=�dE�/���ʇ5�w��<�Qz>�I?�?d�?o�>���>��u����=n�E>7�u?|�?�ߊ?/�>t�?���>�gq>�>�_�>_X?3�?�H?�Zp?  ?��h>=΢<=�I=h�	��򮽅�C�_��=�iA>i�=;�=�Rh�C&!;���;oȞ=��\<" �=�,=���=���=�V�=LI�>	]t>�+���0>�ľ�È��zA>�Q��Q~���i���H:�SA�=�1�>�o?Rc�>a%�֋�=�>���>j�T(?$?�?��9�]b��ھ/K�9&�>�9B?{��=�<k��6����u�se=��m?oe^?�2X�o��A?c?�]?N��k�7�԰˾�/��>�����N?d�
?ewM�`��>�"�?Fur?�D�>�kZ�'{h������Af�	����"�=+H�>����k�Ny�>D�7?�W�>$�v>��>����w��N����?^�?�x�?p��?+A>�np���߿أ߾{M��?�b?am?i���T:?�*�={%�.�������K����Ⱦ,T��1���?侦@S�����Jh4��}>19	?��u?�X?�Յ?j���]b���M��B����w�t�Ga0�dP���N�S�9���l���xR�$����"�=-�~�WA�bx�?�(?I�/���>I�f��L�̾w?>����ݡ��Y�=[�����==t�X=�6i��0�Mp��� ?嫹>��>j�<?��[��w>�n�1�B8�͇���x4>�0�>��>#��>M;�;�>-��轰Ⱦt��(sֽ]c>	�b?�S?9�?��׽���ׄj����֬��ؽ	��w>�A0�E�š
�8[�z�"���H�����׾`/u���턼=�??�hf>�c�=�_�?ܹf?�Q�ˢ�����^���A>Q�A>�ad?���>�a$>�й��!�Fd�>�m?���>��>\����>��x{��T��� �>R��>J� ?��`>��K�rv^���������G9����=�f?A��mc���~>uT?,�+��T�:�C�>T�$���=��3V#���>�O?��z=��B>�R¾��	�^Az��:���'?�?�P���o&��b�>��?���>9�>�?�j�>������5=�z?ka?n8N?��G?�\�>&Xj=��Ͻ�u½��!���=�>��a>[�=q�>$��yY�2�׶K=�q�=�uY��dX�Og�<8�:Nm9��-O=�R>θܿn�W�%�߾�o���Ң���l��� �+���D.���ؾh���r�t��Z��@�<l'���u�����_����?���?�����A��:���䌿��qQ?�d��S��{�Խ� ]��ʽ����i�'���t��+��7��Y�!?v-ľ�o׿"�����3�\�T?<<?�w?�bd�;> ��処����I�8���о�����ܿ�ǔ���u?LV?�W������=��?�>s��>tu�͐�!|>*�>�z�>'�?���=(a�-|ɿ�H�<��?�v@N}A?�(�����U=��>ߎ	?)�?>�N1��F�����U�>�<�?��?�M= �W�!�	��e?�a<��F���ݻu�=�:�=S?=G��6�J>V�>7���TA��-ܽ��4>7څ>��"�����^����<��]>��ս,��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=�n��Pο<�$���%��^\<_b=u�߻�D�������W�侚����)#���=��&>�:r>K��>�y>�R>_?9sv?kA�>~�>:��b���w�ؾ$��=��l�����4�F�\�"��ˊ�����u2۾���R�3��3�M~޾@�C��z<M�X�}݈��ZS��p�3�@�WA?�\M=$A��.�2��Ҽ�|���%;^�a=�ix�j龨0G�KC~��k�?��E?������7�B�(�ZH�����ub?"�?�>��|���>�}��짽���>
K �D'��4S�Z�Z��`>?��"?vy޾?�����=5���ݑ���*?g�?��<��>�V?Z9B���=��>�ʾ>+��>±>���t��R��yQ:?��x?Y����qu��>��ʾ���S�f>�Q�=+�t�:e_�6e�> �f=Fr��J��n�G���>d(W?���>��)��ja��� �fV==��x?�?.�>_{k?��B?�٤<�g��@�S���	dw=��W?�)i?��>T����о6�����5?��e?��N>Gch�f����.�U��$?��n?%_?�}���v}�a��0���n6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?s�;<��U��=�;?l\�> �O��>ƾ�z������3�q=�"�>���ev����R,�f�8?ݠ�?���>���������=�M���ܩ?���?	��2�==\��c~����%���`ټ�N�鹯����F�E���̾9(�" ����=��y>�J@�F�����>ڝ1�S'���Ϳp:��i���l���?�ɋ>s�e�%����|]���j��;���(����QO�>	�>����4���'�{�5t;�������>.����>"�S����<���(�5<��>@��>���>cB���뽾ę?_��?ο2���ҝ�w�X?�f�?�n�?(t?�9<��v�#y{�<��e.G?�s?Z?>=%�G]���7�<g?A��$���w=���&E�U�>�@?�Ev>�xM��ا>s>ɽ-1>.>����ҿӼ���$���?(�?Q(ھx�
?J��?� /?���9���|�]���y>�O?�������~5���k�ySk��vJ?�%7?@s�<j/=�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?  �>r�?�i�=I]�>�b�=�ﰾZ�,�pt#>�J�=��>���?��M?�G�>�H�=i�8�I/�AXF��CR�y ���C�F�>��a?SL?KAb>����2��	!�<@ͽ�a1�K��.F@�̦,���߽""5>-�=>�>:�D��	Ӿ/�?N��ؿZx����'��64?��>!�?0��bgt�Kr�_?j��>���1��6�������?I�?X�?r�׾b�ɼX�>S�>o�>&�Խ�����O���U8>�dB?E�f0��5�o���>s��?��@Lۮ?�h��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?pQo���i�B>��?"������L��f?�
@u@a�^?*C���A���Ӿ�6ž�?>�!C>�i>!.�Dc�=��'�B5G��f(=M�)>gn_>z$1>��s>�,">��r>S/a>H��T%��ɛ����.84����@W����' �O6;b�%��ؒ� �þ�3J��
����,�S���|�8?>�TS?ȓS?�Zr?�f?�B���.">c ��`�<#����5�=�3�>B�/?3�P?�-?���=Τ����a��k���⨾�Ӆ�c�>fmX>��>�=�>0�>Y:���,>XY8>P�x>��
>�)|=(����J)=bfD>�;�>���>o3�>7 �=Z��=����[����f��m���1��V�?7#پ�Ha��Fk����������M_:?q��=T�����ֿ_���]?�����1�:6B��>��d?v�:?��>�!�l���8�y>��i��m�=���&�,ON�ݟh>��N?!�f>�u>њ3�^d8�$�P�"|�� i|>n46?�涾�D9���u��H�Kcݾ4CM>�¾>)D�uk�������ti�_�{=$x:?ȃ?�<���ⰾ�u�C���UR><\>�m=Ow�=OZM>q[c��ƽ 
H�Pq.=9��=ެ^>��>k�?>佀=
0�>�\��J��1�>#`[>��]>0�B?$'&?�H�&���9���nJ�NQ>��>��>>�>�'9�*��=ٸ?�eI>�p�B�c�
��>T��=�>xM�� �.�l��l�T=𷮽��=�}�=��뽭D���=�~?���*䈿��e���lD?W+?^ �=��F<��"�B ���H��E�?q�@m�?��	��V�C�?�@�?��B��=}�>�֫>�ξ+�L��?��Ž.Ǣ�Ô	�D)#�hS�?��?R�/�]ʋ�7l��6>�^%?��Ӿ��>�g>��t������w��0�=��>�`C?aP�n�i������>���>��辢R��xLοY�k�>�
�?�?��j�Å��4�G�=�?���?�|g?{@>����p�;�E>x6?%W?7�>y:�.��?ϼ?�Մ?��>WJ�?��?�H�>|��=�Ͼ\���%��9��l�3��=;=EЩ���u��"D�{5���6j���O�ʻ��~�>�YM=,�>{������؝t=-m�<_b�������j�>�A�=J'�>ǎ�>��=�	.>�r�>��:�U8��l������(M?~-�?���ۅp�ƃ<�)+=z:��;?�Z9?gm!��!���¸>Ys_?�u{?vC[?$��>q��0:���R��Tծ��sm<�A>vs�>N0�>�1����Q>�ҾܨG����>s��>��i��ݾ�pd����آ>�?�\�>��=× ?��#?��j>�&�>|_E��8��o�E�״�>���>�I?��~?$�?�ӹ�{Z3�����桿�[��=N>_�x?zU?W˕>I���/�����E��GI�����1��?xg?�H�]?3�?��??�A?5&f>����ؾn�����>�!?���y�A�<>&�RW��?S]?s�>�ܑ���ս�ռa�����1?�$\?�F&?�T�ka�þ�e�<���(X�W�;F�&�>D�>r߈�c�=�H>ѭ�=�*m��36���h<�@�=ig�>S=�=�6�L!��)5,?C�I�0݃��T�=M�r���D��.>��K>����,�^?j>���{���������U��ʍ?`�?��?��/�h��A=?y �?�8?(I�>�Q���޾Eྣw��>y��^�K�>r�>�c�%u�F{��$����D��JPƽ��Y����>z�>BX�>�8�>��+>ڍ�>*-I;k�ٹ�`����k�1O��6@�C5.��+� Ͼ�Z�x�=N�U+��lq>Jk����>�y�>��>��>|c?��=�h�>�x�>
��>�ѣ>�\>�In>s�>��˽�@���KR?����/�'���辺���j3B?�qd?N1�>Hi�3������x�?���?Qs�?�<v>h��,+��n?�>�>>��Qq
?�T:=e;�j<�<,V��K��`3��x�B��>lE׽� :��M�nf�Xj
?�/?����̾�;׽����?��=\�?��2?Z�#��G��a��e�o�S�g���\
������c+�#o��$��S%���&��l�=��?pg�?ي�+��_�.Am���O�S>-��>�Ϝ>��>� +>Ǐ�z,3�P�M���!�;�]��K ?�m?�e�>C�*?�5?�d?�^S?H8n=
�>�-�����>�z�>�>��G?�o"?��^?"�I?p�A?�b5?]A�=z�\���c��i�)?78#?�&?�}�>�}�>�᤾��S�P]=D����*��AD=]�?�����ҏ�lPl=��^=��*>qW?���_�8������k>"�7?���>���>����%�����<U�>ٵ
?xF�>4����yr�c_��W�>*��?���Y�=g�)>X��=�����Һ\�= ��� 
�=�9��No;�,f<�|�=\��=�&s���t����:�Ї;�j�<	t�>R�?Z��>�ǈ>1����S �,@�)�=��Y>7�T>��>�Uپ�B��� ��i�g��w>8�?�S�?��l=#}�=>"�=<4���^��.���nS�<e?M}$?hpT?�Ȓ?�x>?/#?8>z�C撿����=��K~?�!,?���>7��,�ʾ���3�8�?'[?�<a����Y;)�O�¾��Խ�>:\/�0~����D�"u��m���~����?p��?�A���6��w辽����Z����C?F �>�X�>��>l�)��g��$�i3;>)��>R?vB�>�O?kI{?�\?�W>n}8�j�������l�?�s$>s�??�܁?D̎?Hy?8V�>�c>�[&���߾�7���d!��T�������^Y=l�Y>�ɑ>Nz�>ǩ>�v�=��Ƚ�ҳ�	�?���=�a>�^�>!ʤ>��>x>0�<� H?(�>���w�������n��7�E�+�u?|��?J�*?�==����D�����o��>�o�?<�?n�)?\�U�<j�=�k׼Q���{@r�2H�>G�>�G�>t��=G0D=�>���>{�>������*8�N(G��q?�_F?���=��ſ�q��p�q˗�J�d<����A�d��[����Z���=s�����ȩ��\�\ˠ�Ϛ���굾I���#�{�^��>
��=!e�=
��=��<�Fɼz��<�>J=!�<
�=��n��2r<
9�]xһ���Y���^<H I=gj��ej˾�~}?�1I?˜+?�C?4Ey>]�>_t/����>j���K?+kU>`T�9��Z�;�俨�dW��W�ؾ�.׾v�c�՟��		>�{K�Cg>�B3>��=�؊<+��={lp=�p�=8D7�[=���=א�=�j�=��=��>�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/> �>>�	>՞S�q�2�� ^�{Pj�p8d�^�!?q6�ǭ;���>L��=�׾�vþ��K=gMA>w��=6��_]�X̘=�h{���;=�$`=2~�>��?>3��=B���;��=�6="S�=��Q>�{+��J��k*��H=�`�=�k>Ћ0>��>�?�q1?Sg?�5�>��x�?�ɾ_?��@ǌ>dy�=P'�>�E�=.�M>�><H7?�gE?�aN?�ԯ>HHt=@8�>��>g`)��gn�&�꾺h���ܶ<!�?堇?���>��@<Y9V�"�)9�z
����?A.?)�?�Ø>������2}+���0��w��[��=��>�����T3���)��&۾8�ݽB�;=R��>� �>vB�>��>gۇ>nYg>	O�>l>�`{<g�ʓ̽���=$a�J� =^8$���<��xX��6����=��=,R=���<R��;�j��O�=���>�0�=&��>%�6��{߾��=Mp��AD�=�->�ϾiT�G[�",y��>��䕾"��<Pζ>��ѻ�����?ʈ&>��>0�?�^~?�^>�jb������v�	����L�=�*v>:�ɽFG4�JO��U�����$j�>S��>V*�>:�">[�4�"K�t��<�1�*��l?�֢�הǽ�3� y�h���T��ߚj�8��=v@? ŉ��W7>�K?�QT?�T�?��>o���;����#>���QY�<~t�~|������k"?�?��>����j�<�tp̾�e���J�>\RI�o�O�~���@0���g*��� �>������о�2�P����2�B���q�'=�>��O?ظ�?j�`���i.O�x����?>?�)g?*V�>��?)�?��#�ր�LI�=L�n?z��?.��?|>R��=�g��C��>d�?}��?���?% t?�"9��*�>q <3�>-���T{�=.�>)��=]�=�?�n
?�	?����n �V���P]�(�=r�=>ڑ>,�>j�u>��=��=�]�=)
[>J>�>�Ȑ>|h>=]�>Ŋ>0Ȩ��wݾ� ?�c</tp>�5?�ѓ>�߇=$ȉ>���=���=8Z7���-�6l.�'��^z���<���=�=@��>[ɿ���?uY�>V{��*?^��#a��o�(>z�����l�9�>��A>���> �>��>���=Pܼ=�@>� Ӿs�>�'��c!�0�C��ER���Ѿ{'|>oS��m�'�L�����uI�G������i��M����=����<�T�?�-����k���)�����A	?%�>^�5?f���	w��y[>�^�>U�>kF�� ����0���,⾲�?�(�?\qY>w�>\\?P?I.�!14���T�Ĉ}���C�:�b�#!c��ڍ�L킿�3���eR?Q�m?L=?Y��= �l>_P�?.�c���K�>�@/�B�G��{'=�>*;��^K��.Ҿ�;Ծ��%�xO>��g?WE�?vi?��O�Vs�=��=c�.?I# ?8#s?Q��>1?c��R?Z+?."�>="?5	Q?��^?��!?Э�>+��>'���X�8��%_��pp�2���Z�^�� *>��=\G�=)�=PN<Sӕ�s8��T� Cؼ@���$퉽gni�t�=ԝ=xǦ>Â]?�D�>���>��7?�P��P8� ���!+/?==$h��ڕ��7?���t�\x>��j?���?2Z?��c>��A���B��
>��>��%>t�[>	N�>k��.�D���=&E>��>�a�=OL�!�����	��������<�>'��>�0|>m
���'> |��1z�8�d>t�Q��˺���S�A�G���1���v�8Z�>��K?��?h��=+_龈+��If�d0)?4^<?�NM?��?�=��۾��9��J�	=���>hJ�<�������#��p�:���:��s>�1��`����[b>Z��5޾w�n�� J��~�1�N=?��t#T=��N־�T����=-�	>ȣ��� ��"��eت��!J?^qi=2M����T�쉺�{_>���>x�>�g9��Nu��m@�k��� J�=���>k�;>������qG��V����>�w%?��>?3�?*���b{�N��f,�G���R|Z?!�=�?�T�>�:I>�S^�*��w~�G
t���>�|�>>_/��SA�J���2�7�4�n�4	k>Im4?��>�-?�۝?�+4?��j?�$�?�?���>��[>����9?A��?��B�^�m�پ��u��@��՝G?���>����$c5?0fn?s?�O3?e/|?��B?���>{�þ�S�1��>䚲>�@=�=x��"��>��+?��>0(V?xo?�+>#f��p��DR�)f��h=w�9?a	?�-,?�,�>@<�>���2�C=�Q�>��l?�^�?�?���=�/�>���>�2�>����՝�>�-?��?�[,?]�h?�p ?��>!�=.񑽔\t�[�/���ż�n���gq�|ܛ=4>��B=�#q�
P#;�-�̌U�XĎ=�n�;:�s=JNd=Lh�=�`�>��s>�
���0>��ľ�P����@>i����K���֊���:�ܷ=ƀ�>G�?Ŧ�>%X#�	��=>#L�>����7(?��??�c";�b�e�ھd�K��>2B?���=E�l�����F�u�c h=y�m?�^?��W�'+��K�b?��]?5h��=��þy�b����b�O?#�
?j�G��>��~?V�q?I��>�e�$:n�'��Db��j�Ѷ=Er�>IX�G�d��?�>b�7?�N�>��b> %�=cu۾�w��q��n?��?�?���?+*>��n�\4��`ž���-Dl?��>p1�y�)?K�=��.r��r��d���ﾾ�ݖ�I����ι����M�{�ǫ.<��=�N?Wo?a�t?7ƍ?n��\(x����j���'h�Y/�BmF��O�1�%���:��mk��<��4���������=�{��C��?��&?5<4���>Y]���S�
�̾XfD>iS��N/��	�=Rh��/�.=��,=�f��Z �`���&�?���>��>%�??�G\��`<�C�-�p�:�i���(>:�>R��>���>;w���(��3�Ӆ̾���޽���>*c?^P=?䉂?m�@�^
��OG��&�c޾7}�%��>罧�$���������og7��~C��ɀ�y ��=��.I!�����3?�w�>�yB>���?tDd?����uE/�Z�t��>�o?�U�?b-?�>�▾ya]�E��>!�l?���>ચ>Mˌ�.����z�Q�Ͻ��>�´>O'�>~�e>��J�خ^�Jŏ�������6�~��=�]f?��~�w�k��Z�>uN?�F��:t�<�@�>F"���"�CC꾶����>�?S��= D>h:��wK�Q
t������,?��?�?��4�*��Y�>��?c��>�ٻ>֌�?<�>9w¾t�a=��?�T?F=M?c�K?��>�K�=�}��,ƽ&(��g=`�>�c>\v[=|�>x,1��G�	��7�<�j�=�jJ��H佟|�;�=ٻ�/�>��<5B>��ؿ��E�#Gھp(�����Cp�JH�d���U��%t��-���8��;ｿ�@�OQ�۴O�N����7P���?b��?+BѾ1���%���|(q�����68�>�@�1�,������,�q�x����\9�����)o��!n��]���? ��pԿ�颿q�4���O?O&
?:i?z�<xp�����ՃA>�)=��ǽ;��~���j�DI����?�z?�;��&9��u�>ֆ�>P!�>�-�>�G����#4<=�O�>�/?9S?���(ܿRw���R�;v��??�@�|A?��(�����$V=���>��	?��?>rU1��I������T�>f<�?���?d�M=��W���	��e?s�<U�F���ݻ:�=�C�=F=X����J>�U�>U���XA�/BܽK�4>{ׅ>�m"�	����^����<y�]><�ս�8��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=����Ŀ$!�4\(���g����	ս\��s<%3<u6��Lz��b�ܼ��=���=�KS>r(�>$�*>��d>�W?l@j?��>ƴ�=��5��&��v#ھ�<��.��2��y{���`���A����6���	�Ӄ�!����0�A��̈=6�^�����$(-���S���-��_=?Az�>�<龈iP�LK��S���x��x� ���p�.l>�18S���?99O?����l�Q��3�~A5=�A��SM?��n�i�+�G����r�=����c�>�"�1�P��D��g>��A?�
>?=�׾���8>�E�_�b>�>?�?�s�<��l>�8l?�ŝ�.;�HK�>G
?0ӣ>W�?k�|�	k��%G��)?71l? *�τ��_�>��%U;��o���<@>8��Ks��m��>2Û�w���?ܵ=�����ɼ�(W?���>4�)����]���:��F==�x?~�?�/�>Ywk?��B?6ݤ<Ih����S����qw=H�W?�$i?��>⑁��о����5?�e?��N><gh�����.�fV�%%?��n?�Y?�w��?q}�������m6?��v?�r^�is�������V�8=�>q[�>���>��9��k�>ב>?�#��G������Y4�Þ?s�@���?"�;<!"����=�;?�\�>˫O�6?ƾ�z������m�q=�"�>L����ev�����Q,���8?Ϡ�?_��>�������>r �����?�Փ?��ݾק���߾�	���������A*����"�j�O�*i��{A�r��'v �)V��]s�<G�>.�@ V�s�>-�h��D鿃�ÿ򽅿M���P���Y?V�o>���<��`�n���1�)%���Q���/�M�>��>��������{�wp;� 3����>,,���>ױS�5+��i���+F5<�>1��>���>~@��<齾iÙ?�b���<ο��������X?�f�?oo�?q?Iu:<��v���{��j�R.G?\�s?Z?A%�V<]�8��_n?�����`v�d�Z�E1X�5��>��z>��p>;ʾ:�=zHB�s�>X����@e�ȿ�������Jֻ?���?�쾝J?`+�?;c?��"�����IBվT�8��,>��L?��<������k���T�ܛ��r�4?�#N?�ƽjS�]�_?+�a�N�p���-���ƽ�ۡ>��0��e\�N�����Xe����@y����?N^�?i�?Ե�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>	�}?y$�>��?]o�=b�>)e�=��@�,�Nk#>�"�=��>��?��M?�K�>5X�=��8�;/��ZF��GR�v$�5�C���>��a?�L?�Kb>e��4!2��!�]vͽ�c1��L鼺W@���,�q�߽(5>C�=>%>��D��Ӿ�[,?h�$���Ɲ�NqA��UD?�s>��>�B��ۈ���w�f?o�>���=���}���l̾�6�?��@a?��Ѿ��;��>	��>I״=Ͼ�����X�=�>g)#?b�N��ō��ٗ�4�>u��?���?�?ՎS�'	?x�BM���a~�����6����=�7?��{>���>��=�mv������s�Z��>�=�?px�?|��>�l?p�o��B��2=�3�>�k?�t?#k����B>��?���6��H��f?B�
@�s@X�^?(좿��ݿ:����W���hݾR�=��=�);>j�b�V>q��=����Ͻ�۹=�3�>\Jj>1\>���=�;>�g">�@��t�!������!��6�R�?2�����s����o|���'���־�À�۝Խh2Ľ�N��sX˽�˓�4�=>?BT?^R?��o?�@?�L��&.>t��K��g�B�5�I>c��>uXI?�O?G~??��G>�u�z�h�)����V���BS��>/��<�C�>�>0*d>J9=�9W>W;>`�h> 8��#��<�ܐ�ɑ�c�>�y�>���> ��>�)>n�+>h���C��	�v��i�m�ݽۢ?Hx���FY����������h��9k;=��'?燿=�Y��pmп=@����S?k��Y �rD��(2=��@?�C?4u>��Mb�2w>ϥ���^��	)I=0k&�I����L�lEV><#?9�f>�u>!�3�d8�&�P�h|���k|>46?T붾�F9���u���H��cݾIHM>ľ>I
D��k�����=�7ui�u�{=Yx:?	�?�;���㰾��u��A���RR>=\>7Z=�k�=\M>�Qc�a�ƽ,
H��m.=s��=]�^>h%?z,>E�=j��>}ᙾs�O��K�>��C>��->�>@?��$?����\�����S.��_v>�2�>2��>]=>��I�Q��=SJ�>}b>�?	�N����@�D�>�6V>�ux���]�}�p�[a=�ܘ����=>p�=����I<��A"=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�h�>��۽������n~��P>���>5NB?�l�=�b���'�z�
?�f?&��Fܧ�N{п<E���4�> Y�?�q�?�u�K`��q 7���?��?D_?Q�>�ľa��GL�=�$J?\�a?cd�>��=�;cG��?��??�?�΂>p��?���?H�?��0=X��W,���4��!����A=�if>�����J�8NS����5���WE;���'�Y �>uO�<��S>�;�>Պ����m >��|��4ڽƔ�>���>��>�>�!Q>h��>5�p>˷��P����}��-����K?���?���1n��:�<d��=2�^�|(?�H4?ގ[���Ͼ+ڨ>��\?���?�[?�g�>S��=���翿�|��E��< �K>�1�>�J�>4���LK>}�Ծ�/D��q�>:ɗ>���?ھ�0��R�B�>d!?8��>�Ӯ=*P ?O�#?OQi>�v�>�D����$F�9��>ȏ�>�?�Y~?��?6ܺ���3�l���ۡ�$t[���N>�x?�+?[x�>o;���{����`�kG��2��&��?pg?ͶݽV�?�G�?�??�+A?$�e>�����־H	��룀>��!?aT�M�A�06&�8���?�_?���>�>��{ս8+ռ����F���	?3#\?	=&?��#a�4þ�2�<@G!�"`N�|E�;�`C�2)>h�>�H�����=��>�߰=7m�E�6�O b<G��=-Q�>�.�=�[7�I����8,?�'�Wh���~�=cxs�qD��Du>Y*E>*x��x�^?�E��^{����Jל��+Y�c,�?'+�?q�?Lg��4xi�:>?�?�?Ul�>/;���ݾ��޾"{�j�}�i�����=�Y�>ڱ0��������0��1X��Zuڽ�R��a
?���>.�>q
?>[��=Ϛ���^����Ek$�P|p���W��K���A��$��߮��#�����=`�Ⱦ
Lo��d\>���|�>��?��o>�;�>�O?�M>և�>C��>p�>-��>H��=$�=G�)>̖�������KR?����|�'��辸����3B?�qd?1�>�i�<��������?���?9s�?�:v>ch�/-+��n?�?�>����p
?�R:=�9��@�<�V�����43�������>EF׽� :�zM�of�<j
?�/?����̾:׽|t��KCp=�P�?�)?i�)���Q�$�o��W�a&S��@�h������$���p��U��H��e�(���*=�}*?+!�?����X謾<k�?�ff>j��>��>;��>ՀI>	�	�R�1�z�]��@'�X����=�>AN{?��>A�2?��4?�W?��c?�p��,��>�O��wR�>kt��>��#?�0?W�??v�S?�I$?��U?�]O>p�������о.(?�;	?�c?A�%?�>�����9�d��=��'����������k>�[5�k־�s�����^�:=@X?m��S�8������k>��7?ޅ�>���>����&��p�<N
�>��
?�K�>
����xr��\�$O�>c��?u ���=V�)>!��=?����̺�O�=�=¼��=3����;��d<���=��=~v�m*�����:��;�<��>��?��h> �d>�rf���������=�(�>I!M>ב�=�����t��9l�i>>���?�?E��=i��=({�=R���Ͼ��������=�W
?��$?��i?��?�vG?�1?n��=������p��Ҏ�@�?i!,?��>�����ʾ��ȉ3�Ν?t[?�<a����;)�	�¾��Խ��>�[/�Z/~����:D��򅻬�����/��?࿝?$A�P�6��x������[����C?""�>9Y�>��>7�)�J�g�S%��1;>��>?R?a5�>}�O?��y?	�[?o>��7��릿�����&J�c>�PC?`�?b�?�^x?�7�>&�>>�!��u�����y;8�L.�tRo�bU,<�F>��>	:�>ŕ�>���=ٻ�귽:]�Q�=f�M>�&�>���>��>��q>�|�=�jK?���>�l;�j��Y���5���A�� �?�?�9$?�,$=�:���>;�0�i�>鞪?d�?L�1?�|����=a�	�ԥ��u�B0�>�ٷ>���>��4=�~�=�A>ܞ�>+8�>)��^!�K�5�C괻a ?�M?I��=	2ȿ��r�Qqk��Y����(<�����i�|����8�a2�=�x��bG��L���V����I���0������%ix���>d�=S>*��=D�<�A�u\C=��='=�1= !u����M�E�n<UÆ������:"kP=�%T��}˾�}?DI?{�+?:�C?�y>�e>�\3����>3���@?n�U>-�P�dj���m;�ʩ�����	�ؾ��׾G�c��ß��R>.I���>�G3>���=縇<�?�=ccs=���=TL��^=�<�=��=^�=���=��>�'>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/> �:>n>��R��1�|3[�df�e�Z���"?R�9�4˾2z�>��=~�ݾ�=ƾ�!==}J<>VSg=O���\\����=i�}��&@==�h=k�>��C>��=sU��=�=��R=��=�P>,�j	H�^K.�)�==�)�=�od>I'>�D�>?41?�c?��>�r��;�oƾ]��>�=��>���=�Q>�n�>}�9?��F?x�L?�*�>��Z=�>�͢>DB)��m����&Z���v<H��?Fo�?��>>��9�L�N����;�Q�ٽ\?��0?�Y
?b�>o	��1¿�6Ѿ�<�����f�����)n���ފ>��>�o���X���x>���>n	�>�M�>�^e>� ����=~�>�,�>���=�>O.=r�<�=}� >2�=��$=�i=n8(=�V��t<pL�,���L�@=_,F��>�����=C�>TQ�=:'�>b�<�A˾�<E��d��+�b�<���`S��1��ɼ����5���n��t=�x�>$��<x�����?�=�1�>l8�?ad?r�>l��<��׾�t��R3]�V��Ыֺ��X>P�6�.I��KM��k����?��>��>e��>32>�S:���=�O u��w�����r�>����]��d�������.��f��*c���>aL?����L>�W~?L�P?�7�?g՗>��{��qƾ�;�=���
̂�5Y$��?��gN����(?��?&=�>�����%[���Ǿ|ap�D��>tWj�Y�B�q��uJ4�|��<(��Q��>�b���Ծ$_=��ሿɲ����D���v�(��>�yN?p�?�h���f�`iN��E���&�4?jyf?���>�?��?YQ��q��;Y����=h?�s�?�?��=���=�d�t��>�?�H�?�!�?�jw?��6���>���<>�㪽�4�=�)>�=���=�?��?3'?d{���������:�쾯n\��g�;�̇=�F�>3��>+�`>_��=��v=���=��f>���>�u�>o�^>�U�>V�>WP��J���W�?[��)�>�-?�T>Λ^>B
G=j�P>��{�*��gj�Ju��NှL1$���u=�̉>��=4��>>�ӿ�g�?{��>�����)?)������	��-�=�o/�TI�>�ó>�K>�v�>)�>>+)>�*�>c_����Ѿ��>b���b#�֠H���M�X�Ѿ�\�>%ɘ��*B���ҁ���L�O'����Xj����� @�˲�<'Ր?.�潬�j��)�q[���?ԫ�>x�1?)���S����,>k��>��>3=��k��v������,"�?���?c#s>n�>yod?��9?Eh�}����`@�hՈ�4o��zf�=�t�b���:y�p�)�@�m�]T?(.e?lH?���=X�O>���?��ոԾl0�>�0��Q��K>56�>���9��������������=Οh?SOs?��?��7��җ=׶��n�R?�;?3�?"�T?��G?�=�����>�"?W�?�\w>��? �X?�x?��>�k�>	��������sY����&�K|��ʃ��>�)�;ʽ�����Ȃ=�"<א�;N��<������di^=�e�y�=��6>��>)�]?���>gO�>��7?���,8�l歾��.?F9=������G���I��v�>m%k?�ͫ?khZ?Hc>��A��B�b�>���>)'>
/\>�}�>�y��qD�wu�=��>>��=oN�������	�ȩ��@��<�Z>Z��>p0|>K��@�'>�x��.z�O�d>��Q��ʺ���S�B�G���1���v��Z�>�K?*�?)��=/^�+2���Hf�r/)? ^<?�NM?��?��=��۾�9�>�J��<�)�>xM�<�������#���:��?�:~�s>4����\�]>3��co޾~�s� �H�+"��t�=�����<n��,AӾbfv����=�&>�����"��A��.���N?�!�=*����T���þ[9%>C��>��>.���{{�t�>��C���9�=��>Z6?>�� ����k�G�Л��	�>gB1?�_R?�\�?�K����C�B�;�%������K�=� ?_ڥ>kw?�	t>���=�¾���F}c��a�z?#�>G�#��H����u��z6�J��>/�D? ,�� a?�ە?��?�ʗ?ݬh?�9�>��
?�ݪ�^!�, 9?>�q?:����X���,ƾ��Q�����b6?%�V?�P �~p2?��W?LB.?c^?�w?I�?�s�>��꾢�m��~�>��s>aJ_��ͩ����>�X	?�*�>� O?5�|?��<����dͽ��=j���{�&>�Cn?I�F?��?���>Y��>�G^�\�->txF>
�l?��?~�?gPa=51�>X�d>L�>M>�>?_?�mL?�^y?ǜC?���>�Ǧ;�Hҽ]�+�����Ѯ<��=&D�=��=	տ���J��Pl����=��;<@^żsjf��Yý�8 ��ؼ�xb<z��>S�p>�-���@/>O�¾8��:A>Dć��+��Ql���=9�j�=@�~>D ?�ˑ>?D%�$˔=*N�>�C�>����'?ݾ?�o?�8�c�lܾ��H�4�>�C?r��=��j�殓�]�v�=�e=Gl?�]]?��V�����a�b?��]?�f�=��þ��b����5�O?��
?�G�_��>��~?��q?ӽ�>U�e�
9n�����Cb�5�j��ֶ=�q�>�Y���d��>�>*�7?!R�>a�b>:�=�{۾c�w�l��?4�?��?B��?3*>Z�n�43�2����~�_�H?�?����u=!?HfD�y���?�؝L�H^��O�����&0�p[�w�����O����=}^?Tj?�f?m_y?�����,��B��0��t{�Խ"���+� �V�)�F� �4��CY������kı�H�>�~��RA��n�?�(?͂/�0��>���������̾�lB>���"��9��=o���%9=ĀW=|`h��/�������?�ɺ>i��>�<?�>[�Q">��1���7�}��W�2>f��>>��>+��>KAo:Y#-�����ɾx݄��н�|>��^?�X?@�?��ҽ���z��$�Iac�ۀ�� �P>c�<@�=T�޾dps��y$��Q���w��<��䁾x����-���7?�
�>Xβ>�?�~�>���R�
ž&($��ֺ>�Z�>F_?�p?]rT>1�����~,�>��\?���>	�{>�}��?(�R����~�>l6�>���>Og>�U���>g�m���G��R�4���%>P�n?�
��m�_���:>�u?9��=��>00�>_�5�|�!�fa��Ib�Nx=�?G�X=�\h>����{پtF�������)?��?&���P0+�C~u>"?�	�>䠭>)k�?�ޏ>��^R
=)I?�:^?��K?ݏD?�W�>��N=�Bɽ�
Ž����=.�{>��f>{�M=A{�=�\#�n
\�p���n�<#y�=Z� O��:��ƼΡ��}b=�1;>X1׿;HL�vFӾ����p���2��
¾�Z��Aj��mN��k�\��㍄�����[!<JP����#릾��s��a�?W��?Ԏw�E@M�浩�����Ns�og?�p��|���W�0�\��<ҷ���ྺ���?B��Nv���v� ����?+?b�����׿''�����h[~?�?<��?�PI��p7�����X�a=/ֳ���;~ߴ�����q߿�2���r?�?����U�ʽ��>�?sq>�%�>�2־]m��R=>~7�>C�
?w�>̈́���e�hȫ�_˽���?�L@�yA?��(�����U=<��>�	?I�?>\1��7������Y�>�9�?���?P�M=��W�9�	���e?;�<��F���ݻ�?�=��=2�=����bJ>4@�>�}�LA�֣۽·4>C�>?�"�����u^���<�X]>�sս�5��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=��[�ÿ�8"�*E"���H=���=��L��m�����&<ށ��Xލ�ZmĽ�3�=QO>�}>ت�>��B>�+h>VIY?�1h?A��>��.>��=��夾���(w=�a���c�8>>���<,¾�_�n��f�2�D�6�t��k�2;��G=�KK�Q׈���B�G[�٠I� T=?x�=K��I$�~��<�1��p̏���1=�q����H��t���\�?�J?�����pA���1��4<*$����~?*�z�:Y	��p����P=�7�=|KE����>-������G=�7_c��)??�q9?��ܾ����P>9�����=�f=?^�J?d���վ�>�r?��=Qo3�R��>L�>%��>��*?�Ƚ�ݙ�����&?��\?_��=�lX�4��>�l��gU���y>`M�dB��Sν^�v:�	<�c��m+�k�{��y(=�4W?��>�*�h��}���9&��P;=��x?��?�=�>:�k?FUC?�5�<����.S�ބ
��=��W?��h?�>ѽ~�&�Ͼ�d��N�5?E$e?e�M>�/i���2L.�,���?�@n?W�?�*���?}�;;��T)�N>6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?k�;<��U��=�;?l\�>��O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>��������=+���Ǽ�?���?������!=���s�X �)u�&=���c���:���a=��Bɾ�?	������k;���>L@䀢�ϻ�>�����ݿ��˿𛃿��循^���?��>i�Ƚ�У��mb�
�i��#G���E��d�dQ�>��>$������{�xs;��럼��>6�����>g�S�0�������'8<$��>b��>յ�>kV������ę?,Y�� @ο񨞿Ü�H�X?�g�?hq�?Ms?��6<N�v�,r{�����+G?$�s?�Z?Z%�66]���7�~�l?�*��I�v��U�� +�x�;>�I ?��>��E�f=�p=�x�>�}^=@���0ʿu��I�4�+�?S�?��о9�?��?�'?,뾎p�������T�#��>t�??�ۼ5o��V�N�@3X�leӾ��1?�wc?��6�+^�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?$�>}�?�n�=na�>Mb�={𰾽	-��l#>)�=J�>�Ԡ?��M?�J�>TQ�=�8�|/�zZF�OGR��#���C���>�a?��L?�Gb>���(2��!��pͽb1��\��X@�d�,�E�߽�&5>��=>�>��D�Ӿ�?Cp�i�ؿ�i���o'�274?5��>�?g���t�|��F:_?{�>5��+��\&��@N�Ú�?�G�?��?��׾�#̼B>��>|C�>?�Խ�
��8~��!�7>��B?^�C��f�o���>B��?¶@�֮?i��	?���P��Va~����7�c��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?jQo���i�B>��?"������L��f?�
@u@a�^?*Q�ʿ�٣��M���yپb����>�q>^L+��A�+(�>��νnk�����>���>;{B>���>�nn>evk>̩S>15�s�+���<�����f����S������F�X�}��D@�U���ډ�Ј��e-r� }�=`�����t8�<� �=%�V?\V?>�r?��?#h����*>�g���<U=\����=O��>��9?HQ?Z�+?
��=ω��`�1���)���y���`�>(,)>���>���>.�>
�;�)T>un>>��>;{�=ND=N��;NJ�<۴f>ı�>e�>I��>[�->cw>���>\���:�����wU���?��ھ�~b�S|��������Τ<��/?�ͪ<i���d�ֿ���Lr_?�c�� =��LX����=M�a?g�R?Yp>��ؾ���<�>�{9�j�����P= J�n�����;�+�=>3�V?�f>��t>ݛ3��[8�ͼP�FZ��0n|>736?�ֶ�b9��u�רH�#ZݾD8M>n��>�{E��_����/�~��fi���{=�:?Bv?J䳽�����u��2��)�R>̌\>� =���=ySM>�rd��ƽ�H��Z.=��=�^>U��>!��=��[=�>p���_�����>�&y>�O�>xF?U?4����ƽ�S�� ���R>�F�>��V>s�'>F%����=&?�>!F%��^�ˬU�m
����>К1<��g��ս'�Ѽ!�l�gߒ=`;g��W�p�$��~?���(䈿��e���lD?S+?` �=��F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž5Ǣ�ɔ	�/)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�k�>�}��[�������u� $=��>�:H?^]����O�,�=�/t
?F??X�*���$�ȿ\�v�U��>h�?���?��m��>��V@�G��>���?WfY?�^i>a۾�QZ�6��>��@?[R?��>7A�B�'���?[�?ᮅ?2�o>�g�?��?��?G�<>�e�%���7:�� _��2�a��/>ޗ¾sa�Xg����ĭ|���F��k���>f�=E�>$E<�o��jr�4v�J��z`=��T>�bY>j��>�N�>�oL>rn�>P?�>]0����B�W|G�32��(�K?ڲ�?E��_2n����<c{�=;�^��*?6M4?k�\�ƷϾ�ߨ>ɼ\?9?�[?l�>J���;��翿�{����<��K>�*�>�J�>u3��%9K>9�Ծ2D��u�>�Ǘ>Fۣ�T=ھ4��T���A�>�`!?(��>��=ٙ ?��#?��j>�(�>8aE��9��`�E����>Ӣ�>�H?�~?��?�Թ��Z3�����桿��[�t;N>��x?V?qʕ>[���ო��jE��AI�����Y��?�tg?�S�*?52�?�??T�A?�)f>Ç�
ؾꩭ���>��!?����A�2L&����M?�P?%��>�8����սqSּ���=~����?3&\?@&?����*a���¾{3�<ӷ"�HT�t�;��D���>v�>���͜�=�>c�=Em��@6��f<	m�=�~�>�=�*7�+t�� =,?��G�\ۃ���=l�r�*xD��>�IL>�����^?�l=���{�����x���	U�� �?ߠ�?Gk�?����h��$=?�?�	?X"�>�J��~޾����Pw�M~x��w���>���>��l���3��������F����ŽD±����>�g�>�(*???���>¢�>����3�3�
较���Y��8���9�hT9��������w����=�ͫ��ݚ�5@R>Y��h��>5?N̿>l�>�>hO~=���>��>�5�>�?7��>@W5>���>�����.�@KR?����X�'����Ͱ���3B?Lqd?�1�>~i�����F���?��?�r�?�8v>w~h��++��m?�>�>���!q
?(o:=Ml�)�<�W��]���.��6�����>,;׽!:��M�yrf��i
?�.?^��c�̾9=׽#~��\́=��?��,?�}%�a�L��Bn��K[�GS���<�a�w�M¦���&���r��U��ht�����b)���d=��(?���?�d�������mk���>��c>|��>_͏>�M�>��6>p'��)0��Y���#�������>�|?�u�>�EP?a�B?YT\?��t?�u<�+�>�蟾��?!�>L�>i	4?+�R?��:?>QF?��F?�B?4�@>�٘��|�6־�k?c��>E��>bT?�y�>�w��CX�8җ=��a$���<���>[���Q��쳺c�����=J�?\��9� �����n>�A8?(��>��>���i�����<�}�>1�	?�N�>�y ���q�y^����>Ut�?�y�f�=��->!��=����-�b�em�=a���~��=?@�����~<:�=曓=Y�R�H��/;xQ�;
��<#t�>b�?���>�C�>�>��� �۵�6h�="Y>�S>�>�Eپ�}��.$����g��Yy>%w�?�y�?��f=�=��=�x��
V�����m������<��?sK#?YT?G��?%�=?�i#?��>�*��L��'^�����a�?�!,?x��>���V�ʾ���3�`�?x\?&=a����#:)�h�¾q�Խ�>�\/��0~�5���D�d������������?��?�A��6��w�ֿ��-W��הC?"�>�X�>��>��)�.�g��#�k7;>��>8R?�߻>�P?�{?��[?KY>u=8�7O��bH��@����#>ׯ??�ʁ?�5�?�y?56�>H�>N,%��ྔ���f� ����⺂��F=f�W>��>���>J��>��=��ƽ���6�C�Eߟ=�	b>�h�>�٦>���>[hu>KM�<ϑI?D��>^aǾV�� ���,��QJ�B�y?� �?��?�O�=`���4�?����>/o�?��?��(?�d�pJ�=⧨�l밾�z��>��>.�>T�:=4�B=>8>*�>���>����{�Z43�n�E�m9?�JK?�D�=C�ſ�q�q����݉f<YҒ��d������Z����=�Ƙ����#ũ�N�[�oà������ص�����O~{���>���=*�=���=a9�<Pʼ���<��J=ঐ<��=�]o��n<D�8��QԻ3���0v�L\<Q�I=:��,�˾��}?!=I?Q�+?F�C?�y>w)>Y�3�̑�>V���'=?�V>.�P�������;�Ӯ��I!����ؾ�p׾��c��Ɵ�{I>@}I�e�>�13>n5�=���<#�=]s=iێ=�Q�O=�,�=eI�=�Y�=F��=��>�F>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�9>�~>��R�W�1��|\��d��Z�/�!?<>:���̾I�>t,�=��ݾ��ž/�6=F.8>��j=�a�9D\�J��=)�v�/a==�l=/��>p�B>׈�=ᱽ���=�LP=���=<�O>Oݸ�7A�1n)��~3=7��=��d>8�%>.�>�c?�0?ed?w�>-On�so;���2�>Mt�=.{�>��=@�F>O}�>�8?�~E?�L?��>z��=o!�>ʥ>��,���m�D�\Ԧ�� �<��?���?HS�>�Bn<PJF�8��>��nĽE�?\0?��?�i�>��aR�#���h�ǲ���"=_��>�?��Ҟ��H�>-�1�ڦ��Q�>��>��>K�?�y�>|�>,�>��>3��>��8����=��/>6/="'>�P$<?�=�d�pS˽�y&��E��З�<V�=�<��=��ǈ1=Zm�=.��>���=�~�>�w�=���C�=�c��A@�ʹ=������C�:�c�������5��M��2>�YI>���f�����>r+#>9~�>'�?~N�?f�]>�}��]��I��us��GT���=�%2>��#���1��(M�RR��_־�x�>+��>�k�>��:>�"���C�nu�u�'\ ����>�����<W�8�u���������9c���A=<MK?�U��~��=(&k?�]?*��?;��>}�۽�ʾ%�>k��������8G�i���J?��!?�?�}��)B�bH̾M���޷>a@I��O���@�0�r��ͷ�,��>������оb$3��g�������B��Lr�(��>%�O?��?(:b��W��<UO����,)���q?�|g?x�>K?�@?�%���y�r���v�=��n?���?:=�? >>�=DDͽs��>�6?��?y�?�n?��/�)�>W��(>���)�=�?>$=1�=�
?^�?��?u��M��R�Ծ!�������ߢ<���=���>�i�>�y�>\v#>���=���=N�T>��>�]�>�f>w�>���>kĝ��j
�a?�#�=!�>|�6?���>�N�=/֐��K+=v�C�If8�l1'��Q�����-v;W�/<[�=�s;-�>0����B�?�Q)>�M��?c��9?��+��>���>��[����>��G>�d<>/��>���>2>-��>W>��Ҿ�M>�'��j!���C�sR�{�Ѿ�}>�H����'��X�L6��~�H������
��j�\C����=�J�<�T�?����l�	�)�����#	?�>'6?$2��jt���>Hq�>�>�-���m��aݍ���'��?]#�?�rc>���>/�W?Y�?�*,��F.�0�Y��3w��OA�0�d�Bwa��ٍ�Ɂ��t�B�ѽ/I]??�v?>?v�<Áy>�?\#��ޏ�7~�>�/�;�G�==�,�>n���^�T�վ��¾0����H>dyn?���?)?kM�򆌼��>-G?��?z��?��"?��L?L���!*?1��>��>i�?TG?� J?��?wY�>O�> z�<^^���O������� ���H� ����=��4=�Z=���<��R=��=G�������q`���u<�"<�j=q�F>�t�>"s]?�o�>ƒ�>ܻ7?� ���6�IT���P0?V�:=8��8煾˂����l�>��k?���?P;Z?/�_>��A�łC��>�`�>l�'>��\>G��>�I��scI����=8�>e�>�d�=j"Z�0=���
�s葾���<rd>[��>M'|>h ����'>�z��~$z���d>1�Q��ú�^�S�c�G���1�ߎv��K�>��K?��?#��=�]龰%���Df�t/)?�]<?QM?��?��=I�۾�9���J��K���>AƩ<��{���"���:�R��:�s>�-���۟���c>;����޾g�n�C�I�d���\=E��� O=�d���־��z��#�=�h>�i���� �2:��㲪��I?��i=�ꤾ��T��9���>ď�>H+�>uD�Ur�Ր@�񄬾Yb�=�Y�>F�;>�)���\^G����S�>�!A?��`?��?�ޅ�c�\�2�r�	���|��5[�{�?2H�>**?J�A>�і=t]�����N9d��N<����>���>�����G�:���K���!$��΂>s��>�SE>�A?ݐC?�G?yXb?_�2?¬�>�ʐ>�d����оwB&?��?�=��Խ��T���8�F��>��)?-�B�o��>��?#�?F�&?U�Q?z�?;�>�� ��A@����>�Y�>��W��a��E�_>��J?���>F=Y?�҃?��=>ʆ5�\袾�ة�"Z�=�>��2?z5#?Ӯ?���>�}�>@������=��>c? @�?��o?�O�=R#?��2>���>��=���>ͮ�>u ?�`O?)�s?a�J?�Z�>�i�<Eά�������r���S��Ì;��K<<�y=����t�m-�q �<���;������������pfD��쒼I�;���>�s>Ձ���D5>��ľ������B>O
˼��� C��d�<�~��=�!~>~�?uɓ>�j"���=���>��>�����'?Z�?��?�Ȑ;�ya�>پg�N��}�>8�??{y�=�&m�Iؓ��v��ve=�6n?�w]?A�Y������Y?;�W?���6�.�~�������u��g�f?��?�����>uz-?�7�?֚=? %|���w��@����{�wdW��.'>�ظ>�<�X�e��E�>7�C?���>��?�w[�$������־�Q3?� �?�۳?��p?�]>
�n���ѿyM�����C�]?��>� ����"?��߻_о07��R�����a������씾J`��$�bd���(׽���=6�?�!s?�q?�~_?v �W�c��]�����U�|W�|�&�E���D�-jC�s�n��b��(��v���H�H=8l��Y���?}�?䇆��|6?��6���0~;DbV>I�$�<k.�;�[%�0D�=�y=�,����ٵ�� �?���>�K�>�/?�Zm�&-�!]���3�+����s>���>��>$�?�T��˖v�<���D���������l�q>�a?��N?#o?�R+�Fb1���n�R/$��a�Q7��_>��=B��>jL�ݤ�
�$�+�G�f�n����f������={[,?���>�5�>��?���>3n��}��;����;���C���>}Q?<(�>6�>�ㆽ�W�of�>i?�`�>l��>㈾�#�Js��^�����>���>�>p��>��3���X�����Ɗ�d8��t�=�7i?zd����Y��>�+R?:y���)<r�>H��֊������.�R��=�0?8��=x�;>�F��'_	�.C�~5��i�*?��?Z��ā-�
�>/,#?,��>�s�>6/�?9W�>�žĻ�<�?h�Z?ǽI?�`>?:��>yC=�]����Ľ�@$���:=
��>�wV>�gN=_��=����LQ����̷=�D�=�4-����+EN<����2�<��=��+>kvԿ�WF���ȾԾ��g�۾8$�]@�� �ļ|�����q�о��ʾ��J�#��ֹ���lw�����IP���)\�2��?�@�*c���־8��s��~�m��>8�?�XP���U�Vܷ��5��5;`��T���[��8Y�&M�̔'?^���ֽǿ"����9ܾ� ?�@ ?+�y?����"���8�E� >B�<�-��f��ٚ����ο�����^?���> ��7�����>B��>&�X>8Iq>����鞾�2�<��?I�-?|��>	�r���ɿ���4�<���?=�@��A?%k(�J	쾃�X=���>�	?&	@>(2����/Q��,��>�Y�?֠�?�K=D�W�(���d?CU<��E������=��=�?=���4�J>s�>����G@���ܽ&�2>�r�>E���*��S]�@)�<�]>3ؽTS��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=u6�񉤻{���&V�}��=[��>c�>,������O��I��U��=�����Rɿ��$�&��6�=��o<F&���`��N߼grl�-�ξ�Ɯ������S=y,g>�7�>{�g>{<>Q�@>h�O?��|?*�>g��=��1�A����D׾�)2=V�*�	z(�{�j�7A��ի���ؾ���Jx2�:�'��b�����)=�}+�=$R�8���� ���b�A�F���.?��$>u�ʾ�M�uE%<�KʾU����f��E�[̾��1�!	n��П?�:B?��Z-W�
��{��h����W?kl�,��M����Y�=�j��XT=Є�>ќ�=�����2��YS�ه]?!�?�7�����}�>�T��sM�[u�>��-?�?�>�>�?�ֹ���?���>����r>\�?��?����xCZ��_?�[y?���)4��.e?b���v���a��s�>#{�����|�>vN����������\�zdR�Va?�a�>j�.�{z9��ި�C�.=��۽��v?I��>�4�>iRm?��Q?a�=e�:E�i��o� ;2�R?���?�	4>�<�aȾ����WX^?|݀?�b>d{�f�վ�F��,�_�I?p2V?�I�>v�=QR�%~��KԾP�H?�Z_?��%��Ц�����<z>e�,>&�?��?��Ԟ�\(?��������w����$��_�?'@ ��?�8P�f_��r���?|'�>��������A�Ǥ���	>��>?���xU�������T��?�w?ϩ?_�c��r��X�=�6��ج?O�|?�Y۾ū�=$�ϓh�v��[-�=�o3>Kr=<��F��!1�o�˾խ��"��]wU��D�>��@��I�S)�>r.���"�d¿iy��l��b%�!<?k��>���<߄��n>v���z�>�Y���Q���F���>8�>�b��X現��~���>�G@�d��>|�j��`�>��E�(ݵ����ֹ<r��>|��>��>R�ɽ{~���0�?���+Ͽ�&������^U?�̟?9%�?ϯ?a������S����t�<�hO?lr?5�V?]�
���r�~%?���j?���z�_���3�oE���S>�/3?$��>p-��@�=`'>� �>��>.��xĿv涿�_����?=L�?n�꾨n�>H��?Z�+?�������Q3��r%+��-���@?�3>N4��3!��<��䒾TV
?}/?���OA�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?~��>P��?d�=rX�> ��=Ff���/[>$�>2�P�
� ?��N?�)�>Ϊ�=F?�$P-���E��>Q�_��qC��O�>��`?�K?�}[>����e.�|� �m�Ľ,�2������H���#�ֽl�:>y}:>�>�G�Jzվs+?G��Ifٿ�]��p<;���>|��=�(?�p ��X��=�D?S�.>���A��Ԓ��=����?z-�?�?�ľU`!�>VE>��>�_�>����<��,�����>>Y�$?c{ �LY��d@{��X�>���?��
@2��?�I��'?�L���|��_���1{�z����\���7?;��Mi��z�>�^���������Z��#�>E̷?��?���>��V?�yZ�*�!�V[o>�8�>�Q?���>矖<�V较��<'��>�s �����u��M^?�	@�@�!�?I���TRٿ#V����Ǿ:����=2�=�>FI��پt>Z�=}�]<y�<�rM=��y>�}�>3Vk>�(>���=B��<��bc ����� ʐ�v%@�hd��t�#�f���꾇�^��:�Zݤ�|̾\GJ�}�½`=)�Wi�\D@�%��<J�>�MH?t��?|K�?��>�wO=X�>�ZF��O�=ڿ�;��=���>��#?��7?�S?���>�%���oE���r��T��6�D��6�>���=�*�>��e>���=q��=�&�</�>U��>�8��z�=�{<x0�=�m�>d�>�
�>U�$>��<>�4>O������,�h���v��Bɽ��?Ͼ���J�0��]���'������=�n.?�}>����3Cп�歿�H?*唾j���+���>��0?�3W?H*>����R�6>	����j��A>H���o�l�o])�قP>�A?���>q7�>����Y(��-`�Pd¾�{?၇?��)��R���틿8F\��^@=4�?���>�����>�����vi�#9�Hn�:?���>��[����)�56����=��>���<�7>4�<�P����,�~�	�O,;�u=��c>�?�j>� >4<�>`����J�Y.�>��=Y�e>�&5?�c?fY>�J��I�����K�:>F��>;�m>�F>��}��z�=�{�>�R�>�X;���2�<��� 0�� �{>�S%�of��Vy�դ�=9*��j�>�e>M����q�[�?;�~?w��䈿��f���lD?�+?��=^�F<��"�J ���H��L�?r�@m�?��	�ƢV���?�@�?�
��ܷ�= }�>	׫>�ξ,�L�ӱ?D�Ž�Ǣ���	��)#�GS�?��?�/�?ʋ�*l��6>�^%?˰Ӿ�N�>^9��/������ô]�I���6X�>b�I?ކ�{	�T����>�c�>5N澛/��=�ʿd-q��\�>7�?�"�?/�^�R����jC�
	?���?��S?�n|>3w�2�G��`�>��A?1Z8?g˓>�%�L$*�Ev$?��?tC�?��L>�)�?G�s?��>�񂽰+��s��81�����=���Ý�>su>�{��=�C������O��ޒi�6���md>��=�Ⱥ>��ݽ-��pæ=E���D��ڃh����>�#w>�L>X�>��?���>���>
��<R���Os��� ���nL?���?���B7j�����9�=�D���%?�?���lM��k>:u?�M�?��]?+�B>�c
��۠�K7��]���+�;H[>~�>1��>_"���5>B���ș�M��>y�?>�1�t��qCy���=86}>^6?V��>�=<�?�?+�{>���>.�_��j�����-��>c%?�G,?��? ��>�w�W������WP�L�*j7>7)b?ټA?�ɳ>��j�	e>�9������?iyZ?��Z��p ?��`?-wu?� G?�s>2�X����ȢF�b��>��"?\����@���%��� �&.?�[?v0�>ߠǽ���
X��H���߾�w?ã\?i�?A��gf��7ƾ�X�<��[����;0�<�H�>�>h0t���=Ʌ&>��=�h��Y?�Y&<r��=F!�>�~�==�;�溊��p)?$:pV����=#s��:8�r�4>��<> ���[?���f�z�_g���R��3΄��{�?���?�a�?�[��5Be�F9?c��?��?���>��������h�u�t���R�8����C>c�>}�Y<�t�ǫ���_���Ȃ�S5�� �
U�>(��>!?�X�>��5>�V�>K�Ӿ����+��u���1]�}�eh �(0�l@�����B3��'�<����.����Ks>ḽ��k�>�]�>J�>�R!>�p>ꢥ=[��>�]�=��}=���>R��=T�>��Z>Y�g=N=b:]R?.���@'��g꾿�����=?�<h?��>[���愿��	���?۴�?ෞ?�ށ>�Xi�/M)�Y��>�9�>y8z�yY?�{R=�y�Q3^<���E��y�t���d�6v�>��XW6��L�Kf�+?�?	����̾F?ؽ�]���6�=Oh�?�1??�&� TP���P��\��@H�Ҍ̺n����)о��#�Y@X���:���0˃�W
��*�=ǋ0?�\{?/������䓾�cu�C�T�䝏>��>�p�>�?ZQ>����"���Y�(�!����ri?�&g?܈>FG?$�G?�g[?|�H?#�>W��>��Ǿ3��>F��<K�>)��>7�8?y-?Ч8?w!?σ?�@>@,�"$����վ"@?J]?��?���>�[�>�Zv�L�Ž+���F�����j�t�G	�=� �<����ke�G=
0d>�d%?�����7����2�>A?��>i��>�Qe��L�t!<ܦ?��?cMN>m��,h����ŝ�>��?9���uj=�V;>^�=G��<�iN<c@�=���>uZ�=��a=��T�0��=P-\=	��<��0=�W=��<��>y;	?�)r=0�>�}P���Ҿ/69�V>=����v=�>u�=���h����]�'�>d��?���?�q�=ɪ=�=V���C�p�s�9�[�S�K�=�H�>�Z�>z��?qM�?;�!?��(?R?>��i�������=���?P`/?�ߥ>�,�1�Ǿ�8��L� ��r$?X�?!dy��^�O=5���þ��=om�>�^׾�{r��꧿��b��>�׏�󵇽I��?��?kP��?%�I�����b�ؽ�$/?ݠ�>]��>�x�>a^O�k�I�'��&��I?�H?1C�>o N?���?�[f?��k>�0��¨������D<G2=>��B?'v?�~�?�r?��><_>��'��_ݾv����K���׽}�k���=� c>3o�>���>��>���=^���f'���F�Bz�=fr>���>J��>���>T+�>ٞQ���G?���>F��ş�٦��� ��c3G��~u?�8�?/e*?c�=���mF��&��m��>�h�?wL�?c�*?��U���=ʿݼ�޵��sq�	�>[��>�>!��=�H=�>Uf�>>�>���XE�C98�t!L���?)nE?��=;ƿb�s�Ƴt�p���í�<�s���d��Β���W�m��=i���$���k��`�Y�C����̺�������	}����>-�=���=t��=\2�<Z#��$b<��H=+�<h�=��u��WT<e�(� )������F7<�|Z<4�C=.N���ʾg;z?�C?�$?��C?�M}>�>��[����>�>C?�^>������ʾ�P�`y���n��a�Ǿr�8�p��w��&�>��K�*M>�>"��=�<���=�=��m=�W5�h"=(��=���=���=���=�>�>�6w?K�������4Q��Y罋�:?�8�>�{�=��ƾ?@?p�>>�2�������b��-?���?�T�?[�?�ti��d�>T���⎽�q�=���>2>P��=��2�:��>%�J>����J������s4�?��@��??�ዿ͢Ͽga/>Gj>�O>�zI�/M-�����?� �B�}?x�D�Pv޾d��>0��=����]ﾈ��vi>k��=0c��~e����<�սOW�=z�>=nB�>�%>jէ=�y��K%�=Y��=�0�=so0>,�;�{��;��eP�=��=�~J>��D>�H�>f�?n�0?0�d?$!�>Z�m�N�ξY9¾�9�>���=�)�>]��=q�B>�z�>�38?�E?�RK?�}�>.<�=�]�>ئ>�,��8m����A��^�<���?���?�q�>c�<�7C��V�q>�BjýjO?�71?)�?ҝ>%r����uc5���־{�>~�>�7���:L�s:м�H�����+��>X>�d>6"�>���>a��=P,X�3C�=,{�>¸�=_��$#>�^B=�V	=����k�=3X�,3'�����B�w�=�����s�=�N>j�@=rv�<��I<���=�*�>���=���>�t�,�m�nN�=�P���f����=�"��+���b�����h�F�E0��]��>��>��z��N��FL�>�P>�U�=���?FX?h�>x�#��"��������^��M�<�>=ܫ=b��+�M�q��/�E�1z�>�ew>���>�	�>t�$���9�=j���R
�J�>��:���6>�Y�>C�n��Iە���_�TK=F6C?aą��[�=�?	\?��?���>Zc���
���>n�վYG\���$�M�Q�̲B��?qL?t�>+��#-�v����������>4��dM�{���Z(���(��������>�Ƥ����;�2�H�������,tC����P/�>UQ?ه�?�wf�m6��3R��&	�)꽟k�>�rp?B�>��?�?Kd���FF��B�=kd?��?���?�7>��=$���Kk�>/�?��?\��?��s?��b�_��>FĻ���=��8����=^->q�K=��=�K?M'?��?񿬽�M����-`��^�h&�<��=���>].�>�7W>	5�=�N�<I��=��U>(��>dr�>JNe>��>�w>c��)0��Q2?[��=�\>�)&?��>�B�>?n���H=鎳=�v����q�  ��o�g>�&�=J>�7��>$�Կţ�?YU>5�K�:?������<�ѐ>�Ԗ>��\�`��>��>���>ĕ�>mA�=��=�~>��l>�l�J�_>D\�lH5�b`,�Z�o�@����>��N��җ�������9�Vf#�R磾�$(�3�y��]����+�\��<�L�?*�=ܟ����Y��A<Z��>�h�>�3?举�UN�b�>�
?�E>ց龖��$v��(���]��?��?E:c>%�>��W?R�??�1��3��pZ�íu��'A��e���`��፿�����
����>�_?p�x?�wA?㐒<�<z>9��?��%�+Ώ�+)�>t/�);�oM<=�(�>�����`���Ӿ��þ�6��=F>d�o?�%�?�Z?\WV������V>�,T?xHM?N>Y?��>?^�-?0O��'?�d>���>�x�>��)?)�4?&�(?���>XJ�=�,������9��̢e�����)L�E���%n�=C9�=���!���=w=�y�<���<�H�=%�<�=�!=�G=�GB=Rͫ>ɰZ?���>ht>�Y:?0���a<�3E���},?�=�z������j�� ������=�Bi?C��?��^?ifZ>.0<�u G���'>b��>�&
>�MU>�C�>F����?����=;>�f>$�=W�I�\=��h���獾�j�9�>�n�>�V�>ޱ)=c	g>�n�N`���̀>��z�0U���F�nJ�Y�㻭����>�U?�E�>*��=K��Bk��m�#?8A?,WX?Hp?̔ɻ����nm_�Wi޾��P�cCg>ܣ��j�#�]�������kB(����A2�>��/��۟���c>;����޾g�n�C�I�d���\=E��� O=�d���־��z��#�=�h>�i���� �2:��㲪��I?��i=�ꤾ��T��9���>ď�>H+�>uD�Ur�Ր@�񄬾Yb�=�Y�>F�;>�)���\^G����S�>�!A?��`?��?�ޅ�c�\�2�r�	���|��5[�{�?2H�>**?J�A>�і=t]�����N9d��N<����>���>�����G�:���K���!$��΂>s��>�SE>�A?ݐC?�G?yXb?_�2?¬�>�ʐ>�d����оwB&?��?�=��Խ��T���8�F��>��)?-�B�o��>��?#�?F�&?U�Q?z�?;�>�� ��A@����>�Y�>��W��a��E�_>��J?���>F=Y?�҃?��=>ʆ5�\袾�ة�"Z�=�>��2?z5#?Ӯ?���>�}�>@������=��>c? @�?��o?�O�=R#?��2>���>��=���>ͮ�>u ?�`O?)�s?a�J?�Z�>�i�<Eά�������r���S��Ì;��K<<�y=����t�m-�q �<���;������������pfD��쒼I�;���>�s>Ձ���D5>��ľ������B>O
˼��� C��d�<�~��=�!~>~�?uɓ>�j"���=���>��>�����'?Z�?��?�Ȑ;�ya�>پg�N��}�>8�??{y�=�&m�Iؓ��v��ve=�6n?�w]?A�Y������Y?;�W?���6�.�~�������u��g�f?��?�����>uz-?�7�?֚=? %|���w��@����{�wdW��.'>�ظ>�<�X�e��E�>7�C?���>��?�w[�$������־�Q3?� �?�۳?��p?�]>
�n���ѿyM�����C�]?��>� ����"?��߻_о07��R�����a������씾J`��$�bd���(׽���=6�?�!s?�q?�~_?v �W�c��]�����U�|W�|�&�E���D�-jC�s�n��b��(��v���H�H=8l��Y���?}�?䇆��|6?��6���0~;DbV>I�$�<k.�;�[%�0D�=�y=�,����ٵ�� �?���>�K�>�/?�Zm�&-�!]���3�+����s>���>��>$�?�T��˖v�<���D���������l�q>�a?��N?#o?�R+�Fb1���n�R/$��a�Q7��_>��=B��>jL�ݤ�
�$�+�G�f�n����f������={[,?���>�5�>��?���>3n��}��;����;���C���>}Q?<(�>6�>�ㆽ�W�of�>i?�`�>l��>㈾�#�Js��^�����>���>�>p��>��3���X�����Ɗ�d8��t�=�7i?zd����Y��>�+R?:y���)<r�>H��֊������.�R��=�0?8��=x�;>�F��'_	�.C�~5��i�*?��?Z��ā-�
�>/,#?,��>�s�>6/�?9W�>�žĻ�<�?h�Z?ǽI?�`>?:��>yC=�]����Ľ�@$���:=
��>�wV>�gN=_��=����LQ����̷=�D�=�4-����+EN<����2�<��=��+>kvԿ�WF���ȾԾ��g�۾8$�]@�� �ļ|�����q�о��ʾ��J�#��ֹ���lw�����IP���)\�2��?�@�*c���־8��s��~�m��>8�?�XP���U�Vܷ��5��5;`��T���[��8Y�&M�̔'?^���ֽǿ"����9ܾ� ?�@ ?+�y?����"���8�E� >B�<�-��f��ٚ����ο�����^?���> ��7�����>B��>&�X>8Iq>����鞾�2�<��?I�-?|��>	�r���ɿ���4�<���?=�@��A?%k(�J	쾃�X=���>�	?&	@>(2����/Q��,��>�Y�?֠�?�K=D�W�(���d?CU<��E������=��=�?=���4�J>s�>����G@���ܽ&�2>�r�>E���*��S]�@)�<�]>3ؽTS��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=u6�񉤻{���&V�}��=[��>c�>,������O��I��U��=�����Rɿ��$�&��6�=��o<F&���`��N߼grl�-�ξ�Ɯ������S=y,g>�7�>{�g>{<>Q�@>h�O?��|?*�>g��=��1�A����D׾�)2=V�*�	z(�{�j�7A��ի���ؾ���Jx2�:�'��b�����)=�}+�=$R�8���� ���b�A�F���.?��$>u�ʾ�M�uE%<�KʾU����f��E�[̾��1�!	n��П?�:B?��Z-W�
��{��h����W?kl�,��M����Y�=�j��XT=Є�>ќ�=�����2��YS�ه]?!�?�7�����}�>�T��sM�[u�>��-?�?�>�>�?�ֹ���?���>����r>\�?��?����xCZ��_?�[y?���)4��.e?b���v���a��s�>#{�����|�>vN����������\�zdR�Va?�a�>j�.�{z9��ި�C�.=��۽��v?I��>�4�>iRm?��Q?a�=e�:E�i��o� ;2�R?���?�	4>�<�aȾ����WX^?|݀?�b>d{�f�վ�F��,�_�I?p2V?�I�>v�=QR�%~��KԾP�H?�Z_?��%��Ц�����<z>e�,>&�?��?��Ԟ�\(?��������w����$��_�?'@ ��?�8P�f_��r���?|'�>��������A�Ǥ���	>��>?���xU�������T��?�w?ϩ?_�c��r��X�=�6��ج?O�|?�Y۾ū�=$�ϓh�v��[-�=�o3>Kr=<��F��!1�o�˾խ��"��]wU��D�>��@��I�S)�>r.���"�d¿iy��l��b%�!<?k��>���<߄��n>v���z�>�Y���Q���F���>8�>�b��X現��~���>�G@�d��>|�j��`�>��E�(ݵ����ֹ<r��>|��>��>R�ɽ{~���0�?���+Ͽ�&������^U?�̟?9%�?ϯ?a������S����t�<�hO?lr?5�V?]�
���r�~%?���j?���z�_���3�oE���S>�/3?$��>p-��@�=`'>� �>��>.��xĿv涿�_����?=L�?n�꾨n�>H��?Z�+?�������Q3��r%+��-���@?�3>N4��3!��<��䒾TV
?}/?���OA�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?~��>P��?d�=rX�> ��=Ff���/[>$�>2�P�
� ?��N?�)�>Ϊ�=F?�$P-���E��>Q�_��qC��O�>��`?�K?�}[>����e.�|� �m�Ľ,�2������H���#�ֽl�:>y}:>�>�G�Jzվs+?G��Ifٿ�]��p<;���>|��=�(?�p ��X��=�D?S�.>���A��Ԓ��=����?z-�?�?�ľU`!�>VE>��>�_�>����<��,�����>>Y�$?c{ �LY��d@{��X�>���?��
@2��?�I��'?�L���|��_���1{�z����\���7?;��Mi��z�>�^���������Z��#�>E̷?��?���>��V?�yZ�*�!�V[o>�8�>�Q?���>矖<�V较��<'��>�s �����u��M^?�	@�@�!�?I���TRٿ#V����Ǿ:����=2�=�>FI��پt>Z�=}�]<y�<�rM=��y>�}�>3Vk>�(>���=B��<��bc ����� ʐ�v%@�hd��t�#�f���꾇�^��:�Zݤ�|̾\GJ�}�½`=)�Wi�\D@�%��<J�>�MH?t��?|K�?��>�wO=X�>�ZF��O�=ڿ�;��=���>��#?��7?�S?���>�%���oE���r��T��6�D��6�>���=�*�>��e>���=q��=�&�</�>U��>�8��z�=�{<x0�=�m�>d�>�
�>U�$>��<>�4>O������,�h���v��Bɽ��?Ͼ���J�0��]���'������=�n.?�}>����3Cп�歿�H?*唾j���+���>��0?�3W?H*>����R�6>	����j��A>H���o�l�o])�قP>�A?���>q7�>����Y(��-`�Pd¾�{?၇?��)��R���틿8F\��^@=4�?���>�����>�����vi�#9�Hn�:?���>��[����)�56����=��>���<�7>4�<�P����,�~�	�O,;�u=��c>�?�j>� >4<�>`����J�Y.�>��=Y�e>�&5?�c?fY>�J��I�����K�:>F��>;�m>�F>��}��z�=�{�>�R�>�X;���2�<��� 0�� �{>�S%�of��Vy�դ�=9*��j�>�e>M����q�[�?;�~?w��䈿��f���lD?�+?��=^�F<��"�J ���H��L�?r�@m�?��	�ƢV���?�@�?�
��ܷ�= }�>	׫>�ξ,�L�ӱ?D�Ž�Ǣ���	��)#�GS�?��?�/�?ʋ�*l��6>�^%?˰Ӿ�N�>^9��/������ô]�I���6X�>b�I?ކ�{	�T����>�c�>5N澛/��=�ʿd-q��\�>7�?�"�?/�^�R����jC�
	?���?��S?�n|>3w�2�G��`�>��A?1Z8?g˓>�%�L$*�Ev$?��?tC�?��L>�)�?G�s?��>�񂽰+��s��81�����=���Ý�>su>�{��=�C������O��ޒi�6���md>��=�Ⱥ>��ݽ-��pæ=E���D��ڃh����>�#w>�L>X�>��?���>���>
��<R���Os��� ���nL?���?���B7j�����9�=�D���%?�?���lM��k>:u?�M�?��]?+�B>�c
��۠�K7��]���+�;H[>~�>1��>_"���5>B���ș�M��>y�?>�1�t��qCy���=86}>^6?V��>�=<�?�?+�{>���>.�_��j�����-��>c%?�G,?��? ��>�w�W������WP�L�*j7>7)b?ټA?�ɳ>��j�	e>�9������?iyZ?��Z��p ?��`?-wu?� G?�s>2�X����ȢF�b��>��"?\����@���%��� �&.?�[?v0�>ߠǽ���
X��H���߾�w?ã\?i�?A��gf��7ƾ�X�<��[����;0�<�H�>�>h0t���=Ʌ&>��=�h��Y?�Y&<r��=F!�>�~�==�;�溊��p)?$:pV����=#s��:8�r�4>��<> ���[?���f�z�_g���R��3΄��{�?���?�a�?�[��5Be�F9?c��?��?���>��������h�u�t���R�8����C>c�>}�Y<�t�ǫ���_���Ȃ�S5�� �
U�>(��>!?�X�>��5>�V�>K�Ӿ����+��u���1]�}�eh �(0�l@�����B3��'�<����.����Ks>ḽ��k�>�]�>J�>�R!>�p>ꢥ=[��>�]�=��}=���>R��=T�>��Z>Y�g=N=b:]R?.���@'��g꾿�����=?�<h?��>[���愿��	���?۴�?ෞ?�ށ>�Xi�/M)�Y��>�9�>y8z�yY?�{R=�y�Q3^<���E��y�t���d�6v�>��XW6��L�Kf�+?�?	����̾F?ؽ�]���6�=Oh�?�1??�&� TP���P��\��@H�Ҍ̺n����)о��#�Y@X���:���0˃�W
��*�=ǋ0?�\{?/������䓾�cu�C�T�䝏>��>�p�>�?ZQ>����"���Y�(�!����ri?�&g?܈>FG?$�G?�g[?|�H?#�>W��>��Ǿ3��>F��<K�>)��>7�8?y-?Ч8?w!?σ?�@>@,�"$����վ"@?J]?��?���>�[�>�Zv�L�Ž+���F�����j�t�G	�=� �<����ke�G=
0d>�d%?�����7����2�>A?��>i��>�Qe��L�t!<ܦ?��?cMN>m��,h����ŝ�>��?9���uj=�V;>^�=G��<�iN<c@�=���>uZ�=��a=��T�0��=P-\=	��<��0=�W=��<��>y;	?�)r=0�>�}P���Ҿ/69�V>=����v=�>u�=���h����]�'�>d��?���?�q�=ɪ=�=V���C�p�s�9�[�S�K�=�H�>�Z�>z��?qM�?;�!?��(?R?>��i�������=���?P`/?�ߥ>�,�1�Ǿ�8��L� ��r$?X�?!dy��^�O=5���þ��=om�>�^׾�{r��꧿��b��>�׏�󵇽I��?��?kP��?%�I�����b�ؽ�$/?ݠ�>]��>�x�>a^O�k�I�'��&��I?�H?1C�>o N?���?�[f?��k>�0��¨������D<G2=>��B?'v?�~�?�r?��><_>��'��_ݾv����K���׽}�k���=� c>3o�>���>��>���=^���f'���F�Bz�=fr>���>J��>���>T+�>ٞQ���G?���>F��ş�٦��� ��c3G��~u?�8�?/e*?c�=���mF��&��m��>�h�?wL�?c�*?��U���=ʿݼ�޵��sq�	�>[��>�>!��=�H=�>Uf�>>�>���XE�C98�t!L���?)nE?��=;ƿb�s�Ƴt�p���í�<�s���d��Β���W�m��=i���$���k��`�Y�C����̺�������	}����>-�=���=t��=\2�<Z#��$b<��H=+�<h�=��u��WT<e�(� )������F7<�|Z<4�C=.N���ʾg;z?�C?�$?��C?�M}>�>��[����>�>C?�^>������ʾ�P�`y���n��a�Ǿr�8�p��w��&�>��K�*M>�>"��=�<���=�=��m=�W5�h"=(��=���=���=���=�>�>�6w?K�������4Q��Y罋�:?�8�>�{�=��ƾ?@?p�>>�2�������b��-?���?�T�?[�?�ti��d�>T���⎽�q�=���>2>P��=��2�:��>%�J>����J������s4�?��@��??�ዿ͢Ͽga/>Gj>�O>�zI�/M-�����?� �B�}?x�D�Pv޾d��>0��=����]ﾈ��vi>k��=0c��~e����<�սOW�=z�>=nB�>�%>jէ=�y��K%�=Y��=�0�=so0>,�;�{��;��eP�=��=�~J>��D>�H�>f�?n�0?0�d?$!�>Z�m�N�ξY9¾�9�>���=�)�>]��=q�B>�z�>�38?�E?�RK?�}�>.<�=�]�>ئ>�,��8m����A��^�<���?���?�q�>c�<�7C��V�q>�BjýjO?�71?)�?ҝ>%r����uc5���־{�>~�>�7���:L�s:м�H�����+��>X>�d>6"�>���>a��=P,X�3C�=,{�>¸�=_��$#>�^B=�V	=����k�=3X�,3'�����B�w�=�����s�=�N>j�@=rv�<��I<���=�*�>���=���>�t�,�m�nN�=�P���f����=�"��+���b�����h�F�E0��]��>��>��z��N��FL�>�P>�U�=���?FX?h�>x�#��"��������^��M�<�>=ܫ=b��+�M�q��/�E�1z�>�ew>���>�	�>t�$���9�=j���R
�J�>��:���6>�Y�>C�n��Iە���_�TK=F6C?aą��[�=�?	\?��?���>Zc���
���>n�վYG\���$�M�Q�̲B��?qL?t�>+��#-�v����������>4��dM�{���Z(���(��������>�Ƥ����;�2�H�������,tC����P/�>UQ?ه�?�wf�m6��3R��&	�)꽟k�>�rp?B�>��?�?Kd���FF��B�=kd?��?���?�7>��=$���Kk�>/�?��?\��?��s?��b�_��>FĻ���=��8����=^->q�K=��=�K?M'?��?񿬽�M����-`��^�h&�<��=���>].�>�7W>	5�=�N�<I��=��U>(��>dr�>JNe>��>�w>c��)0��Q2?[��=�\>�)&?��>�B�>?n���H=鎳=�v����q�  ��o�g>�&�=J>�7��>$�Կţ�?YU>5�K�:?������<�ѐ>�Ԗ>��\�`��>��>���>ĕ�>mA�=��=�~>��l>�l�J�_>D\�lH5�b`,�Z�o�@����>��N��җ�������9�Vf#�R磾�$(�3�y��]����+�\��<�L�?*�=ܟ����Y��A<Z��>�h�>�3?举�UN�b�>�
?�E>ց龖��$v��(���]��?��?E:c>%�>��W?R�??�1��3��pZ�íu��'A��e���`��፿�����
����>�_?p�x?�wA?㐒<�<z>9��?��%�+Ώ�+)�>t/�);�oM<=�(�>�����`���Ӿ��þ�6��=F>d�o?�%�?�Z?\WV������V>�,T?xHM?N>Y?��>?^�-?0O��'?�d>���>�x�>��)?)�4?&�(?���>XJ�=�,������9��̢e�����)L�E���%n�=C9�=���!���=w=�y�<���<�H�=%�<�=�!=�G=�GB=Rͫ>ɰZ?���>ht>�Y:?0���a<�3E���},?�=�z������j�� ������=�Bi?C��?��^?ifZ>.0<�u G���'>b��>�&
>�MU>�C�>F����?����=;>�f>$�=W�I�\=��h���獾�j�9�>�n�>�V�>ޱ)=c	g>�n�N`���̀>��z�0U���F�nJ�Y�㻭����>�U?�E�>*��=K��Bk��m�#?8A?,WX?Hp?̔ɻ����nm_�Wi޾��P�cCg>ܣ��j�#�]�������kB(����A2�>��/�����Eb>�v� �ݾ~[n��I�SG��wI=A����S=���R
־ !��=��
>�i���� �����Ъ�a�I?�f=]����U� ع���>�>_
�>�=���y�L@�[p��S�=��>%!<>}��Z�cG��N�
�>��9?��`?iՉ?��,�U���+�	�8,������SL?��>j}�>���>KS4=�괾U���]��:�E=�>��>1��W�C�@h�Ԩؾ�*���>'�>p
>>M?y�:?�V?EaW?
�:?7?m��>O1����ʾ%D&?���?W��=V�Խ��T�K9��F�V��>W�)?��B����>��?��?!�&?ҀQ?$�?z�>2� �>;@���>]�>��W��e��O`>��J?>��>�3Y?3؃?n>>�5�Jߢ�ͩ�K5�=�>T�2?S1#?�?��>�[�>�w��1�=u6�>R�k?Wg~?*Bp?Bg>�>�U*>u��>�}g=�f�>X��>6h?�UP?��h?ͧ@?��>2�<�D׼ZA���
C��j$;U�a=�A�;�-=<"��5���H}�t7<���\��i�f�6V�p!׼�&���o!�> �D>�<�ˤ�>$��T���k�>LV޽��h���%�;(�(�%>�&�>!�
?�<>��R�X�L�� �>���>���Ba(?��
?+!8?oo�=�`��K'�"IپBr�>~:?�K-�po�r{�����������f?:�O?Tj�\�澗`Y?�tQ?o 	�mK��_����ѽ�/ܾsJR?�3?=w��3%W>���?5�?�C�>�И�����>��I�U��Ǔ�=7Um>���}�c��Vs>u-=?"?��?>*=��ǾGS���w���p?���?z�?�΀?��1>�WY���ݿ�?���ț���d?$Կ>��ɾ~y0?�rn�m?Ҿ��V����?龮�����.b������ ,��Д���ؽ��<�0?�#�?�Fb?6�]?����~\p���\�۬��9'H�7�Ҿ����5N���E��<5�V�o�{y
�j��0O��jl�=Ć�N'd�)�?��?(ń��#?�Z��Q����=F;>w���%\�n7=�� ����=��b=�ǅ��y-�Z�ξ��$?��>�6�>*�5?KPX�RA�%�-��V=�0pؾ!�|>���>�?Q>���>'��<��Y����Q�̾�V��^����>�_?9-O?f��?X�:�K<�
�[��b>��s�jσ�)�A>�n>��{>n4�y^O�� �Q\5���q�@�����L��lXY=N�(?�|�>�w�><R�?%?XO!�澭�φ>�q<����=/��>�5e?���>���>Ϫ'�Wz ��!?I�?�d>hs�><��A1 �+C�W�����?N��>,�>X?�>n�P�#��Շ�`׌���2��,�>�ғ?�)}�ؒ��(h>��m?�i4��½m7�>��P>��F�/J��#�=x��>���>���=Xg>�o¾`"��T�����9*0?0?���9�,��8�>=*?f��>p�h>��?�=�>��Ͼ�EZ<??��[?yV8?��1?���>r�=�n.�w´;���l�<
]�>��F>ɇ�<�  >���m�?��%�q�=�a�=%���o^��%��<S�ü�-Y<�<D�1>��֒V��Tξ�
���:�	{���r�=?�x��F���������H�`�6��b��V��p��j�,�t����?Cf�?�������#����
]� 4¾���>/CF���#� �۾<���.n:��Z~�f����1��V��=e� 	K���'?,���k�ǿ����+;ܾ[ ?�7 ?U�y?"���"���8�Ŭ >\�<᜜���#�����ο���,�^?���>���g��|��>F��>ՠX>s1q>P������<��?/�-?t��>[�r���ɿ�������<���?�@q�A?az(���ӯV=e��>B�	? �?>��1��������V�>b4�?�݊?�yO=_�W��S�#e?�<&yF���໭?�=�=�`=�����J>��>�Y���A���ܽp�4>J܅>N�"�v���1^��m�<�]>��ս�|�o?�xN�{Ct��MD���g����<9E?��>��U�x�?�B�}�տC�g�4R?��@ĵ�?�G?p���ڭ>.�Ѿ�\G?Ym6?�[�>Z�2��p��j>P<0�o%�=�����M�똔=��>-��=Іg������S8�=��ͻ����ƿ�#����eZ�<��N��^��U�̽R����$y������q���罛$C=���=�O>C�>[�V>=�V>�V?��j?U��>{�>/��;��N�ɾ�Aƻ����$�Ng��5�����:L��Dܾ��
��S�����	ʾ�FM���1=B�Q��-��e�"�f�b�Q*F�vB6?##>�+�(�K�e�;ES��Lݡ��`G�ӈ����Ѿ_�/� ci��{�?��C?�拿��a��
�����!b��lTS?����[���N[>�3��=^w�>�=�v羏x.���E�t�1?��?����G��C�*>a� �#/= )?j?%��;�t�>j�)?O�(�v�ӽ��P>�Y$>��>$O�>��>��������g?j�U?����:��B�>򹾔��_�F=&A>V/����ԉ_>uI�<����L�5����v�9��^?��>1p���)���ȼ\�I=K�y��a0?buJ?�a�>6w<?$�B?�ć=����=V���+�|Ly�-ux?�?<U>'F��3�QT�^:?��?���>�὾�������R:�"v0?�Tf?�[=?{b�����i��M0����?^;b?�J^��O����4��G~>e"�>�[?��<�C-�>��3?� @�+����㾿(s"�ܩ�?ln@T��?�n�[t��8==�&�>��>��:�j$���_r��䷾Κ=C��>0���~���(�^�Z�DiU?���?Ǉ?���.��s��=����;��?z�t?�LӾ�	<cQ� n���Ͼds�=e�=]�Ž��޽���8.� ��r�����������>	t@��Y�:��>���Db���ο�7}�����&���1?��W>�@;�ş���v���]��&�Zw7��K�?M�>��>ͨ��5���v�{��s;�������> F�Y�>��S��+��ɝ��;�5<��>��>���>�%���۽��Ù?�Y��=ο)������X?yc�?�l�?
q?��:<��v�w�{��,��%G?6�s?�Z?_a%�\*]�ֱ7���j?�h��� `�LR4���E��T>�3?�#�>mI-�_�}=%>���>�k>�u.�jĿ�����$��Y˦?IT�?�P�W��>���?%�+?Mq��H����\$+���{��HA?�x2>q�����!�3=��>����
?On0?v���=m^?�Ja�	�q��1/�Sl�����>�-1�|FW��%���"��d��v������s�?���?-��?���?$�]%?gv�>(G��ىž�k�<MV�>���>�Q>h�W�,/r>�����9��E>��?TF�?w?	���=���>��~?�I�>j&�?��>t�?��J�=(��C�=*J`�]�;>ݮ��p}
?ty?ի>"]a>��j�@+6��<�I!��̾�OC�{0)>0��?��U?H ��U������a<���}���:�
X�.�����߫�b%>{��>;7>9щ�������>����ڿ���B���1�?D&�=�Q?��=T��9��;�?K?��U>�����(R�����n�?B�?�_!?l�ž��w���S>�
�>�R>�a ����D���}��>��L?���Jѓ�.���<�>�3�?�B@(
�?�HO�$r�>���Ó��d~�>y��4V��=Ї���K?���y�>޴�>��`=~�v���-^�S��>�\�?3��?�h�>��e?�Z�:2�� ��Bt�>��E?�U�>
6#<8��C>���>�d�f� �##�?C@y�@�U?Z����忰���Su�����C_=�	L��tػ9��==��=�$E�uY�=�&��X�=�i>�?>B�z>[�M>pSd>�K>�����n��͗��o���(O���-���.�cPw�\����"��S���~˾�Խ�ZD�Dν���&7���}�����Zl>^�?:V?�7�?��>��>+�=��Y�+�a(
��{><�d>�)5?�`?�&?�o�=���a�}��Z��ݖ�3q�:ȳ>�v�=�^?���>�)>�2�=�ej>Y�&>T��>>5�=��->*�=]�>�{�>%��>�O�>�+�>/B<>��>7ϴ��1��:�h��
w�\̽�?ǁ��n�J��1���9�����Nh�=[b.?�|>��� ?пH����2H?���p)�&�+���>[�0?�cW?$�>����T�:>���j��`>�+ ��l���)�O%Q>}l?XC
>�s{>iE5��9�Ӝ@��O���f�>/?E߾�f�Lf{�	�_���Z�>e_�>��=���W`��d�u��o�3�=@q8?�`?�H���^��B�p��S���n>Z�P>f��<�.�=�p>���j�
���e=�b,>M�>�V?;i(>-�=���>1"���\�͒�> �>
Y+>��??��?&	�����\��|@��p>���>��n>�F�=*N�	ݳ=��>O�S>��;S@��+���.���<>� |�O�f�z���so=^Jý=��=��=���C6�B1=@�~?y��V���c�mᶽ�mD?'B?&J�=�G<"�p����(��#�?��@Ge�?X�	�p�V���?�:�?����n�=���>�٫>�8ξ`�L�5�?�Rƽ�¢�U~	�i�"�I�?�?7�/�UƋ��l�	=>?P%?o�Ӿ�o�>��ט��膿G�o��S=�p�>o�I?ϥ������A�N�?�:?#��������ɿO]y���>���?��?H�l�Q���9D��&�>^y�?�T]?*j>9g߾C�a���d>��C?�V?5��>���L<���?�g�?��?��?>h�?��u?o��>�蜽�s0�E�������s=*:ʹ^��> p�=)Y��o�D�����=҇�Ygf���HLi>ٶ1=V{�>ul½����4��=�ʟ�̯��)<��\�>l,`>�Q>���>���>��>yI�>��=�D�xn�/T��}�K?q��?���k2n�}M�<桜=��^�o&?1I4?l[� �Ͼ�ը>Ժ\?p?�[?�c�>/��O>��D迿&~��ͨ�<��K>�3�>�H�>2%��EK>��Ծ�4D�-p�>�ϗ>����G?ھ�,��;���B�>|e!?1��>�Ѯ=?��7?��j>n��>L�*�%���(Uk��ڼ>�?D�?[��?I�> e��2[a��-���Ɖ�Yj1�
��>x|?��+?+�>;��ᷯ�I|�>g�3>�>�1�z?xZ�?5;�����> ~�?k�f?ك�>��>3�پ���>h�>�A?
�1��cW���@�*���K#�>I��>Hr�>�a���)���T��y<�&����?�u�?N�N?i��Ҿt��򃾭�<c�T=���<<�<�V��?�=�fV>�Z���K�=*�>AV�=:��7���G�ȝ>��n>i��=�KZ����; =?�:�;{-��J^�x<~��_�K�z>׍u>�x���2R?����1��6m��P��)ڧ����?�\�?�S�?��=�G�c��O=?��?�s?f��>�B2�6�Ǿ+��//����P�JV���j>-�t>9�����웿ia��kf��H�X]��P�>��>��?_e�>� >♬>�R��l� �!e����=EX�TS���<��x"� ��� ����l�dt�J���D�o�~��>�H,��e�>+�>6v�=�G�>��>�/��B˄>�}>�Pq>��>��S>�>��>qV�<���d�A?+���l��$�뾲
��&E?���?�e	?�/=�r����F�5?ƛ?#Ơ?�9>��q��E�r ?7�>�q��r�>��>��>ó~��kҾd�N;��c�k������>�>�=�2�w�T������>��?�|=�Ӿ�\��o4��6Օ=��?z�??k9�
\�J&r�AoV�fr'�M��=�x�'rž73�]*m�������h�m q�@�t+R=	�*?c͗?����ž�9����~��O�㞦>H�?� v>�l�>��Y>������3�A�h���(��JZ���>��?�΍>�fI?�&<?O�P?[WK?A��>���>����>��<(^�>���>�9?��-?�[/?��?��*?��`>����(���ޮؾ?Y�?N&?��?�\?#셾�ɽ+���3i���}�B�}��~�=���<��ӽU�q�l&J=8�R>��?����@H�A���Ƹ=�GM?�#?!�?�+��Ǔ�Rؾ A?��?p�>|��ƨ��x�6�ul�>�bA?���e�G<�2w>W�><�9�e�����>4�=�#P�)�����y=+̎���;陁>H >PE�=�n);H�=[Չ�C@�>��?���>*�>y䆾�����G�=�Z>��T>��>X�پc����&��E�g�Yy>A�?X:�?gh=���=��=ꖡ��5��gy�#n�����<��?ԫ#?��S?H��?j�=?�b#?4�>Wl��P���<��>���=?��)?���>_y�qľ�o��2�+�x�$?a�?u?W�����="����ώ꼟<G>�.�w�{�^访�A<���F�����8��&�?b��?��y)@��D��+K��Oʨ��G?$�>rƑ>��>�g+���i�a ���F>��>�WI?QN�>��@?E�y?x4]?��\>^]/�ɵ������M�>�)>NL?�!w?�>�?�~x?�6�>�\*>��&�XG�����ͼP#-��8�����<�-j>`��>���>oֲ>$�Q=�檽���GCF�6Q�=}"e>��>�^�>ܶ�>:~>ʉp��B??N�>G]Ͼ ������������.w?��?�$?�)<"^%��AJ����l��>dө?86�?Bj?>yI���=f�>�����29��Ӕ>1�>�>ZJU=�(�=�;>�"�>���>����+�g�>�M����?�&M?�� =j�ÿ��n���J�������]K����o�O�����T��!�=5ϛ�8��7w���*^��ܥ��E�����ʙ��8k����>�=�\�=?Ƕ=jS�<��
�R4<]Tn=��<%��<�==��H&�)b/�祾<=�u�R���}�<��r=�.<�̳�q�m?K*N?�9?�?�>��:>h���i>D������>>8>������ྐྵQ��	T��R6����Ծ����˪e��Z��$$�>��μ/&>���=��}� � >B�l<j��=�==Ջ��e����=��=|��<�]H>G��=L�D>�c??�=~��<���#u���7=�q�>(��=��n>��	��]?��{=���}ÿȝ���?���?NA�?�|�>CJ����>�h�����]�~�"��&>惁>G�b�P7>�k>�Q�)���Ȣ����?H�@SMi?�H��U�(l�>y�,>�&>��S�O3�pvV�8Cf�� V��!?��=�V�Ͼ�}}>B��=���d}ƾ��=�J>�܍=�*�zDY�n�=
5u���N=f}=�ن>=>��=����=�\@=�T�=�L>u֯;m&)��&�i�=6(�=Ʃa>v%#>�W�>L�?��5?p\f?�/�>fl��/�Ӿ�U����}>9�=���>#�	=�<+>Q��>G%?��7?�5F?���>ҍ�=,��>D�>i�4�Uu��޾�$9��ּ���?�y�?F"�>�Ȩ=*0#�F�i�E�I]P��?5�/?e?���>(X���࿵R&��.�������H�fe*=5;r��bU�U���va����)�=�[�>9��>��>uCy>�9>�N>��>ǳ>*~�<P��=����<Ny��b=킑�u�<f�Ƽ#��	 ��c+�C��&m�;z��;B�[<���;������>B۩=]h�>�FE���rN>,���_~;�;$�=�:�&�S��>���!��� ��gx�J>1�=I�C�b���D ?��>.�[>���?���?��%>/Ef������ւ�������=�j�<��h�ѧ.��h��[�Y�����"��>{g�>�٧>���>ӌ3��
C��6�=
��,����>��a���m��1�i��뤿�����g��J����=?�#��o�>Ww?��G?5e�?�\�>����Z޾!,>�+z�K
�������d���g�?9�$?�|�>!1羐�<�	þ�Y��ߵ�>l�|�M�����/�i���U0�>(��v*վN�/��\��{��/�?�%�a�T�>��R?EԮ?�@����rS�a�������p�>P�h?J�>t2?,�?����u��0��o^�=��j?���?���?�>�^�=z0��r��>�S	?兖?�2�?E�r?�*?�H��>2��;��&>���A��=�>>R�=t��=0�?��	?�
?�	��#f
�rX�f����[����<0@�=2�>O�>��r>���=4	b=�ۥ=�"\>�Ҟ>ϐ>ld>�x�>Iˇ>��)}!���?i��<�(>�,4?�NJ><�`;1�	�Y���T)��Im�$���Trc���`=L�>��<��ͅy��?,X�#�?��d=��.�V�(?�Z޾�=fe?F�>:��=�"??�>�e>	>�g�=����A�>{��=�I��d�=P*��<��>�:�K����$��>���G��D2�׽�p�c�[���
���h�_��+�ཛ=K��?�㖽�'��ޫ#�=�;K� ?�@`>»?�C���?����2>Ig�>�&>Y)���<���[D��^�?ΰ�?p8b>u��>�EX?�(?�X3���5��#Z��%u�J�@�j{d�*`�ⳍ��E����	�
8ǽ�^?//x?m�@?a�<m�|>Cc�?�%�x6��B��>/��2;��7I=q�>0ï�PK[��Ӿ�yþ����G> o?��?*�?�rS�D� >�F_��W?�pC?"�?�� ?�!?uC�����{R>��Z?wׄ>��U?�N+?�m�>���>�k�=����
���\MսR���*��,��5��;��<;��=�s�=r]�� �ռ�J缀�ܼwK���i��Y;��}���=C}�=�N�=ga?jj�?���>��2=�mO?�"
>h@��&���l?3�?k���Z�"�8��������A�� �?|*�?]�?DC�>���q꽞�+=\��>���=���=~�>�T-�j����R�<_�A<:�Y>7c}=p>q=�1O����l��e^�QF>v��>o7v>�#����>�������Og>�<�ܿ���L���G��w8��Y��ӂ�>��P?��!?��=�d꾓J��݅c��D(?�g=?DP?�os?���=:cؾ��:�f�>�`g�j��>(��<DH	���������6<��)v�Dׄ>+ǫ��٠�gZb>;��l޾Q�n��J�����GM=}��PV=K�.�վ�(����=X1
>����� �q��kԪ��-J?��j=q��FiU��p����>���>��>��:���v���@�ݴ���E�=1��>��:>��������}G�05�D��>6�D?'�`?���?mˁ�`Xi��=�3P�3��{��A�?���>я?b�D>P~�=����*��?af�C,B�
`�>M@�>���'fF�l���L���^$�ߙ�>��?��#>}�?�O?�V	?!�]?f&?��?Z�>U{��g��VN&?��?�.�=#�ѽ�0R���7���D�Z��>!�)?bsB�lp�>]�?H?K3'?H�Q?�?�>E� ���?�YM�>�8�>ݱW�Aȯ�a>�IK?F)�>S.Y?7w�?,i<>f5�����<���Y�=��#>�c3?$e#?sJ?�W�>���>�o��/�p=�"�>�b?Ur�?�,q?�|�=�5?�+1>��>�Ŧ=��>�$�>[�?�O?!�r?H�H?s�>��<3��������y���@�LI�;n2<q~=���$�z�վ-���<���;9���=!����X�>��W��B;��>�
t>Z���Tb4>��ž�w���A>Z��&������`J9����=�~>,�?���>�&����=�ߺ>OU�>���&?33?8�?�F;�`��Qھ�eP��'�>��@?�{�=��l��f��Zv���m=¿m?��]?�W�������Z?i�c?V�������ć�� ���u�mJd?\?��8��M?�}?[?
w?a˒�l�K�����ʄ\��u�T@>�Ӧ>�2��@7���>4d?�?t3�><��=z��q�g�F^��)�?�݅?�}�?�Z�?�s>~5U��mͿc��ZK��7$^?���>ȟ���"?�����Ͼ�p��𘎾M%⾜ت��(��������{2$�XՃ��]׽�x�="�?�s?h�p?�w_?_� ���c�`/^�y��V�%�����e�E��,E�\C�ֶn�qt����2���kH=NTw�g�n�2�?�%?�[���?�[}�c���k��vJ�>+�Ⱦe���b�,=�sɽ|�<]��=��н�\���о&S?��?�U�>FI?X�:B:�	�Q���V�/��>���>���>���>�|�=.���H�S��^ؾ)�Ӿ��ku>d�b?<�K?�n?���0�ˀ�~�!�B�7���i�=>;&>̘�>�DV�!���%�C/?��r��>������
�+�=R=2?�z�>]f�>zD�?�|??F�𛰾kE��C1��;�ɲ>��g?>��>���>��ɽ ����>��j?e��>���>5Z��ܡ �
�y��н[�>���>�h�>�q�>
�/�
V�$@�����:z8���=D�k?c����b�O$�>.�U?r1���6:W��>�+k���#�. ������->>�?�ߡ=��B>Ofþ��	�a�z�?��ck8?�C? ����^��D�>y7?�>?��?Nkt?�Q>�AA����>�F9?�q?9څ?� ;?�/�>�^��	S� �&����N��=�=[=v�>U7���>��.���!X��&�������=��=�H�=����%μ:Hڼl�<�Qۿ�WK��(پ|��y��M
���H���?�����ߴ�h����x������(���U���b������=m�[u�?�^�?�������6�������a��$ɽ>��p�s'���[��������4�߾�謾}�!�"#P��;i�Ve���%?@�����ǿ�ԡ�\�۾~�?�?�Ly?����#���7��s>�C�<�j��ȏ�1��k�ο$i��c_?=w�>B"������>z��>.Y>�n>�l��'���L!�<1F?
�,?�-�>�cv��-ɿ:+��߼<���?:@�A?��(������U=k��>��	?�?>�Y1�'.��۰�sB�>�?�?��?�ON=��W�D���je?<��F��[޻:��=���=��=���bJ>�b�>!��M|A��vܽ��4>>Ѕ>��"����`W^�6g�<s�]>��ս<���5Մ?,{\��f���/��T��U>��T? +�>R:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=u6����{���&V�|��=[��>c�>,������O��I��U��=�˾ƿI�$��~��S=�)Ӻ�F\��o������T�+$����o�7�轾[g=���=(�Q>���>�NW>VZ>@dW?��k?W�>�y>�q����wξi/��7��|��������c���8P�N�߾~�	�������R�ɾ�Q�Hz==JX��f���p�fzc��PG�Ϗ-?V#l>bb����J��c���?������5�T�l�n��Zؾ(��s�W��?� .?\�����`�\q��Й�n�'{R?��սO��4̪���=,�����<�r>'޶��X��td!��q8�W�8?�?T;����<7>�����<��"?�b?%b=GX�>�2?W/��}���>��=TN�>/V�>_�O>������@<#?B�^?,R;�2�����>yW���%��%��<�)'>f�7��/��XI>aP@=�.���뗻��������i?�He>υ*��0���ֽݕ*=�*��k?a*?�@�>�wk?��E?ڃ>�fȾ�bU��(�lj��bS?E~?��@>ߍW<�1�����.Y?��{?ٱ�=�2��z�Ѿ�:����9�o�5?�l?��+?�d�������u����bX?��V?�h[����3�k�3�ff>ɛ�>�O�>�@9��w>v�"?�ό�q���¿��"�ӹ�?�3@Iu�?N�����¼�M�=�?��>�j���:ϾY��;ɱ��v>lE�>Յp� �d���{�5v%?w$�?wG�>��T�4��#��=v&׾³�?�v?d���}�T������e�����>t
>#bg�@����@����5��_��~�쾭Y��>{��>7@�hh�d��>�>��������s�����E�R�g�*?��>�Ž�{X�oEq����	H]�W�R�<��4�>��>Ze��`D��`>z��<��D@�/��>�6ɼ؉>*^>�8F���Ӛ�~T�<�x�>��>eـ>�ս����/��?cx�ο�V���� �� \?Π?�?A?ܠ�I@u� �i���B<�I?"�v?��Z?�+�#�_������s?F ���`��� ���6�G/>�S#?��>�%��=�m>
�?G|�=��Ŀ�e���6��*m�?���?�5�g��>|�?A�@?H.&��;��va��)#�����w)?�p^>usʾb�9:7���C�Z�?R�'?K��2D1�_�_?�a�G�p���-��ƽ�ۡ>k�0�me\� M��2���Xe����X@y����?Q^�?^�?��� #�Q6%?�>X����8Ǿ��<���>�(�>*N>^G_�M�u>����:��h	>���?�~�?Cj?���������U>��}?j5�>"�?x�
>F�>fw=z��&<�<��><w�=7Q����? R?�K�>j�=��H(���L��R�� ��7D���r>e�\?}O? �t>������K��*��$��y,>�޵�p�,�0ؽذE�/8>4.1>�@>��)��ʾ�>���N�ٿb����aݼۋ?0�<p��>R�ƾB�Ѿ���=�!?6�Z>�,(�������´���?���?�?�Ž��`=��>���>a��>�\��v���Ǿ��>!?S�;��'���������>��?�@���?�~H�_K�>Z����|��]����W�Ow�Ǻ�4N(?=���h(=��>ć��	�t��<��"	K�̗�>0��?�[�?���>�R?�aI��9	�]B�=���>��??��>d��=l��Nd�=���>|�F���m��E�Z?N�?p
@�DQ?���~����Rs�崢�J3ƾ��=�N=�w>M\�֛/>a&����ѻ��L�i>�u�>�K->v*�>��1>��>�e9�@������Z^��f���xwA��)(�J&7��Q��Kt��V��\��Gľs�վ��
���n��8�H����=�p����>,!c?VSz?6��?��>��T>Ԛ>�(��r�=/�;�>'�~�>��$?�#?X�?Rv>����s���>�ot��) ���>��=GȦ>��n>�Yy>Y+�=?��=�6�=�W>2#�>�����̀�W5>��>F˺>��>>%"<>�>�ϴ��2��9�h��w�r1̽  �?t��A�J��0���;��v����m�=�\.?�v>����;п�����/H?y����,���+���>��0?^W?��>���U�S>>����j��X>�= ���l�.�)��/Q>�r?��i>Atx>��2��)8��=P����Ȼ�>h(8?�u����9��<t�uG��b׾�U>�O�>rqP��[�D	���v~�e,j�f�w=;?_�?����̏�� �v�3i���VI>E�_>xD+=ײ�=�L>ҝY�pϽߌF��$"=���=Fp`>%?{,>�*�=�t�>$<���[M��Щ>`�=>�9,>�??��#?�@��ԗ�����_�,���u>�?�>��}>6|>�J���=W^�>\a>��銀�����?�ЋW>�$|�b�_�|��u=�ۚ����=˕�=�6��4�<�9W$=�~?�~���㈿<�`^���lD?�,?��=��F<��"������E��[�?I�@�m�?�	���V���?@�?�����=Q~�>�ӫ>�ξn�L���?��Ž�Ȣ�h�	��)#��Q�?��?V�/�	ʋ�wl�4>�]%?��Ӿ-D�>���Y��@����u�~�!=0*�>�6H?�����SQ�5 =�\[
?7?6A򾜫����ȿ#ov����>���?3�?��m��8���@���>���? !Y?i>RP۾��Y��N�>��@?R??�>S(��	(�P�?�ڶ?7?��I>�L�?�s?g��>ψt��,��I������2��=�}<��>�|�=)c���qD�rm��Cʈ�j�����'a>�m%=���>�۽�껾9�=漏��˦�]�U�L��>�p>��K>(e�>4�?d��>cǙ>��=n���h�����ÄN?,�?�����d�l�<��X=QkC�P�,?+=?�r=�밶�N.�>�x?��?J/t?v$}>|�+ ��g���1$�����;�d�>��>֒�>GF$���*>�{��E��D֠>T��>�t���/���K0�hث���>y2?��>T�=�?T�?
nP>j��>�\�5Ò�N#��d�>T}�>�&?v��?N2�>$︾��#���h��lmL���=^U?�@?��>���U����>7B�=�üx��?h�p?�����8?=�?�u?�7a?\�I>�V�ϫž#��;���>�`"?���E�A��7$����G�	?	?�|�>{2����ֽ����h���S��&?�^?rS&?��Da��¾92�<*!7���V&;�M� >��>̀�N��=�>���=�`m�q�2�Ze�<T��=:ڏ>���=}7��5��Ϳ�>i��v�c�Z�c=�Z{���g�N�>��7>|�����,?�Խ�O��Vⲿ������\��O�?K�?�ء?����2�W���'?�ņ?��?�Ĥ>�����F7��~�T���'F��!��Px>�M�>��>>^��%��_6��)Й��@�O.���>���>�%?!�>g�>��>�����F��I�4R2�TW���'�P���M�A��R͛���]�>�Ľ�Ҿ��U��,�>W啽z��>��&?�K>P�+>��>�=z�>U�W<	��>Kɚ>U>�> +�=4g��!1�z�S?����$�W��Le���=?�@m?��?�YN��E��r���� ?���?J�?�>�>p�b��*�m#�>�A�>hW�}�?Aѧ=��
�wMӼ!�ž��4�>�5��<��>%���D�?�iYB���C��� ?Ĕ?����о�IϽ8�����m=�.�?��"?Wh?�U�J�t�O�"�L�<I�s��=~۽?����*�39d���z�x�o�Н|�F� ��{�=!:7?��?\T�iT �͇��;Qh���K�|�>P�>Ԍ�>�i?��=�~�������f�L�-���f��,�>eVn?:
�>�AJ?�o=?��Q?[�I?��>�W�>ٲ�ٴ�>U�a<o��>m��>�9?x�+?E�0?�?�'(?�T>�������׾ '?��?��?�v?� ?����Fʽr���������|�I���@&[=w��<��ս5�_��d=pQ>aI?C��A�Q�7�VS�>�^A?�'+>=j]>��U��=ȗ���"?j�>�z�>��4�.���4���>쿢?�_>;mo7=ͦ�=�S�>������B�aہ>�>���Y>���6H��S�=�F���6>���㑽�^��	��,�<��>z#?gʉ>׏�>UɆ�.\�Y��'��=I�X>�lP>N�>�ھܨ��NN���Kg�n�|>��?�ô?$�W=���=���=�垾B����b��1��|e�<޹?�$#?uuT?���?(�=?{�"?S�>�B�{������P?1�+??�>�Ͼ-q�������7�]�6?J&?�n����Ծ����4>�w�>��ξ�KV�-�g�U�/�ڻ���YY��[h�?� �?%�y�+����c!���R��n�G?1��>�.�>ܵ�>@yD���l����()�<���>6T?��>�cP?��{?�k\?ʜU>W�5�O謿�� �����#>+>?Uр?^��?�x?��>p�>}�)��v�z����_�DP�`Q��_�M=��W>JB�>�S�>��>
�=v1ʽ�T����7���=��_>�[�>t�>V��>��x>�/�<��G?
��>!`�����I褾?у��h=���u?���?I�+?�"=���[�E��X���H�>^o�?���?.?*?��S����=�ּԶ��q�/�>�̹>n8�>l��=��F=Lq>��>���>s.�EZ��o8��M���?�F?���=��ƿ��o��C�,����=�z�VL��Eٽ6J��(�=tܧ���@�[���A�e��]�l�Uy���Z��^����>�C����=��{=M1=L�&=��_;�oK=� ;w��<3!��i{Q=���<e1��i��LW�=�i=K٤<͟�<oʾl+|?ēI?�T,?�A?�dy>�� >��M��|�>�y|�H]?ȉX>C�Y�g1��Z�2�^����瘾ڡھ}�Ӿ�Y`�lp����>�)Z���>��2>�8�=�ɑ<�$�=�o�=e�=�Y��<�<��=�ó=�?�=���=�N>��>�6w?X�������4Q��Z罢�:?�8�>k{�=��ƾo@?}�>>�2������{b��-?���?�T�?@�?Fti��d�>K���㎽�q�=W����=2>z��=z�2�V��>��J>���K��E����4�?��@��??�ዿϢϿ4a/>�\<<3�:�dQ���5���3�
5���JȾ��#?�LL�9F��ܲ<�a�+����"��w�=���>-��>�Ij>��Y���=��Ͻ���=�s0>�@�=���=�J<>y�Q�&z6>`��=��*>�w�=G^����2��%��lh> �=@j�>��� �>uS?�U2?9Fd?��>־`�4�ǾH!Ǿ�ʀ>#��=���>3#�=C�;>�	�>E�8?�D?�G?��>�=�>�T�>".+�Ymn�H�\����c��ۯ�?�,�?K��>on=�L��
���9��޽�?f�1?��	?��>�T����R&�n�.�:U����6i+=�wr�/.V��c���y�]�㽌��=�g�>M��>��>�Qy>��9>ɱN>��>��>A�<�O�=c��T�<�C����=y����-�<��ļg��f����+������;���;HE]<?|�;(u��DD�>cF>���>��<rKʾ8`>C��[�Z����=>I��@E��q�C�o��L%���
���S>��o>,� ��a�����>ќy>�;>�#�?�ȁ?��J>S�7��y�&���L����P�ޮ.>�[>�=�S>6�l�Xfo������ ?{'h>��>M��>ӏ&��n,�v�#=��	�Ħ����>��K� ��=�����_3��������]W�d�ּ .?�˅�����3)�?��R?��?,
?Zp���l����=C볾��eM����t�'�S�3?��R?�2�>�%�C_�y~˾o����>/H�ĽO��ᔿ��/��1�ŷ�(�>����Iо�[3��셿s�I�A��Ju�ㆹ>Q�O?�?Qoc��Ӏ� fO�����s�����>��g?I
�>�>?��?�䭽�a쾔��7͢=��k?�?��?�T	>Jp�=�?�����>O�	?�'�?���?(s?��D����>�ۇ;w�>�n��\k�=�>.�=,Y�=�?�F?��	?#k�����s5�ץ�jh_��*�<'�=�F�>�>��s>���=�U=��=$�Z>��>)u�>z�f>���>�>�7 ���P�+^-?��=�%c>�,8?f�=>�@估�Ⱦ�Z���f��ǳy�L�%��<�Qý�j>v=*>Yr�=~x�]	?�Ͽ��?g4�=��#�Gc	?9�	7e=�?�>�k�>,�"�-��>�B>\�=���>S�>l:�>u��>�w�=�<�Z��=�C=���M���3��(^�C.��S_�>�ӽ��������D�2�<������s �ܜ]�|��K���.={��?�'-��Wh�7�
�a���>�U>@�?`殾��*�P�o>g��>��I>����ݑ�G<������﬍?#��?��^>⫝>��U?��?�p+��95�V[��t�޾A�Dme��a�%�������������^?y#z?�`B?H�<��y>��?u�$��Ӎ�>D�.���9���D=~��>�V����a�:Ծ��þ�J��6F>:�o?c�?]n?=_[��zɻ�v�>�N?J�I?�c?�Q7?��9?Zc��?7�>j,�>č?͏;?ߊ?G?�?�>���=Nn���������H^�n�۽Г⽿�׻$�=vF>=L������R��=��=�DϽɧ�<��8���e���)=e��=���=W��=z`�>��[?H$�>#/�>�6?Z!���8�'���6.?��&=X�������9v��"���H>@yk?�v�?L\?�P]>l~@��A��>�1�>�>��W>ٚ�>�����@���=�N>��>�=��@�n�������z��w��<~G>���>ѯ�>����i�?>�7žI[���Ǉ>�4@���Ⱦ.%�S�0����
*����>P�M?r?�����<��ėC�P f�B?<�7?�IV?D3x?L��=p��.Q�\!4�m��]Di>�,�=���i��iS��u�1�	뽼�/�>���۟���c>;����޾g�n�C�I�d���\=E��� O=�d���־��z��#�=�h>�i���� �2:��㲪��I?��i=�ꤾ��T��9���>ď�>H+�>uD�Ur�Ր@�񄬾Yb�=�Y�>F�;>�)���\^G����S�>�!A?��`?��?�ޅ�c�\�2�r�	���|��5[�{�?2H�>**?J�A>�і=t]�����N9d��N<����>���>�����G�:���K���!$��΂>s��>�SE>�A?ݐC?�G?yXb?_�2?¬�>�ʐ>�d����оwB&?��?�=��Խ��T���8�F��>��)?-�B�o��>��?#�?F�&?U�Q?z�?;�>�� ��A@����>�Y�>��W��a��E�_>��J?���>F=Y?�҃?��=>ʆ5�\袾�ة�"Z�=�>��2?z5#?Ӯ?���>�}�>@������=��>c? @�?��o?�O�=R#?��2>���>��=���>ͮ�>u ?�`O?)�s?a�J?�Z�>�i�<Eά�������r���S��Ì;��K<<�y=����t�m-�q �<���;������������pfD��쒼I�;���>�s>Ձ���D5>��ľ������B>O
˼��� C��d�<�~��=�!~>~�?uɓ>�j"���=���>��>�����'?Z�?��?�Ȑ;�ya�>پg�N��}�>8�??{y�=�&m�Iؓ��v��ve=�6n?�w]?A�Y������Y?;�W?���6�.�~�������u��g�f?��?�����>uz-?�7�?֚=? %|���w��@����{�wdW��.'>�ظ>�<�X�e��E�>7�C?���>��?�w[�$������־�Q3?� �?�۳?��p?�]>
�n���ѿyM�����C�]?��>� ����"?��߻_о07��R�����a������씾J`��$�bd���(׽���=6�?�!s?�q?�~_?v �W�c��]�����U�|W�|�&�E���D�-jC�s�n��b��(��v���H�H=8l��Y���?}�?䇆��|6?��6���0~;DbV>I�$�<k.�;�[%�0D�=�y=�,����ٵ�� �?���>�K�>�/?�Zm�&-�!]���3�+����s>���>��>$�?�T��˖v�<���D���������l�q>�a?��N?#o?�R+�Fb1���n�R/$��a�Q7��_>��=B��>jL�ݤ�
�$�+�G�f�n����f������={[,?���>�5�>��?���>3n��}��;����;���C���>}Q?<(�>6�>�ㆽ�W�of�>i?�`�>l��>㈾�#�Js��^�����>���>�>p��>��3���X�����Ɗ�d8��t�=�7i?zd����Y��>�+R?:y���)<r�>H��֊������.�R��=�0?8��=x�;>�F��'_	�.C�~5��i�*?��?Z��ā-�
�>/,#?,��>�s�>6/�?9W�>�žĻ�<�?h�Z?ǽI?�`>?:��>yC=�]����Ľ�@$���:=
��>�wV>�gN=_��=����LQ����̷=�D�=�4-����+EN<����2�<��=��+>kvԿ�WF���ȾԾ��g�۾8$�]@�� �ļ|�����q�о��ʾ��J�#��ֹ���lw�����IP���)\�2��?�@�*c���־8��s��~�m��>8�?�XP���U�Vܷ��5��5;`��T���[��8Y�&M�̔'?^���ֽǿ"����9ܾ� ?�@ ?+�y?����"���8�E� >B�<�-��f��ٚ����ο�����^?���> ��7�����>B��>&�X>8Iq>����鞾�2�<��?I�-?|��>	�r���ɿ���4�<���?=�@��A?%k(�J	쾃�X=���>�	?&	@>(2����/Q��,��>�Y�?֠�?�K=D�W�(���d?CU<��E������=��=�?=���4�J>s�>����G@���ܽ&�2>�r�>E���*��S]�@)�<�]>3ؽTS��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=u6�񉤻{���&V�}��=[��>c�>,������O��I��U��=�����Rɿ��$�&��6�=��o<F&���`��N߼grl�-�ξ�Ɯ������S=y,g>�7�>{�g>{<>Q�@>h�O?��|?*�>g��=��1�A����D׾�)2=V�*�	z(�{�j�7A��ի���ؾ���Jx2�:�'��b�����)=�}+�=$R�8���� ���b�A�F���.?��$>u�ʾ�M�uE%<�KʾU����f��E�[̾��1�!	n��П?�:B?��Z-W�
��{��h����W?kl�,��M����Y�=�j��XT=Є�>ќ�=�����2��YS�ه]?!�?�7�����}�>�T��sM�[u�>��-?�?�>�>�?�ֹ���?���>����r>\�?��?����xCZ��_?�[y?���)4��.e?b���v���a��s�>#{�����|�>vN����������\�zdR�Va?�a�>j�.�{z9��ި�C�.=��۽��v?I��>�4�>iRm?��Q?a�=e�:E�i��o� ;2�R?���?�	4>�<�aȾ����WX^?|݀?�b>d{�f�վ�F��,�_�I?p2V?�I�>v�=QR�%~��KԾP�H?�Z_?��%��Ц�����<z>e�,>&�?��?��Ԟ�\(?��������w����$��_�?'@ ��?�8P�f_��r���?|'�>��������A�Ǥ���	>��>?���xU�������T��?�w?ϩ?_�c��r��X�=�6��ج?O�|?�Y۾ū�=$�ϓh�v��[-�=�o3>Kr=<��F��!1�o�˾խ��"��]wU��D�>��@��I�S)�>r.���"�d¿iy��l��b%�!<?k��>���<߄��n>v���z�>�Y���Q���F���>8�>�b��X現��~���>�G@�d��>|�j��`�>��E�(ݵ����ֹ<r��>|��>��>R�ɽ{~���0�?���+Ͽ�&������^U?�̟?9%�?ϯ?a������S����t�<�hO?lr?5�V?]�
���r�~%?���j?���z�_���3�oE���S>�/3?$��>p-��@�=`'>� �>��>.��xĿv涿�_����?=L�?n�꾨n�>H��?Z�+?�������Q3��r%+��-���@?�3>N4��3!��<��䒾TV
?}/?���OA�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?~��>P��?d�=rX�> ��=Ff���/[>$�>2�P�
� ?��N?�)�>Ϊ�=F?�$P-���E��>Q�_��qC��O�>��`?�K?�}[>����e.�|� �m�Ľ,�2������H���#�ֽl�:>y}:>�>�G�Jzվs+?G��Ifٿ�]��p<;���>|��=�(?�p ��X��=�D?S�.>���A��Ԓ��=����?z-�?�?�ľU`!�>VE>��>�_�>����<��,�����>>Y�$?c{ �LY��d@{��X�>���?��
@2��?�I��'?�L���|��_���1{�z����\���7?;��Mi��z�>�^���������Z��#�>E̷?��?���>��V?�yZ�*�!�V[o>�8�>�Q?���>矖<�V较��<'��>�s �����u��M^?�	@�@�!�?I���TRٿ#V����Ǿ:����=2�=�>FI��پt>Z�=}�]<y�<�rM=��y>�}�>3Vk>�(>���=B��<��bc ����� ʐ�v%@�hd��t�#�f���꾇�^��:�Zݤ�|̾\GJ�}�½`=)�Wi�\D@�%��<J�>�MH?t��?|K�?��>�wO=X�>�ZF��O�=ڿ�;��=���>��#?��7?�S?���>�%���oE���r��T��6�D��6�>���=�*�>��e>���=q��=�&�</�>U��>�8��z�=�{<x0�=�m�>d�>�
�>U�$>��<>�4>O������,�h���v��Bɽ��?Ͼ���J�0��]���'������=�n.?�}>����3Cп�歿�H?*唾j���+���>��0?�3W?H*>����R�6>	����j��A>H���o�l�o])�قP>�A?���>q7�>����Y(��-`�Pd¾�{?၇?��)��R���틿8F\��^@=4�?���>�����>�����vi�#9�Hn�:?���>��[����)�56����=��>���<�7>4�<�P����,�~�	�O,;�u=��c>�?�j>� >4<�>`����J�Y.�>��=Y�e>�&5?�c?fY>�J��I�����K�:>F��>;�m>�F>��}��z�=�{�>�R�>�X;���2�<��� 0�� �{>�S%�of��Vy�դ�=9*��j�>�e>M����q�[�?;�~?w��䈿��f���lD?�+?��=^�F<��"�J ���H��L�?r�@m�?��	�ƢV���?�@�?�
��ܷ�= }�>	׫>�ξ,�L�ӱ?D�Ž�Ǣ���	��)#�GS�?��?�/�?ʋ�*l��6>�^%?˰Ӿ�N�>^9��/������ô]�I���6X�>b�I?ކ�{	�T����>�c�>5N澛/��=�ʿd-q��\�>7�?�"�?/�^�R����jC�
	?���?��S?�n|>3w�2�G��`�>��A?1Z8?g˓>�%�L$*�Ev$?��?tC�?��L>�)�?G�s?��>�񂽰+��s��81�����=���Ý�>su>�{��=�C������O��ޒi�6���md>��=�Ⱥ>��ݽ-��pæ=E���D��ڃh����>�#w>�L>X�>��?���>���>
��<R���Os��� ���nL?���?���B7j�����9�=�D���%?�?���lM��k>:u?�M�?��]?+�B>�c
��۠�K7��]���+�;H[>~�>1��>_"���5>B���ș�M��>y�?>�1�t��qCy���=86}>^6?V��>�=<�?�?+�{>���>.�_��j�����-��>c%?�G,?��? ��>�w�W������WP�L�*j7>7)b?ټA?�ɳ>��j�	e>�9������?iyZ?��Z��p ?��`?-wu?� G?�s>2�X����ȢF�b��>��"?\����@���%��� �&.?�[?v0�>ߠǽ���
X��H���߾�w?ã\?i�?A��gf��7ƾ�X�<��[����;0�<�H�>�>h0t���=Ʌ&>��=�h��Y?�Y&<r��=F!�>�~�==�;�溊��p)?$:pV����=#s��:8�r�4>��<> ���[?���f�z�_g���R��3΄��{�?���?�a�?�[��5Be�F9?c��?��?���>��������h�u�t���R�8����C>c�>}�Y<�t�ǫ���_���Ȃ�S5�� �
U�>(��>!?�X�>��5>�V�>K�Ӿ����+��u���1]�}�eh �(0�l@�����B3��'�<����.����Ks>ḽ��k�>�]�>J�>�R!>�p>ꢥ=[��>�]�=��}=���>R��=T�>��Z>Y�g=N=b:]R?.���@'��g꾿�����=?�<h?��>[���愿��	���?۴�?ෞ?�ށ>�Xi�/M)�Y��>�9�>y8z�yY?�{R=�y�Q3^<���E��y�t���d�6v�>��XW6��L�Kf�+?�?	����̾F?ؽ�]���6�=Oh�?�1??�&� TP���P��\��@H�Ҍ̺n����)о��#�Y@X���:���0˃�W
��*�=ǋ0?�\{?/������䓾�cu�C�T�䝏>��>�p�>�?ZQ>����"���Y�(�!����ri?�&g?܈>FG?$�G?�g[?|�H?#�>W��>��Ǿ3��>F��<K�>)��>7�8?y-?Ч8?w!?σ?�@>@,�"$����վ"@?J]?��?���>�[�>�Zv�L�Ž+���F�����j�t�G	�=� �<����ke�G=
0d>�d%?�����7����2�>A?��>i��>�Qe��L�t!<ܦ?��?cMN>m��,h����ŝ�>��?9���uj=�V;>^�=G��<�iN<c@�=���>uZ�=��a=��T�0��=P-\=	��<��0=�W=��<��>y;	?�)r=0�>�}P���Ҿ/69�V>=����v=�>u�=���h����]�'�>d��?���?�q�=ɪ=�=V���C�p�s�9�[�S�K�=�H�>�Z�>z��?qM�?;�!?��(?R?>��i�������=���?P`/?�ߥ>�,�1�Ǿ�8��L� ��r$?X�?!dy��^�O=5���þ��=om�>�^׾�{r��꧿��b��>�׏�󵇽I��?��?kP��?%�I�����b�ؽ�$/?ݠ�>]��>�x�>a^O�k�I�'��&��I?�H?1C�>o N?���?�[f?��k>�0��¨������D<G2=>��B?'v?�~�?�r?��><_>��'��_ݾv����K���׽}�k���=� c>3o�>���>��>���=^���f'���F�Bz�=fr>���>J��>���>T+�>ٞQ���G?���>F��ş�٦��� ��c3G��~u?�8�?/e*?c�=���mF��&��m��>�h�?wL�?c�*?��U���=ʿݼ�޵��sq�	�>[��>�>!��=�H=�>Uf�>>�>���XE�C98�t!L���?)nE?��=;ƿb�s�Ƴt�p���í�<�s���d��Β���W�m��=i���$���k��`�Y�C����̺�������	}����>-�=���=t��=\2�<Z#��$b<��H=+�<h�=��u��WT<e�(� )������F7<�|Z<4�C=.N���ʾg;z?�C?�$?��C?�M}>�>��[����>�>C?�^>������ʾ�P�`y���n��a�Ǿr�8�p��w��&�>��K�*M>�>"��=�<���=�=��m=�W5�h"=(��=���=���=���=�>�>�6w?K�������4Q��Y罋�:?�8�>�{�=��ƾ?@?p�>>�2�������b��-?���?�T�?[�?�ti��d�>T���⎽�q�=���>2>P��=��2�:��>%�J>����J������s4�?��@��??�ዿ͢Ͽga/>Gj>�O>�zI�/M-�����?� �B�}?x�D�Pv޾d��>0��=����]ﾈ��vi>k��=0c��~e����<�սOW�=z�>=nB�>�%>jէ=�y��K%�=Y��=�0�=so0>,�;�{��;��eP�=��=�~J>��D>�H�>f�?n�0?0�d?$!�>Z�m�N�ξY9¾�9�>���=�)�>]��=q�B>�z�>�38?�E?�RK?�}�>.<�=�]�>ئ>�,��8m����A��^�<���?���?�q�>c�<�7C��V�q>�BjýjO?�71?)�?ҝ>%r����uc5���־{�>~�>�7���:L�s:м�H�����+��>X>�d>6"�>���>a��=P,X�3C�=,{�>¸�=_��$#>�^B=�V	=����k�=3X�,3'�����B�w�=�����s�=�N>j�@=rv�<��I<���=�*�>���=���>�t�,�m�nN�=�P���f����=�"��+���b�����h�F�E0��]��>��>��z��N��FL�>�P>�U�=���?FX?h�>x�#��"��������^��M�<�>=ܫ=b��+�M�q��/�E�1z�>�ew>���>�	�>t�$���9�=j���R
�J�>��:���6>�Y�>C�n��Iە���_�TK=F6C?aą��[�=�?	\?��?���>Zc���
���>n�վYG\���$�M�Q�̲B��?qL?t�>+��#-�v����������>4��dM�{���Z(���(��������>�Ƥ����;�2�H�������,tC����P/�>UQ?ه�?�wf�m6��3R��&	�)꽟k�>�rp?B�>��?�?Kd���FF��B�=kd?��?���?�7>��=$���Kk�>/�?��?\��?��s?��b�_��>FĻ���=��8����=^->q�K=��=�K?M'?��?񿬽�M����-`��^�h&�<��=���>].�>�7W>	5�=�N�<I��=��U>(��>dr�>JNe>��>�w>c��)0��Q2?[��=�\>�)&?��>�B�>?n���H=鎳=�v����q�  ��o�g>�&�=J>�7��>$�Կţ�?YU>5�K�:?������<�ѐ>�Ԗ>��\�`��>��>���>ĕ�>mA�=��=�~>��l>�l�J�_>D\�lH5�b`,�Z�o�@����>��N��җ�������9�Vf#�R磾�$(�3�y��]����+�\��<�L�?*�=ܟ����Y��A<Z��>�h�>�3?举�UN�b�>�
?�E>ց龖��$v��(���]��?��?E:c>%�>��W?R�??�1��3��pZ�íu��'A��e���`��፿�����
����>�_?p�x?�wA?㐒<�<z>9��?��%�+Ώ�+)�>t/�);�oM<=�(�>�����`���Ӿ��þ�6��=F>d�o?�%�?�Z?\WV������V>�,T?xHM?N>Y?��>?^�-?0O��'?�d>���>�x�>��)?)�4?&�(?���>XJ�=�,������9��̢e�����)L�E���%n�=C9�=���!���=w=�y�<���<�H�=%�<�=�!=�G=�GB=Rͫ>ɰZ?���>ht>�Y:?0���a<�3E���},?�=�z������j�� ������=�Bi?C��?��^?ifZ>.0<�u G���'>b��>�&
>�MU>�C�>F����?����=;>�f>$�=W�I�\=��h���獾�j�9�>�n�>�V�>ޱ)=c	g>�n�N`���̀>��z�0U���F�nJ�Y�㻭����>�U?�E�>*��=K��Bk��m�#?8A?,WX?Hp?̔ɻ����nm_�Wi޾��P�cCg>ܣ��j�#�]�������kB(����A2�>��/����"_2>�?&�,Z�}�f�4G#�����7�3=���'/>�'���t��z�y��<D��=)��m���2���c���.^?9�<����&��FH��RX>�I�>�˝>�,�v�U�=�"����40<��>
�>q�;R�侟2X�p��m>�`R?��R?W�o?S"���r�ǹS�~q��Q��O�;_�?��>��?oO�=+���,ᾛ����n� ID�vZ�>]�>cj�x�W� ۾6Ū�BQ��lm>j�?�;>��	?AW>?8X!?YGm?�/?O�?B��>�3����߾�&?[σ?��=`�ݽWiS�!�7�P�F�N�>�*?,@�=�>�?N ?�H&?_@P?��?H�>�����@�s��><T�>��V�6S��
�Z>�{K?<�>(X?�7�?�>?>w�4�}���� �����=P�">�3?��"?�%?���>0��>筡�M�=��>oc?�0�?'�o?���=�?o;2>���>���=���>,��>�?XO?��s?��J?w��>��<�8���7��OBs��O��Ă;�tH<�y=!��03t��I����<x	�;�h���G�������D� ������;3��>��%>��~�g�>mN��=&���r�>1 ��N��A���1V��31�=d��>wp??�>����A>=0�>���>�/�G?�!�>Ps?rS >	~{����|h�ۍ�>��<?��;>��Z��T������~uJ�*Bc?�b?Pπ�h��]P?��x?�ľI<N�va������9��54?��6?�Խ8��>���?��?�.�>RD��H�e����r�x��`Ǿ��>�ѝ>����x�u�F�G=B�\?�8?��>>z�=ܩ���D��u���"?,��?C��?�H�?�N$>��N�y3ҿ7�Ծ����cل?���>�����4?5s=<�՜��W��G˾��Ba����d����'��+S��B�go�=�9?��w?R�y?��]?z�ᾼ.a�p���̠�#P����_S'��wP�]�J�$�D�8 c�KB��H?��n�V�W��n9~�Q�A�6õ?-u'?�]/����>����ﾫ\̾�7A>Pb��������=�����A=3#Z=h��.��#�� ?�Ϲ>��>U�<?C\[���=��2���8�\�����1>���>˒>���>y�/9�.���齱Ⱦ�΃�a�Խ\(v>�yc?��K?z�n?�C�~!1��}���!���/��J����B>�q>���>��W�2���>&��V>���r����v��5�	� �~=��2?}�>��>~N�?�?R}	�O��9Yx��x1��܄<�(�>�i?p/�>�ӆ>�Vн�� ��`�>�Z�?���>���>�}0= �=�2⇿4�>}��>��@>&�-?���>G�����p�����[��F"�|�j>�Hn?)���5�0��-�> �R?qZ�=�XM��i�>;#���+�������+>�D�>`��
��=@���I�?�����&Ĥ�Ux(?v�?Vs��^�-��5{>"$?33�>-^�>��?Q�>7���w�;:?)�^?��H?c�=?>�>���<�`νJoʽ��-��G=���>�U>��q= ��=n^#��zf���h(H=�v�=���!t��x�G<~ؼ��<z�=�'4>�Lؿ��G�ؾ��,}��
�>4��	|�����`�����`��n\�O��W�9�k�T�Pok�`匾W��z�?>e�?_7��j���c����bo�/�p�>)/u�a)� \���齽%���/ݾ�)��}� �J��Th��Gd���(?_���uϿ�u��L���; ?�J1?9�`?���6��7��u,>Š7=p�t��+��S��ۄɿ>�Ⱦp�`?�P�>�������{��>��=2�>�E>w�\�l���L[A�Գ?��?n�>X�j�ʿ�`�����=չ�?a�@�zA?��(���dyU=(��>j�	?��?>�`1��A��밾�]�>q:�?P��?��M=��W���	�%ye?�� <��F���ݻ�=|R�=�1=���i�J>0b�>���ccA�/"ܽ�4>�х>�"�ǚ�,o^����<~]>Ϩս&A���Մ?�|\��f���/�AT���[>D�T?C,�>J@�=�,?:8H�~}Ͽ=�\�-a?�0�?!��?�(?Aۿ�`ݚ> �ܾ|�M?9D6?P��>a&���t����=���<n�����&V���=��>�>c�,���ދO�� �����=o��A\ſN%�w�W��<IT��kb^�m!ݽ[���S]�tʞ�P�j�(����_=sb�=2�Q>�"�>+�S>��Z>
�W?�ej?���>�4>M1ٽ�*���@Ⱦ(U�;�{���u$��1��<g��C�����s�߾���P���H�k�ƾ8��S=��Q��m��lq���S��&,�Q-$?�x�=���%0E�x�=�G��?���v/��KӠ��'ϾG�0�#Y�p��?|�8?����a����h.�=fC�<\@@?.����E��B�>ںJ��=y<о�>.��=�$ѾF/<��4Z�is0?	b?.v��7r��$*>� �n�=E�+?i�?�]<5�>M%?��*���H][>ً3>�Σ>��>�	>���e�۽M�?��T?$��������>�o��-�z�)a=�5>�%5�"�'�[>���<����k�V��"��ij�<Y!W?��>*�)�~��J���@���;=�x?��?�@�>��k?a�B?���<4w��=�S�$ ���w=��W?�2i?M}>}/����Ͼ�a���5?0�e?��N>�Th�9����.��?��/?��n?.V?e���z}��#����[p6?�rp?��W��צ�Oa����3��>��>h?�U.�og�>�k0?5(��D��n�����8�K��?'@�C�?pՁ<ZO-�1�]=��?u�>�Xd�ɾ�����>���E>>�5�>e7���q����$�W���1W?J�?�(?W3������U�=*\���W�?��?4}��qL�<%����l������;�Z�=g���!@�mF�)7��qľ���/���oԼM�>�@�-����>	81�0�⿚�ϿGy��FkվȚt��W?�<�>[�Խ�M��zsh�&�p��C���F���&}�>�>>f���]����t�B	8�y�X�S��>}l~�OË>!�T�;���!��� ��&��>��>Baq>{3ƽ���<�??{���Ͽ�Ѡ�!
��`?Q��?�6{?�?G�+=D�~�I�S�w#K<>?��k?�qU?���οx�����i?����Oe�m�5�|�I���O>W�3?K�>n�-��&=�)>�%�>e�>�/�R�Ŀe��)����?��?����K�>�D�?��.?E���ƙ�E1����"�|�<�3>?�{1>��Ⱦ�#�ʈ:��'��1�?�8?Z Խ�k �vv?B����x�p��򉾶��>!J==��=�eW>�4u�5�v�w��}Ѿ"��?E�@2̱?Z�P���&��N?��>+�ƾ��N�F$8>�[8?,~�>S�>����,�����h_/��C罹��?�4	@_��>����替��S>��w?��>r��?'z->.��>��=�s�0:~<�'=�*�=ԛ=�? �K?���>Uj>U����2�a�A�^N����g�;�c�:>Mk_?��N?v�:>�������M*����_�"���W�XH�̶�=`�%(3>��>l��=��E�ľU� ?�	�RC޿�g�������&?�-�>M� ?a	
�������^�Z? D>���Y��'����r�?Vm�?���>]��-� �u��>��>��>*�/���=�/!��7�=�:?ݾL������`�H̉>�~�?��@lJ�?�j��1	?4������SH}��,
�Wr9�j�>|�8?6�L�c>��>:Ю=^ev�0T��fu�P�>�)�?�?�K�>��g?�j��>�l߂=gם>x]e?��?H#�<A1߾�fE>C?e������;K��ɕj?�m@Pg@7^?6���ؿ:���p��糟���9=���=E�>�L�[���<<
��9�I�<�q�=���>�vS>cA>��0>�*�>�GA>cE��?���0��*-��q(����pC�ϛ����jH�O��Hk�������.�PT�xݾ��|6�G-��)ς��6�=��P?:�O?HDP?t�>�E�<�Z_>?���n�:&��>bH�>j ?��F?$"?�Þ��z��j�Y�p��0������=��>)�j>�'�>#
�>��>'κ��<>�)>Ȇ�>9�5>~�&=%�J���!=�Z>v�>�2�>�n�>��J>�'�=9����9��eol���/��
���?����[C-�b����X�,����  =�?��	>�����Կ�����P?s������RD�'�=�#?Y�J?��>�㞾n��21�=[�\��8��Q�>rK�����5.�9�R>\*?a�f>m
u>��3�88���P� f��c�|>�=6?;'���$9���u���H��/ݾ2pM>翾>_�F��l����� �~�7pi�hz=�f:?vj?8O������@�u����vR>��[>8=��=�aM>�]c���ƽ��G���.=��=C�^>u&?D->�ő=/��>.1����M��ԩ>��?>*^*>q_@?�X%?�K����겂�
�,��$u>�R�>�}�>�)>RhJ���=�-�>��b>�b�i���<��X?�8W>�A��u�]�7�o�߇w=�%����=�=� ���;��](=��?f��@&Z�ܧ��Ҍ��B�V?c/;?$|=�hk�)��j����\�y��?G@�#�?GTξ�n���)?�ƭ?��%��&�>з?��=��4���>��_����3��f{�c��?)��?�;X��\�{j3�`~>��?�5����>B���K�����V�u���"=̰�>�#H?Au����N��>�z
?q"?xY򾃕����ȿ�kv����>0��?��?��m��N��7@��!�>/��?�Y?1�h>?]۾��Y��W�>|�@?�R?��>!��L'�S�?��?w��?��=)�?�-e?���>%&�>�d�\r���F��^V=R0>a��>Ӡ�>~|��ek�P���n��g__�dC�ڝ\>�}=7z�>�N�-#�	.>r�=_0��8������>)�~>�>ǆ�>�g�>���>��a>��Y<-� =�����þ��6?'k�?����/Î�#��<���>#�X���>�-?Y]�>�Aս䐮>p,o?�t?�5?�� >B� �qۜ�%��p�۽��>�к><��>g�<vx�>S���Fվ\�>��q>�}�5j"��W�{��=��@>o��>���>��=k� ?��#?8�j>��>KCE�8����E���>���>NF?:�~?T
?X���[3�j	��衿f�[�p�M>[�x?BY?�ו>㌏�Z�����K�m	H�F������?�zg?KP�W?c)�?ܖ??��A?�Pf>s4���׾񭭽���>D�!?9��R�A��9&� ��iz?�\?>��>N���:dս��ռ����I��%?9\?�"&?L��*a� 	þ�w�<�'��N�s��;UF���>�k>�������=E�>�ɱ=�m�:6���f<�z�=ዒ>��=�6�)��1<,?@nF��փ�dۘ=O�r��uD�t�>aYL>����Я^?�R=�H�{���7x���U����?J��?�l�?�ⴽ��h�i&=?i�?u?��>$O��$x޾Z��Rbw�ϓx�)j�m�>���>�}l�4�Q���S���FG��>�Ž�^�n�>��>�p%?4�>x>O��>���6�;�z�ᾨ$	�@�V�Xr�Q �n	����r���!�_�&�t���ƾH)s��~>�����>z?o�>�a�>sI�>`R:��֠>S��>Z�>�h�>K�6>0L�=��L=�z��Č1��&S?"�ž�F$�8M�� ��%�??�|f?�b�>O�|�_φ����E?f��?��?�-�>�Ue��*��?�e?)D��Q�?�1=�8:���<�ž�)��ƞ���W��>o1�� �2��+U��?��o?e*?^�:хξ�4��Y�����n=�M�?��(?��)���Q�P�o�t�W�S�{��O6h��i���$��p��쏿�^��%����(��u*=܉*?N�?�������!��<&k�K?�lcf>��>�$�>�߾>�uI>K�	�H�1�+^��L'�)����Q�>[{?�w�>�I?�6<?(*O?��K?�8�>��>뱾`�>L�9<ᙢ>#��>
 9?��-?��/?>�?@�*?P�a>���������ؾ}�?��?X�?g�?G�?�47Ľ���=aX�/@w���}=2��<�ֽzv�	4[=�YT>�P? ����8�����uk>�z7?���>���>	-���&����<���>ߴ
?=L�>L����yr��d��=�>Λ�? &��%=�)>���=OɅ�Ϻ*�=������=�F��ߎ:��( </��=z�=*	t�Q���g�:�|�;^*�<W�?�e.?�o>�K>�K��N�ǾW�?� g>��?&�>��>/�ž��z��Ԗ��t��$@�>X�?���?�(�u�ƻ��>��J��㚾��#�!ʾ0ؽ��	?r��>[�1?J��?;�@?� �>��/>�̾Қ�����~��2�?L!,?Ë�>�����ʾ���3�˝?jZ?l<a�q���:)���¾��Խ2�>f[/�b/~����)D�X?�����肙���?ݿ�?A��6��w�߿��C\��*�C?"�>MY�>n�>Z�)��g�u%��0;>���>R?j»>)P?5{?R�X?�S><<5�,ì�����EK��*>r3A?+��?� �?��w?z�>�:>Ka,�M!߾���� �����ӂ�U�l=�Z>>�>�E�>���>-{�={�˽�?��J�:�˅�=Q�^>�b�>lަ>��>f�w>@�<*�C?Ձ�>O���0��:ѽ
#T��J'��o[?j��?�	?F施kJ�"8��X�Vu>�'�?��?$H?(����$�=��^=�Ǿ=;�t�>x��>��>��h>�tT>�(�>T.�>5л>��1��d�)�Y��^�X�2?��T?���<����)�V��|�|�9�&�O;Ö ���U��� =�k�Yh1<��z�Yҍ���e���h�A/����f����Q���b�^�?�>��G>�11=S�Q=�=��=��=]x��{�@=���֋=�v =�G��{�߽�0y�S>�Dr���>=(����:a?�G?e�?V�?��>*�>L6���H=�Y7>a�*?�ѻ>�$���P�wh����)�ƾgfǾ���p�Ԫ���L�=��=��>C�=	�>S>��+>Q��7�>&L�=��>�l��h�=�9>z[�=1�5>�o>�o?��~�-꥿o7@����o(?�r�>W�>U\���~
?y�=�J���Ⱦ�k��ހ?���?RK�?(S�>���	�>vP����=�?=�A��v��>�]i=�됽E�	?�p1>L�/������<��?a@�e?7���/�׿�b�>�Q7>d>R�81�VB\��lb��Y�~�!?�m;�̾n��>�F�=h�޾ 5ƾwZ/=}6>	�_=v���1\�鏙=RK}�U�;=aj=��>UD>m4�=LK�����=�	H= 5�=WP>J܌�!�7���+��[6=��=W�b>�a&>���>�<	?	^)?]��?�~�>����}�������>F]ݽ��,>4����P>�/9>?'?'k?�a?]c�>�֕����>��>��"�c^��[鞾�J���&b=�.�?.$�?��>�k��)���L��2��}��
��>{T?�@#?�z&>�s
��ƨ�i�����(oʽ����Y����F����>M��=��M�i7=F�t>��7>5$>Ww�>�+�>h=�E�>	^�=��<�f=%u��oC��5H=�kF>��c=�ԽX�׽p�.=C�g<���7<-a=�o>��>սY�8=��=���>Ku >��>PC�=��Ͼ��T>�zs�Z�G�`E�=������L��Ao�Je����.T:�	H*>�W:>���?����]?�]>�t>��?�
t?NNZ>C��ڲ�j�N����F�t��=�� >pO9��d@�ł^�gGM�RC���>�ގ>��>J�l>�,�$$?�
�w=��a5���>�~�����42�d7q��>�������i���Һ��D?�F�����=� ~?c�I?!�?���>H����ؾ'60> D����=k�K.q��k���?w'?���>2���D��T̾2/��&ʷ>�WI��O�ؾ���0����޷�%��>s���о�3��a�������B�#ar��>�O?��?b�']���gO�d��
1��\�?�_g?��>PT?v2?�����L�wn��o�=��n?h��?�*�?��
>���=���v�>�6	?��?C��?Q�s?@k>� ��>�Q�;
� >7����=�'>��=0&�= ?6B
?E�
?2����	��t�N���]����<�ʟ=���>���>�q>2W�=��j=���=V�[>���>�N�>R�d>���>w��>��y�U+?"@> @�>Y~.?�u�>C�>V	�5����p=��Ľ��⽣v;,=�+��=�}�]�C�|�:g�>0̿��?�B�=�\�Kg-?�1z-�v�>�s�;�lI=	?��y=M�5>��>�.�>_Cb>9��>'�!>j%Ѿ'�>ܞ��&#�XnC��^P��̾��z>���G`!����wED�𬵾{���3h���{�>����<[�?8�d�k�V*�M
��[?�x�>��4?�&���~���*> ��>1͋>����n������2R����?���?��>V��>��r?p"a?'��=;�о��k��B���H[��܎��;:�'b���u�����լ=��?�?)�?��3��>�
{?N�e�P���>�X��V�u����l>�6�����G�����A�ƾ*>q>�?4PZ?�I?��������u>��E?�?۟O?Ŀ@?5�=?���, ?Ӹ�>�j/?�`7?D?n�?�*?�@�==dP�{W�;����x�ɽ͞��ʿ�3�Z=�;��-�/��=�>xP�=	����1<hB=���<<㉽k3�Lz�=��=���=�K1>u��>�UZ?�k�>�>��B?��$�%x>��ө���:?��==s%�� ���㉜�'�.Ɯ=�u?��?'�d?/0>a�/�J:>���=�,�>�$	>��[>TҢ>s����
�T>�>o�>A��=)$G�kj��Z=�"=~���=�%>M��>h�D>��'�eTQ>B/��𣳾9}�>��X��ս�m���NV���/�.�����>�B?�R?j�=S�Ǿd�<i8{�W_H?n%?��g?sS�?Z ;��h��{���>;�{��<=y�>��+�2�����Ɯ���.��,�<�_�=�����^��A�d>Ĉ
��S�?���(�V�k+��/�>e�� <=&��qоh�l>W��=�ڴ�q��f6�������M?� �=�Գ�&3��m���c�=���>>K�>�v���L+�`��^��=���>]>5�����𾝛C���޾X�>�~C?}�t?���?�m��(�q�փ1��ɾ����Q�u�\�&?_"�>��+?9�z>O7K>?�޾�2��K���'����>��?��.�#A=��pW���پq�5����?�z>}'?��l?�S?�FI?�>c�?���>B�ɽn�q��u ?A��?�	�=΃�h�̼E�J��VE�c҄>�R?����Jh�>�3?�	W?�,<?��:?%�>���>���_,b����>�L�>��`�6���
k�>�,9?B.�>��S?V�?C��>�i6�Ԭ������h>R:_=k�,?tm@?>�3?埠>���>6��!U�=�L�>�c?�1�?|�o?Q��=7�?�v2>���>��=Ѥ�>� �>F?�)O?ҿs?�J?IV�>�?�<e���p���o���O���;�*K<$�z=�'���u�֪��,�<r��; =���|�h��K(F��n�����;�]�>J�s>�
����0>-�ľ�P����@>�p��Q��ي�E�:�
�=|��>�?���>�W#�N��=笼>�G�>����6(?��?M?� ;E�b�t�ھ�K�*�>:B?���=f�l�Ă����u�y�g='�m?t�^?��W��'���b?��]?M�F�<�R^þYgb�<7��%P?��
?��H�v�>��~?| r?���>�g��]n�����`b�n�i�A��=4�>o2��|d��u�>?[7?qM�>{�`>C��=^]۾զw�O��P?8��?9�?�ъ?��*>��n��H�6KԾ򠘿ƒ�?C��>����R�:?���<A�龼�B��x��?վ�瀾E־E��㩈�z�5�2_�� �G�<�C?*.�?Ru_?�v?�2�bj]����������E�u	����yJ���=���S��~��ԡ)����<S���=tp~�>B���?��&?vH/���>�ɗ�����˾Y�@>W���^��,�=vх�&�D=�-Z=��f��a-�e����a ?�>'o�>�=?�\���=��s2��7�����0>x��>�	�>�h�>�C�90��S�[ʾ#^����ӽ�qq>#�V?9�D?؇?�M��8��i��v�����=�����5�=�=�=���>?c��;f���M�y�B��@���"������V��>��:?��=ߦ�=[$�?�6�>Z~,���Q�&+ɾ�J�bA̽��?a�?��>ag�>����h���>��q?;��>��=�ݼ>�LL�������"?}�&?v�b�dc�>*�?�1e����e���Z,�������S�<{��?8�2���+��I�=��1?2��3��=�_o>��>a���]J����$�K�p>�3]?�cI�J,>>OžKW��̾��Z���y�?J�7?�셾��<��e�>Ü�>�-�>5N>ɟ�?�,�>ir^�J�>��1?r�p?%�.?�r?_?�'�=�����-�I�n�1��=�U/>J{>��f>,x>,�+�������0��7�=��=
���|��p&
=�����Ai����=���>��ſ��9�P��_�+�����J��\簽]{P�lоd�A=�s����_�_�I����.#J���X�~�`ؙ�_��q�?}]�?:����|��<���k����+?l��_@������jP� w��\~��l�ľ��<�9XX�#e���'?�e����ǿ݇���)ݾ�]?Z� ?يy?�[�L"�Z�8�J!>ߢ�<0��CO�~����ο���_?��>��y�����>J��>{�[>��r>�c������T��<2�?�-?�O�>�6t��sɿ�`��Xg�<Z��?�@}A?��(�����V=���>�	?5�?>mS1�I�Y����T�>h<�?��?M=L�W���	��e?�~<��F��ݻ��=�;�=�E=�����J>�U�>���3TA��>ܽ=�4>�م>v�"�ƪ���^�;��<]�]>G�ս�:��k�?q�a�RD��^�[���+E�>X?���>��=a�[?�D`���߿	��P3H?Xo@�s�?Z�.?+�վ[Y�>S�辆�b?�
4?xƝ>��)�ĕ{�T)����=
��>JE�Zy�־�=ܪ�>�h>��D�e�=�J�|��<KI�<����/��4������s �m�=N�ּP�D�ԊD��\;=|���tp�xd��ϸZ=ܘ�=$q_>�.�>T,E>�z>��^?�n?ǧ�>Q^?=t1�*e�9��v՝�e6U���4�홙�M���Į�)U㾱�վ���@��I���ξ+�:�Q	~=eaQ�#���G;+�q�_��u8���+?�	>���zP�>��<ǥþ�:��κ�R�����˾h�0��"g���?�IB?���f�K����mǽ�Ͻ�>b?�*��!��$��p��=����Z=�>u��=h�ھ�Z2���T�G0?ȹ?G���S����,>����%=�+?�?5�q<���>6^%?(�Nܽ,�[>x�2>���>���>�>u宾�ݽ:o?�<T?r������Y�>F����}�N�\=�>��4�������[>#��<�Ҍ�l�a�*�<��V?�j�><V)�YE�6����>(��:,=fOx?\�?B��>0�j?�B?|"�<N���RT�rU��+k=b3X?r{i?��>�#Fо2�����5?��d?��M>u�e�?x��6.�Og���?��n?��?�'���h}��=��6��$6?�?Q�t����E��N��Er�>¤�>%�>��E����>��?�.����>:��!W=��k�?A�@H�?��U��N���HW���?�q�>/o�4���3�#&¾�?3��	?����i܋��);��W��U?ʛ�?{�>�^��$��`>󿜾Uǲ?�i�?� ���/o=�o�28w�J��,'�� H�=�e�cm齃�ݾ�8��̾�_��g^��(2��@�>��@ddL����>��9����p׿ց�V�;ȫ���S?�pE>td�پ2�{��k�J�3��+�f�F�>K�>�>)�������N�{��p;�%���#�>�(��
�>��S�g%��왟���5<��>ȭ�>��>|2���潾ř?/`��:?ο����Z��6�X?�g�?o�?�p?$9<_�v�{�T~�v-G?)�s?.Z?Ux%�*?]�"�7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�_�|=�>���>g>�#/�y�Ŀ�ٶ�@���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�b�_?0�a�J�p���-���ƽ�ۡ>��0�f\�O������Xe���Ay����?Q^�?o�?���� #�d6%?�>L����8Ǿ1�<���>�(�>�)N>�G_���u>����:��h	>���?�~�?^j?���������U>�}?�N�>K��?_��=N;�>�==߲���4�rP'>�=e�L��3?�L?�]�>��=*$6�1�/�"hF���R�ҡ	�?C�H��>�b?{K?��`>�f��!3�����N׽��-�#�bZ@���?�l�ؽ�9>�=>�>��C���Ӿ�90?�$���ݿ����&?��;?h�>��>)�9
��� h���^?Ƥ�>k��7�������k��?��?E�?'{��/�N�6>��?,��>�u7��ѽ��i���S>��5?1�ս����ӂ��2v>�S�?�@7^�?&~}�q~?�� ��n���|5��%*>�*,?f����>'h�>:G>Q�o�x���r)x�+ź>Ea�?��?G#�>۹e?�?s�� 1�Yk=���>�Jh?���>͛;����=>�c?N�'�����f�_?ӌ@�@#�T?�]�տ�����殾[��x��n1=��->����[��=�V�;�]�>�Ir=͡(>�E�>�H>�:'>�02>і@>|��=@��T��Y���i���m���Q{ �i�
��޾wTe��r�:���`E��-����Aڽ�Mo�_6_��/�bG�_`�=�yK?vd?
�?�G�>���t�=*��#��hfZ���k;M>��4?�>?1V&?w�������wi��5��*���f�|�(4�>W[%>&��>��>6�>54���=t�>��>� >[V�<^�z<l�=��h>Y<�>~�>﷗>�{;>3�>D�������Ri��_y��ɽ �?<'��OtJ�\vI��R<��
?�=<�-?��>�푿'пAĭ��aH?�����k��*�R�>/g0?�QW?��>7��BgR�u>�~�kh�}!>�*���m���)�"0P>��?nmI>~am>H�1��:��1^�Yd¾D��>��8?m����2�6~p��S?��fӾ�A>��>1��
�����x���F��޻=�I3?��?սʾS�����f�A�B>Q�>0!�=�-=�`O>`�����M�T���=b�=�8>]J?`,>ُ�=ܣ>\I��sP�瘩>��B>�,>a
@?�$%?�q��&��+����-�]$w>G�>?��>�8>mjJ��}�=�_�>��a>�����������?��:W>g�~�~�^���t�u�x=iK��+��=�8�=�� ���<�l
&=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�G�>�R�� ��'���!�y�_gV��s�>�6<?Ⱦ	��n�;������
?2?.�ƾGR��y�����x����>o��?ə?Qv����-)��H?tn�?�1R?ȕ�=9dϾ[Ƚ�>^CH?��H?��;>� �˚5��T?H;�?\�?�}N>�?&
q?IU�>���7�0������~��[�=ya�/�>2w�=�Kƾ!(G�_�����&k��~�]kz>�0=1�>�����K�����=R3������	*�R��>��z>ɝ5>���>v
?f��>�/�><�n<X�ս�9���A����K?���?����n�7��<�2�=� `���?�5?�\$��ξ2��>�]?�ʀ?�XZ?�>���r���S࿿6��H�<{�I>)��>��>q�����M>f8Ӿ�@����>���>"ȴ���ھV���&����>�>!?��>% �=ʱ ?m@%?]jj>���>̦8�������L��/�>W�>��?)Bw?��?�����9�%���ܞ��9�a��I>�!}?�?t�>�֌��w���Å���ʼl��]��?ovf?�b޽��?S�?��C?MC8?��b>�� L׾4��sց>ߞ!?���&�A��!&�����?(o?d��>U���:}ս)�ּ�������?J\?�@&?^��@%a�� þ7Y�<�A+�9�f�O��;9H;��X>�>�̈���=��>�ٳ=�pl��B6���_<�=���>s��=��6�.'��6,?�;D�dł�Ⱦ�=s���C�m�>��H>�x��޸]?|�?�#a|�a������N����?pK�?Iɕ?�����i�}
>?���?L
?<��>�����cݾr%⾤}�חy����j�>��>�}��{��R���^/��@ƃ���ʽ��L�+?�e�>z?F��>kl�>�?������04�����Դ���5��K��a�q��ZZ���G�����cԾL����:>������>e?u��>qTE>��R>���MV?*\�>d�;>ϫg>o�>�	G>%��=���<R낽�KR?����#�'����²��e3B?�qd?Q1�>mi�:��������?���?Ss�?=v>h��,+�n?�>�>F��Vq
?�T:=p8��:�<V��x�� 3��1�*��>�D׽� :��M�=nf�uj
?�/?����̾�;׽}n����n=7W�?l )?M�)���Q���o�K�W� S�a���h�倡�T�$�Q�p��쏿,Y����s(�GU*=�*?l,�?ʩ�!��>k�H<?��kf>.��>��>E۾>��H>�	���1�^��='�����>b�>�d{?�-�>��G?!:2?��@?��\?&;�>kj�>m7����?k�=��?{� ?�x.?R�W?7g0?5��>�?ѽ�>��Ľ
 �(z�O?�
@?���>)��>�9�>-�Z��Z�.�&���#>B�X�p::�3=ⓧ=C���/��a�<��>�X?X����8�3����k>��7?T�>���>���`+����<i�>��
?J�>J  �V}r��a��V�>ꡂ?� �{=n�)>���=+�����Ѻ�[�= �����=LB���m;�Z<�}�=���=��s�f�����:F��;���<�}�>ˎ$?���>��0>�	�!#�E'4�f�6=&ʙ>��w��>��2�������y�<�>��x?x��?�a>���=��5>��۾�������S���LS�v<?`#?��e?6)m?ʩK?+�-?J�=Vj�Qw���Ӓ� %����#?s!,?��>�����ʾ��׉3�ڝ?k[?�<a����;)�ِ¾��Խȱ>�[/�f/~����>D��텻���A��3��?쿝?wA�Y�6��x�տ���[��t�C?"�>Y�>��>P�)�|�g�r%��1;>���>fR?�1�>NP? {?DY[?�9U>�8���Ϭ����tT">[@?<��?��?py?�d�>��>��(�@�p������w���LT=23Z>޽�>�5�>��>��=X�ƽY.���.?��W�=�Tb>4H�>M��>��>,%x>|[�<��G?���>�]����=社�Ń�e=���u?M��?ӑ+?R[=Ԁ���E��B��xJ�>Gn�?f��??2*?��S����=��ּⶾ��q��%�>_ܹ>43�>%ʓ=5�F=�a>��>���>�-�H`��p8�LM���?�F?��=ȬĿ��o�o�u��x��/�Q�&����T��1����u�[/�=�����Ţ�q�T��������稱�Fě��5m���?�^�=��=�=(0�;��ܼ]��<p�h=���<�]�<4t��oa�;�H�0� ��V��6�!�m:��=u���þ��v?�O?��7?��=?��K>�]>��;�i�>�"��`�?&�/>���勳�/g��9��Et�����{��^������>4d�.:>�>>r��=9<��=�=B��=il<�Q=���=y��=zQ�=UG�=�`	>�g�=���?JC��㽜��D/��I%�f�\?sO�>�En��X� �r?M�U�������L��N}?Lp@�z�?�?5oB�{>yqS���
>$[=�秾3~�=~�1>�,"���>��>}�	�\�����ǽ?^k@��3?�˗�d�߿f>�.>G�	>�Q��z.��]^��nZ���F�V."?�U:���Ⱦ��>y��=W%�*ʾi;=��;>�VU=�"��Z�H��=����,O(=��v=p��>�G>�F�=�Ȱ�2'�=��=�M>��U>]$� $8���<�|;=�=��^>�1%>��>��?=^0?�Nd?A=�>�"n��%Ͼ{A���\�>��={F�>�=�B>B��>��7?��D?a�K?���>�~�=?�>��>]�,��m��R�Qǧ�X|�<�?�Ά?�ظ>�9Q<��A�6���c>��BŽt?�Q1?�n?��>�7���vK,�G�!��|�����= �}=���(K���^>��x>�x��=>���>���>�<�>\6	>�N>aS�>k��>jO1=(��=�H>S�=E��=�=�4��ə�R��>�W����a��d��3N�cX8�h4�=m�E=��	<b6�=FG�=|,�>�'#>�j�>Zv<�Z����f>�g��Q�:�X�=��ؾn�]�,{f��[|�."���½;`a>��>͠�=o��h�?Ï>��>���?�Oj?�*s>������㋿<�r���|��>"�9=krp�}�A�Ȉd���L�Ծ���>��>6�>��l>�,��?�[/w=���W5�'��>�r���`����<q��@��
���Ci�8�⺃�D?^E��ȉ�=�~?��I?�ڏ?��>����+�ؾl#0>J���=7�Qq�^!��U�?='?��>*���D�|H̾B���޷>AI�D�O���+�0�$��Bͷ���>�����о`$3��g������ӍB��Lr�D��>�O?��?�9b��W��4UO�����*���q?}g?G�>�J?�@?!&���y�r���u�=��n?���?1=�?5>^�=���v��>�%	?r��?�?��s?*?����>k�;��!>������=��	>+��=K�=B5?�(
?�m
?�p��s
���j��f]�Ͽ�<�ϡ=2��>a��>i�p>�F�=oNn=�g�=w�\>�y�>�ŏ>5e>bA�>�5�>�䵾�|!���+?XC*=���>�TI?R��>Y����+���νw�>`�K�����c<�rO�<� >ı�=!?,=C�ý��>-�ѿ*-�?[1ؼU���>���z����>qv�=�F~��d?� >�?��>7H�=�8G>�T�>�?�=���e>�`��e �>rZ��{]�:��d٭>�Iþ {��	������#vj��|���_�&f��uI��(?=���?b +�6?��3o�7��;<?L��>�$?Ė��W�$=�Y1�0�?SY�>?������)��.ﾖ-�?���?Qt>|��>�fk?i�?RH8��ZG�9e�N���%� ����D��I��.C���'�0�h�q�:?7ko?��X?�!F=:�i>!��?��H��K���,�>s�M��X�!'>rݼ>+���5���Mٰ��� c�=KsY?$�v?�7?v��Rak���>g�0?�?(�|?�X6?)�+?w��G�?�V>ӏ?h?�(-?-T?U_?c�>oC#>#�~=��!=��ҽ����sj<��>")9��M ���=A�O=rZ������'>jl��b��y둼��=l�&=`+ɼ-W�=��E>V�>�$^?��>"�>�!8?�j��7�l����n0?k�C=�b��4��]ԟ��ﾭF>`j?\�?�Y?�M_>��A�BD�m.>+�>	�%>l�^>\�>1�𽨖G�(g�=|?>��>83�=xvI�[���	�}����C�<(� >=�?C�V>�zK��1b>%(ؾ�{���>.�U��s��+��p?���H���þ&'�>YX?d�.?)~B>��ž�$��M���1@?�\4?�1?�X�?zS=A�̾I�E�T���l��h> l�=�C��ns������S�K���U��FW>Y���&���aE>U�.d � �d�/�F��С��о��U���=��#��!̾�~2�7o�=��=���bm�Ğ��Q����Y??�>���8y�{��=��>#r�>����r���T�����
�P=x>�>8".>!"� ��@�!���`�b>�:?�/]?O�?�q$�������J��.��y��LT���>EM�>��%?X�n>�y:>:���]9�;c��yn���>d�>Rv�)F�$��O���j/�	�>j�0?�3C>���>�O_?c*?MVR?x?{�?�z�>�C#�甡�I�?rބ?�]M>o\g�f���>���F�L[
?p�j?gy+��Ў>��%?��H?�v@?�h-?R�?Ga>�оÉ_�<x>#M�>N6B�{�Ŀ�%9>�f?m5?g�n?��p?��$?w1�j�;,J���>;N�=�?�EM?8K?,�>ً�>C��yK�=qg�>,�b?d8�?��o?18�=��?��2>=N�>_͖=[��>� �>?�O?�s?N�J?ځ�>�Ō<����J��$�n�LR�6�b;|�F<� |=���y�u��F�Q��<;��;~����
��g����D����AU�;/;�>+@t>�n���O1>J�ľoꈾ#-A>�ͣ��ԛ�ʒ��!�8��W�=���>B?bƕ>h\#��	�=�Ѽ>�>�>j����'?��?�M?^&;��b�u۾�K��>��A?�7�=�ol��O��q+v�.�e=�m?�w^?��W�*�����b?�]?�g�|=�=�þ�b����O?��
?��G�G�>��~?��q?X��>��e�s:n�5��Db�S�j��϶=�q�>'X�C�d��@�>��7?bN�>k�b>�)�=�v۾��w�r���?5�?��?���?�+*>��n�*4�R���ϒ�q�i?�"�>tP��2?K�M<Bξ�Os�����ʾᙾ�]��1���F���%>��|b�K��[n�<��?�D|?��|?�a?�p����o�?R���o���uK�8�y--���4���/��BR�,�u�ݑ�S^��:����<�=��~��B�:h�?��'?�p0�a��>���ܗ�*�˾&�B>�������@�=����VH=]U=9�e��.���+A ?kz�>���>[�<?6�[��2>�SB3�8v8�����f(0>	;�>�(�>�V�>r��{0�ܱ𽜰ɾ�焾1ӽ0+>�;S?d�-?��?陛>�M�χ�&6�A�A>[�.���>���>��?�����5��7<���M�r	p�����u�������R>T1?��x=�p�=�?H��>/�5��K��8t��6���2��q?�Mq?</?�A>�,���5��9�>�t?a<�>i�i>FZ'���抿BvE����>�Xl>�L�>��>�Ľ�S�*�� ��>XS�D)=wŁ?��h�F�_�e!>ԂC?�h�<DS��P)�>E�p�#����C�!�AyV>�=(?@�O:\��=����a������j���T?D&0?v&��Hq���g>á>?m��>:_�=�ٖ?�Y?��9���~��/?T��?$�,?�>e�>'�>&z<�_q�kI���= $�>�d�=��>�?�>��龱��`���>	L�<�����=Ȍ>�%�!kC�%j&<v��>=�п��I����;	�탾��3�L�v�K�縯�1���о����5�*q�}L��3�j+Z�2����c��Z�?���?�3�~D���m����p�_���8��>�jG�G�:���Ǿ�;���W���Y����|�÷P�-v�=�z��K"?����jȿ�읿�����?�&?e��?R��>���RH��FX>Z��<ی��[�)�����ȿ�����X?OD�>����-ɽ�1�>�+�>ň>��f>m?2�)>��z�3=`�?�\<?��>𻟾�tƿ����ƚ=���?��@ }A?��(�c���V=��>#�	?��?>�S1�rI������T�>c<�?���?�~M=d�W�<�	��e?2�<��F�V�ݻN�=<�=H=^��B�J>\U�>���SA� @ܽ&�4>]څ>�}"�ͫ���^����<��]>)�ս;��H�?�av�
�p�k>%��R���=6�U?�>�<���> )c�r�ֿ��y��?�@3��?%*?z����>T�ݾ�Q?�A^?T�>��H�۵���>J�a>�=�y)�s!q�A�d=�l
?R�=�ࢾa��HM7��h��2�>)l���ƿI��-d���=��F��.���k�G�G�o�����S�t4���A�=��=�U>-��>��3>_k�>"�g?ƛv?���>:�>����
 ���m��}��׊�+���j_�������4��z,ᾇM��.����OWվ��;��!�=��R��q���4 ��Ab���B��*?g>@�ž��N���<�3ƾ-M��WG��飽��̾��3�`>n��<�?_�B? �����V����F���1��uW?� ����~&�����=��J�=���>�ĝ=)w㾧-3�S�[a0?d?���*\����)>�d ���=�+?�?ˁa<�z�>e9%?�X*�J�ώ�[>ee3>��>���>�%	>�	���ܽ'�?�T?��� ��;��>Y����z�o!_=c2> �4��@���Z>��<�Ȍ�j�U�"c��7u�<i'W?���>b�)����\��w��"9==��x?#�?�.�>�yk?�B?;Ӥ<�d��h�S�G ��Uw=��W?\*i?��>D����
о肧���5?��e?�N>`ih�z���.��S�U$?h�n?x_?Y����v}�������o6?n��?9Wr������Ͼ���<�>�'�>B?��:��^�>NF?�hʽf��� ��haE�ƣ�?A�
@���?`�̽�z<�����>r�>���m����J�8��;�t=�`�>zU���x����%��:9�ܼR?R��?���>h����d����=a������?��?���Q��=���jo�;��d���X]=4,��xý�����2�˕־����PΑ�JXH���>��@J��V��>_ɽ�s޿�eܿ�ق����Qv���u�>َ>�=��{!۾s��Aj�HrE��i%�i��@K�>��>�֔�������{��q;�(���"�>�1�=�>��S�M%������H�5<��>��>Ѳ�>�\��0�Eř?�Y���?οߩ������X?�g�?bo�?�n?K�9<l�v�.�{����,G?�s?�Z?��%�K>]�R�7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*�{�+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�n�_?E�a�`�p���-�$�ƽ�ۡ>��0��e\�(P��$���Xe����Ay����?^^�?�?e��� #�o6%?��>9����8Ǿ�<D��>F(�>�*N>uH_��u>���:��h	>���?�~�?_j?ݕ������oU>�}?9��>)�?bI�=�l�>��=�ϱ����O�!>_�>��X�٫?�6N?��>yv�=�*?���/��F��PR�����/C�^r�>��`?FM?�\g>����ޕ*��i!��(Ƚ��6�pa�NhC�v���6׽�t3>�@>��>\lB��վ%�"?���K<ٿa0���[o��-?�;�>�D?x�$�8�μ�Jl?�ga>M�3$��t,��K��.�?�Z�?�?R���dQ��f�/>���>/�>���w�j�X���0�L>��R?W���X���p��?>��?�	@��?,�[�!�?[+��|���'i���ĳ�U�4>#[Z?���˼>6^�>7�M>�u�s������7K�>I)�?��? �>��j?f����4���>���>gas?�Z�>>�w��"޾�4>�e�>�b"�;���� �E?��@�5@Ga[?7u��w�⿪`���ԣ�@6羂2+�6Y���	 >ׇѼ�!�<]U�;��=0�(�L>��>U�>��P>��>�a>~c.>&Y���}��C��х���c�p=��n�`-C�k��������Ad�����O�J��f���L��A_��2ʽ�����=q�T?n*R?4dq?�?�ϑ��>�����A=91�t��=���>\x2?(�K?*?��=l����e����줾p��L��>09G>f4�>��>N�>Oqq;�1N>�C<>�|>5]>G�,=B\K;��'=>]U>��>n�>T�>�p<>�R>�p���鯿H�l�a�����~��ם?	֤�c?�Ue���凾$ά�`H�=C�(?M
�=1J��ՍѿEW���IF?�0������7�la�=)�)?�T?�k>�*����,���=�&��X-����=�
�qc��A�&�c�j>L?aIf>|�t>�4�dr8�^Q�����!>��5?ɻ���{7��@v�f^H���ܾzaL>�;�>JC�i��)����.�g�I�~=p9?�U?mù��P��ϝs�5��(�P>��[>��=�6�=Z�J>,)f��{ǽ6JI�Y�*=��=2�`>?}1>��=VZ�>A�����E���>��>>W�2>#�>?�B)?6P������xo��:%���q>_��>I��>�:>�J�>ę=7��>��q>mN��什����k6�58W>�Ӕ��_��<�im�=V�Ľ���=�	�=����<�,�=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ?��>������7����~�<g�>�rU?������:�c���?��>����ۇ��b�ſ!5n����>O��?ĥ�?��l�!{��Z3��?�#�?D�K?��w>J�ԾZ�5�[�>S�A?�0?/y�>M� ��:�4)'?ų�?�.�?0�O>���?��E?��j>6~�>r+��!P���#f��/>�߼z�1>п�>�:\�2B6��ؙ�������|�[˾z�*?���<�l�>y]������J3M>_s�n���H=o9?�/�=�H�=��>X??�j?>7>N���G'�����sF�V�K?޳�?3���9n����<"��=��^��/?�T4?Q�X���Ͼ�Ш>��\?�À?��Z?�d�>���5��d翿�|���Ė<s�K>��>�G�>����qK>P�Ծ$4D�f��>e��>�����Gھ���a��p7�>4b!?���>߮=�� ?��#?C�j>�G�>7"E�����F��g�>�q�>�'?��~?��?�幾wW3����ޡ��{[���N>Ey?>?;�>A�������s�8�ŒH���o��?fsg?����?��?�v??!�A?X�e>@���ؾL-��72�>�!?&��_�A�A&�j��|?�a?���>����6�ս�Լ]��K���#�?�\?t:&?��'a��þ���<��"�[�U�, <#�A���>ܛ>h���e&�=Q�>�d�=�m��!6�+h<4��=ё�>�
�= 7��!��W�0?C���Ҿr��q�=X��/�W�x˝>�x�>�z��Pl?�ʺ�O���+������T�½{�?�?b��?��$��Dt���O?�?��?s� ?�c��y7�ty��ێ���ߜ�:���>&��>������և��ȓ������"m�UxY�T��>�φ>��?�(�>�]>]F?�]X��������|��C���G��$�"�/׏��Q��1/������-�i>��;}Q�>��?Ir>��(>��>��Ľ1%�>A��>��>D��>:�>ũb>�[>\��= m0��KR?���� �'���辰���y3B?�qd?�0�>�i�!������s�?���?`s�?K=v> h��,+��n?�>�>B��Aq
?�T:=#1�e:�<�U��H��%3��Z���>�C׽� :��M�,nf�sj
?�/?����̾I;׽0#����=��?)9?#��s6<��;t�Be[�ږM�1ܽ�lv�D5��f&�c�n���������y��t��=�!?;�?_i��b��K ]��^�YrU��b>���>�>ʘ�>e>���� �(��CY��_�\z��l�?��?-�s>287?��Z?W�\?#)"?�q�>��>������?���;��?���>{�=?�eE?%�!?"��> >?T��>[O��������8?!N:?�??0��>���>X�	�p�%��NC������@˽�D =;�����i.���_=70�<�'>V?�x��8����?
k>?�7?�m�>���>��`#��T��<��>��
?�F�>� �or�_f��K�>L��? ��y=�)>��=Vo���OغVM�=<����=�낼^;� <���=�Ĕ=�Cs�E#���=�:�+�;rE�<��>TE?bҋ>��>��������N�=�sW>p�Q>�>�ؾ�L��Aї�)�g�1u>�ʏ?5w�?�{=�M�=�L�=8��o¾-�t���(��<�?g�#?��T?�:�?�<?�#?G�> ��C��4���MB?s!,?��>�����ʾ��Չ3�ޝ?k[?�<a�����;)�А¾��Խݱ>�[/�b/~����=D�����X��/��?뿝?�A�R�6��x�ο���[��t�C?"�>0Y�>}�>\�)�}�g�t%��1;>
��>qR?�4�>��O?{?$c\?��V>�\9��̭�硙�H'���>H�??se�?�͎?�?x?�>�@>��.�-⾍���8��~�𽥢��	Q=ϳW>�Ց>_�>�g�>^��=y�ƽ�����;�ٝ�=�&e>ы�>(��>��>��t>O��<_�G?��>������A��������4=���u?��?ȧ+?ً=�k���E������/�>�^�?R��?�9*?�TT��l�=�ּ趾Bor�W*�>�:�>���>gc�=�F=�F>���>��>����:�Z8�|�M��?F$F?ֻ=�1ʿR�s�r�t����D�� ��$
d���y���_�#�=�ˊ�Ҵ�Aq����U�Vz��7⓾�n���֒��w�4��>���=4��=Bӝ=tǥ<(���j�<D9=�9�<^�
=e��ñ<��R�d��;X1����]�|'<��=�K~�P�˾@3}?@�H?m+?�TC?g�y>��>G�.���>r���Z?R�Q>c�^�Q���_:��ާ�O'��O�ؾ�ؾZ!d����k>�SE�x�>�P4>!��=+?�<��=�#n=��=�Ҷ�� =�c�=�ݽ=�q�=5��=��>nM>=��?:��ݥ�S|8�ߐ��\]?�`>���=���Q?� ">}M��HV�����Ie�?g��?&��?�p?����@ho>`Ҍ��;\���=P���1<��(>֖\����>H�=�{��Z(��t#�U��?1�@��[?�����̿j�>��>ǲ>M��-&���N�*}D�Bg��� ?��G��Ⱦ�"�>G6<���4gؾ�@L=��;>�7*=D+�m�\�z@f=k�����&=�!�=��>��[>20�=�Vƽ��k=t��<�'>��f>{{�<s[��R�	��l�=�/�=w>a�:>�s�>�?�q0?�Rd?|:�>bIm��_Ͼ�I��Q)�>s��=c<�>��=��A>(f�>V�7? cD?�K??ֲ>�J�=�ߺ>z<�>��,�Y�m���來���&"�<���?�?���>oU<[�A��q�K*>���ŽS?5#1?,�?O.�>�4�&�߿M����*�.�y����=�	���kJ��c��v����c_�=?�>n#�>��>���>*u4>�fW>@��>gv�=cE�� �=8s>ߟ�=ԩN���`<.�8=��>t�	����=��]����h��C�=��3<|�B����=Py�=���>	M�=�"�>)���]�оx�>=讽'�^�)�h>Z��ٴf���r�{�����&��$T>��=��'�����?>ޕ=R>�g�?]́?ȍ><����
��
��'��=��a���	�=N~��s[�3Vf�z�A���	����>
�><�>3�l>�,�#?�t�w=}�]5��	�>�|��.�����:q�L@�����_i�g�ֺ�D?�E��Z��=f~?;�I?��?ֈ�>���0�ؾ@0>�M����=��Eq�t]����?'?���> ��D��D̾g��@ܷ>{<I�M�O����Y�0�i��ͷ�l��>-���:�о�#3�Eg������C�B�Mr����>D�O?��?�4b��W��BUO�9������n?�{g?��>�K?^B?#��q{�mr���g�=��n?ٲ�?�=�?�>_%�=�ϳ��,�>X	?)��?C��?�~s?Et?�m	�>�;I�!>?�����=�#>Q=�=���=R?Ò
?��
?̓����	�i~�sm��]��v�<���=���>���>�1r>���=z�j=�4�=�I\>﫞>�я>��d>���>gR�>�h��T�-�?A�b>�ٔ>��V?��>��>�;W��f��|>�^�?����짽Eϖ;��0=���=+�=^2�s��>��˿*l�?>e7>7j�[�-?u��ˆ���?��j>� c�"�?@��>���>��>��=i>�[C>��=����h>�"�QC'��&Z�V��Y��॔>0�����f,��%���&��\������϶\���~���L��c��[��?��dd�A���J��@?��>{Y?�.���#�!�$>:?�1>��	�^ᑿʿ���̾��?M��?��b>�Ġ>3X?K�?��,��\.�0w[�Squ�̒@�ޢd�d�_�R㌿Q������˽|�\?��v?f�A?IY�<My>bJ�?z!'�����#��>b�-���<�C=�>��]�^XԾ�'¾E���8A>]`m?�т?�?�NH����#�x>��[?z&,?�\F?|<?��1?Wl5�7�?Ȫ?>q1C?�z�>x�5?�3k?��?
��=�@�=��!>���=�ﺽ����ZW=��,>C����Z�Qk=B�&>�+��U�Ͻ��=n�<k���ͼ�	���!�= �)=��0=٥=࿦>5�]?���>KF�>[m7?���+�7� ����R0?~�P=�����"��9.y>��i?���?<�Z?)�_>��A���B���>��>��%>h!`>y�>����qF���=FS>�w>)t�=��<��π��
�ݬ����<�">���>?w>ӊ���'>��nх���k>��.����31�~�L�q5��d��N,�>6�I?��?qL�=��1q����i��,? �7?�I?톂?�y�=��׾J�;�B:O��N"����>j}<���4'��7���b�B��xc���_>N���9+�=,�M���+��3S��1%�'L`��٧��,�3��>7�5�b'}��,޽g�!�˕>�~���#��f��9(����`?,[<<��ľ��	���	?�=>{�>n~{>�����f�/�4�����bk�<�G�>��H=PN������M�څ��v>�~I?Gnt?m4�?�Ya�F�t��b2����������E#�4?���>�k ?���>$�>�Aʾ0;�~V�(e�2��>(�>�*4�o|L�)���KϾ�6#���>�N?�O�>���>�]?��>�4?Wf?�?dظ>��)��G��a�?���?)�=>3�Խ��&�:�$��C@����>��9?
ɽ��>��$?Fn8?)Y;?�D?���>��c>�9ľ� J�d�>#�>�Nk����G\>MTY?M��>4�F?�{�?�ȩ>���oؾg��)��=�Y�=۽%?�??�>?�c�>��>=����=���>��b?S��?�o?{�=�?�%1>���>��=O��>���>+�?I N?�xs?E�K?���>b�<P?������`�v�<�X�r;Y�t<v=�W�L{�n��a��<�a�;GH���u����E�G�����9�<���>Q�u>���]5&>�lݾ}ᔾ<�R>�n=���?��SE��6�=ng>�q�>J��>Х:��]M=�T�>]�>a��h.?�???6O):�j��B��g�\^�>>�<?Q90>�p�֗��q~�q>=�8l?�i?���w��za?�a`?����l>�績��f��L����K?v?ͣ=��+�> V�?;�t?���>��{�:,o�Uԛ�s�c�Hf�VƯ=AϘ>K��9�_�eӚ>��4?뇼>pY>xD�=H�ؾg�u������?�J�?�ȯ?XO�?�/:>�n�/����澐���01e?'|�>�}u��5?0��<����&_���~��lA��'���{�ʾf~u��ʎ�1}��4m���э=[�?[x?wFx?�Y?��_Wj��4r�9E���BP��.�K�-�-�{8��B�rh|����S�IV��;"�=�t{��iC�^9�?��%?� �8B�>�����7��S̾�P7>�o��^����v=�x���X=�\=�Gc�S5� �W ?��>�K�>��;?��W�2�>��5�f=;��p���~">4G�>.W�>4�>�8"�Q5>�57�)�ƾL���̽�:[>K0s?�qQ?1�X?�Q>�N�\2���o����=�Ό�=�X�>��?
	;�r�Y�@�J�ޜ0�����4�E������h
��S�>�O?Ŗ�=��>��?���>��R�����Z����=�ʌ���I�>�x?�W�>o,=�
����$��>i�n?� �>6(�>����� �[#�S��D�>	��>$��>f��>h(�$BZ�)������<�Ƀ�=��k?T���J�Y��>\^M?�n���<�J�>����- ����U&��W
>bt?��=�)9>�ľ�����{�C}���9?��'?�x���:��d>�~*?i��>��>�u�?�2�>h�u����<�?� �?]*0?r?� ?G;�>�L�օ�Y �匸=�r>#QP>��=�.r>�D�{Um�}�Q��ɡ=%��<���+Ԝ=��0�ݳ��\�y}q=\K�>�ϿKmG��6��)8���־��	�J�x�P���ro=겾�����.5�����\$��6�6Ђ�������O�?�Y�?��tX׾����?yq�=I��Mq>�D׽��>j�Ⱦ�-ż(�A����R����k��>�ӡo�\,-��{0?37����˿�	��n��4?�`5?I"I?׸�-���FR���Q>��=��
��h�T����!˿f��ċ^?�w�>ۗ��u�;3��>4t=4�2>P�Y>&�L�sI�өB��?Pj'?F�>P%���ſ[��Y"�<�l�?�	@�|A?��(���쾆�U=��>!�	?_�?>�Y1��H����[Q�><�?���?"~M=�W�Z�	�*~e?�<1�F�Y�ݻ7�=�;�=IQ=�����J>V�>�.PA�(DܽW�4>�؅>ax"����^��e�<e�]>��ս%7��4�?
^�c�Y���ޒ�����=��??b�>���=w?߅Y��}�"}��?:#@5�?T�?У����>��ݾ��;?�\?��>ilx�1����$=�Ɛ>��]�g)˾]�X�o�'=DkY>Fݢ>7�G��a/��0%�C�=��-��F �J�ÿ� �^b��o<o�U�P�߼M��Q�o&������q��fݽI�V=���=gHM>j�u>ȩS>��I>��Z?��k?�^�>cA�=�������ަϾx
�	�T�Vۢ�Z���n���̞��?��^�Ǿ�K���.��ٰ�u;�Z�v=�T�������_��A�4"'?v5>O��'&N��<����-s���!V�����u�̾�82��Ze���?XA@?�ꇿ�[Y���&�˼+���+hO?����"��Г���9>�aw�bs�<	��>��=�]ݾ�2��6O�A@0?�?�<���I��m*>?����x=t+?]?��n<�P�>&%?�v(��S۽m[>��2>���>�'�>��>�ா�D۽�O?��S?9*��웾V��>�n���|z�9�\=!�>l�5�֭�,8]>�'�<\����c�����j�<4'W?.��>n�)�)�3V��*;�w�<=��x?��?w#�>wk?�B?�<-k��`�S�d!���v=��W?R/i?�>x��	о3���6�5?��e?�N>Zh������.�GT�)?}�n?{a?�Ý�\t}�������[n6?�|?�;Z������⾐�����>a��>!!�>E�,�؛�>}�?"F�_A��ν��U1�C��?��@��?b��<h�a<�,���?%�>=��	�[��D��B�ݾ�<6��>�>s����@u��+��P����B?-�?�>�r��yv��h�=Uޜ��e�?x�?Bm���=�gf�{5�n��1�.>����1f�]վ�1��
ξ��� [��צ��N�>$e@L[����>�%=��� ~�`�����Ǔ����>�^�>"�_��,��t����΂�.
O��"��t����>�D>Uz������=�{��N;�Va��j�>B�	���>�pT��յ��9��-<UԒ>`�>�U�>�߰��D��Vϙ?K����Dο����V��4�X?�B�?�(�?�??'
C<e?w��<z�����F?J_s?u�Y?��$�w�]� 7�ch?�8��OUm��2�']��r>�-:?-8�>ʖ"�Kk=�MP=���>�$>X#��ʾ�mޱ�51���?�u�?������?�՘?MqC?�<��=��ӛپ���h��=�*?���>pX׾ �2�
I�]䡾�&�>��C?�C�=c���`�_?,�a�N�p���-���ƽ�ۡ>��0�/f\�N������Xe��� Ay����?N^�?n�?���� #�k6%?�>_����8Ǿ��<���>�(�>�)N>|H_���u>����:��h	>���?�~�?Qj?󕏿�����U>
�}?0̴>.Մ?o�>>7�>��>dX���yȼ��(>Z�=�p��$�>��L?7��>#��=I~6���0��G���T�H
��B��Ƅ>\zc?9J?TN>������^�!�jOｏ�!�v��T�H�AqP�<KϽ�c;>7>>,x>�fK�ՃоAR?����ֿ��گ��i�?���>�?Kzᾶ�e��a<4`S?�rk>��X4��ϥ�����h��?���?�O�>XԽ���h���]>84�>�Q6>t���0A��F�-�]>��J?&�Y��A���N��ঀ>��?�L	@s �?�
k���?�Ҿ����U2:�88������	9>8hW?Aԕ����>6��>v�r=;�}�!���.�r���>�p�?~y�?�k?�i?����:6����=P��>q>�?J?B��X�x�>s6F>2m��������C?@�@�kA?4�����ڿ���_��HϚ�_|��y1�=-f�>^S��?����<� >��d�}g�=W�g>l|<>��b>�;?>�D>O(>���L; ��ʟ��%��Qg.�_
�����@ý�Q߾6Y?�X��~���٤�L���.�v徽0�P�g|8�/�ҼB��=)cV?ˠn?O�}?iR�>��.����=���L���վ��pv=�%x>[07?�AR?�?k���˾�m�</��Ql����y���>0N>\aO>[�>,e�>EX�#0�>��=>/e�>�a*>��>��&>���=�d>��>>?\�>�R<>�>�д�2��=�h��w�|�˽���?ي��X�J��2���2��S����C�=�].?,}>x��@п�󭿶2H?����'�X�+���>��0?LfW?��>����U�;/>ó�M�j��o>�= ���l���)��Q>&q?��d> �v>��2���6�?4P�M���P�>��6?�l���9���s��I�ྜྷ�F>`r�>
��g��G����z6j���s=29?xY? ���(��Y�q�����{V>�\>�A?=)��= uO>V�[�w��}@�|�*=>��=ξa>�3?�_,>d�=��>�Q��T:O�б�>�@B>z8,>D�??�C%?��o���Kd���>-��<w>#�>���>��>?uJ�ȝ�=�9�>�Sa>?���-�� L���@�8�W>��}��]^�6Nr�+{=�s��Ln�=[��=�n �]<�el(=�~?���(䈿��e���lD?S+?] �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��L��=}�>	׫>�ξ�L��?��Ž5Ǣ�ɔ	�-)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�e�>
z��Z��5��K�u�+�#=N��>�5H?�V���O��>��v
?�?�^򾂨��_�ȿ){v����>��?��?!�m�B���@���>9��?_fY?7gi>�g۾�\Z�e��>!�@?�R?��>8���'���?Fݶ?���?�X�>7��?}l[?�������>Id/���ο�M4�\J�>�n��d>��#?�����1!��yۍ�����#R��3/(?�f�<�H�>X��]�;}��<9I=͒�FA����>�?��C>�`�>{9p?4$?:1i>Z���9#>���k���K?���?B���2n�+e�<#��=Ƿ^�o&?^K4?�[���Ͼ�֨>��\?~?y[?�a�>����<���翿�}�����<��K>�/�>�F�>����LK>A�Ծ�-D�'o�>�ϗ>�I���@ھ;*��xk���A�>�d!?7��>�Ю=��?z�,?2R�>���>��!��7����_�2��>0u�>��>��l?$2?r�ž�H@�K���]���df���h>�b�?�?��>ݍ�l����N=1ՠ��q � Ӄ?�Mu?W�����>�%�?��B?�7?� >̜��0��?-���,�>� ?�~��@�L�$�����?�?�7�>�����1ؽ�X��8,�=k����?�[?t+&??����a���ľ�W�<�E�4p��<��;@�;��R!>�3>� ����=��>�5�= f�{[1�"�<>��=(o�>I�=�6������0?,[G��R��=�=�>��B�J�x�|>6��>(�ƾhA]?�!��"݅�[���ѭ��}1 ��Տ?���?K,�?b¬�K�t��L? ��?�S?��?Je}�N1��S��
���-���~��>hJ�>C+D�
G!���9ə��p�/;h��0��p�>�S�>(a	?u�>=�w>G��>�1׽:�4�[N㾒���c�w��c9���G�9`��O޾�V��&㤾��=�6>ƾ�99T>X���$��>[�?'�>�����>�g�<�o?F��>���>���>�im>�ܡ>���=�$�����<�MR?������'��������YB?�yd?/B�>H�i��|�����1�?�~�?Bd�?w�u>��h��5+�K?ք�>z3��Ë
?z�;=�D���<<���K8�'V������>��սc:��M���f��G
?�?4:���˾�.ֽ�����p>`��?Z�$?:����O�t삿��S���?��h������O���,.��t�Wk��8ʄ�	��l���r�=h�"?��?������O�[������v��>�>�?��R>��K>}�>�ѾĻU��2v���)�c�Ǿn& ?�{�?��>pF7?W0B?�_?u�d?tb�>E5�>���Rf!?���L ?�_�>�K?$r?�?�P�>V_*?�W?�XC���Ҿ����[-?ҸP?���>�ܢ>=��>}�-��I��ay��ޙ=
��Uҽ�2A;�H>�R1�%�ؽ\����#>3X?�����8������k>�7?�~�>���>�	��M)��J.�<��>��
?vO�>����|r�5_�]�>!��?8��v=��)>���=l���Ѻh�=����ܐ=3m��.m;��_<쀿=�	�=�t�Uo��4��:3]�;�ɯ<�t�>Z�?瓊>�C�>�?��g� �Զ��f�=|Y>�S>8>REپ�}���$����g��\y>mw�?�z�?��f=��=���=R}��.V��G��Z������<�?�J#?;XT?��?��=?rj#?е>.+�HM���^������?�r,?:.�>p��/̾�X����2��?c�?q�`��\�J*�l��Gν�>�/�x"~��̯�N`D��.�;f&�����'�?#�?O�Y���7�|!�e(������C�A? ��>մ�>5��>�)���g��6�c&A>|�>��R?���>f�Y?�gv?��D?gņ>��5��V��Xo���О=v?>�f8?,;�?��?րt?�ٖ>�ɠ=��!�����6��g�c�8���G{�W/�=(?2>��>�>�>��=�Z��'���v�,	>��[>�K? C�>1��>̺f>�<����G?#��>�R�����䤾ﺃ�,+=�͚u?���?��+?�~=�{���E��0��K�>]j�?���??7*?��S�G��=��ּ�߶�i�q�� �>��>n=�>���=��F=�c>��>P��>4>�qX�^p8�M-M���?�F?���=a6��Úe�����>)澏1�����.l����ʊ�*Gu>�8��D�ƽ�����s��;}�ߓ������6��3���?���=�{��3K<��<8�<�7=)�?�*�?�����١=u����o���jo�<Qn�;m��<� ���˾I�|?��H?�,+?1�B?��|>y�>��A�P0�>�o���/?�S>FLY�����8�&������l%پ��׾rd�����3�>�/N���>�4>���=4�<��=:5r=�R�=	�f91&=�
�=WR�=,0�=���=��>f>>2�?�N{��I��C�뜘�{K�?u��>
똾;q��z�?g���8����Z��wG���o?C��?�f�?pC?��н�u>�l�����=��*�w��=)�8>(w�<n琾hz>Q�4�Ā�������i�a֐?~	�?$Y?���1��S9a>�72>�-	>�P���-�z�]�9�X���I�I>#?�;���˾Ҋ>C�=���6˾_N=in;>e==-M'�v�\��B�=8@����+==�Q=�߈>4P>�Q�=��ܽ' �=��Z=3=	>��Z>8��;~x ����7q=���=ك`>X�->���>?�i0?^d?��>�n�/Ͼ����'��>�?�=�T�>ػ�=D�C>��>��7?�ZD??�K?�|�>�=6�>Q��>/�,��m��#徆
��霮<Es�?�ц?�!�>��P<�B�%���!>�ӤŽ'l?ie1?	�?>�>�Q�Jɿ�㾖���KU�%�����9>1�=�K��:����PR<�b�>=�G>�g.>�K?>���>���=���>��Y>P��)MB��'=B=HR��;�<4���m��=�5ٽ�g�M&;���;��9���=۟��ϔQ��⼿��=�'�>�	0>:�>էF�ӻ�7�0>��%���o��i�=� ��_�\�Vas��Ex�{��3�;�2>9w>�K������E?�v�=��>D��?�Ue?&1�>{�I���/w����>�y~��<� e��-���QE�Ӻn��of�!��2��>&ݎ>ɢ>��l>#,��$?��x=$�ᾕT5����>��������X-q��=����i��7ݺ*�D?]D���c�=:~?B�I?;֏?'@�><ߙ�s@ؾ`�0>C���{=7���q�_`���?i'?���>F��2�D��	̾oZ���\�>�I�� P�(ϕ�׆0�w�� ���W��>�Ҫ�<�о�3�	e��e�����B�0r�{�>G�O?Ԯ?��a��P���O�����V��j>?�kg?\K�>�T?A[?녣���#��Rj�=�n?���?S�?�i
>�3�=����(�>tY	?9r�?k��?�Cs?>#A��H�>�v;�6%>T�����=��>��=#F�= ?�B
?�(
?x���:
�ϟ���x\���<g�=�w�>]�>��q>
��=cyp=�q�=Ⱦ\>Z �>ԅ�>�Ve>��>pԈ>�7���t�X�?�7>$;w>|�^?-)�>���=�#�� ����>	S��}���A����=Cy�=#����Ľ��5�mS�>�Tƿ�?	,�=]�H�c?�� ���>@�T>v�=N���ʎ?���=g[�>�b>�O�=x�U>��>w%>�dǾ�>S���	&�n�C�T�N�R��� .W>�ʠ�W�����W0ܽ<�}ݴ�s���f�H���n�B��T=�?���\�f���%�|��
j?�<�>��9?n炾�U��p�>(n�>���>������R���D߾C8�?5�?�;c>��>I�W?�?ْ1�33�vZ�,�u�n(A�-e�V�`��፿�����
����.�_?�x?2yA?�R�<-:z>R��?��%�[ӏ��)�>�/�'';��?<=u+�>*��.�`���Ӿ��þ�7��HF>��o?<%�?wY??TV��6��tI>�??��f?���?47?4�(?���oD<?6~=h�7?g��>ȡA?^?�� ?!d�=�#>NQC>�A�=+l��,a��^V�_>�6u=�$��Δ=c ���Τ"<+�;=E&��a ��]5�{&����K=A��=���=�,8=�ڦ>y ^?X��>dM�>�7?���C�7�C\���0?CD=I���鿉�ݽ��:��=�>h{i?O��?�O[?w�`>��A�faB��>C�>�%>��]>�*�>���E�Kσ=��>��>�=�=�:����	�Z����P�<��">�&�>	u>�/{�< 0>N.���Z����`> 7��ÿ���>��M�N�4�*.��C'�>��L?K?�'�=�v�$'��~Qi��,?�;?\HJ?]&�?�^�=�r۾:5���N�M���S�>�0=���o���3��l<E�Y�-�˶b>?U�������4^>;��B�Ᾱrj�>N�q�Ӿ8vQ=x��s=@�7�پ�+d��*�=/�>)2��c�#��ɘ��ʩ���M?$ڥ=�U��σ���rо@>��>��>P�4��J{��B�zʖ���=E��>3�;>#�����.�C����ȯ]>z�??�W?{o�?F拾���w�7����챾ҩd=�I�>&��>i%F?*�
���������L,��%w�!(�ݭ�>Y� ?;׾'�Z��¾U3�Q�^�c�~=�g]?x����%>??i�?޽�>��j?є?}�?c�|>�ȣ�~!��� ?���?���=��!��Vo��=��R����>��=?l�_���>�`%?��0?��9?��F??���=a� �p�U��P�>��>ȕS�;8����|>8Q?���>�#Z?��c?l�-> �@�sϷ�Gsƽ�� >F�d>��0?�?K�?>d�>]��>�S����{=a��>�a?Z@�?��p?���=�?w44>��>w�=I��>oS�>?�K?<�p?�L?��>�2u<Fṽ2���5��?�w(ٻ��/<��w=G1�'�g��g�(��<я�:�Ҽ�Cn�B{���C��wq�<�t<���>��t>9o����,>��˾L#��_!G>y�l��*���}����A���=h��>�� ?��>��$�J�=� �> ��>�)��g'?��?��?
���Ga�6�ݾW�J����>��B?NT�=+k�͆����w���O=U�m?�Qa?��L�-A���h[?q�f?	�ӾB�8�
�о�I���)��:?JI"?' `�4��>r�?��|?�7?�Z���h�N����~[��$���H�=���>�Hu�֧>�7?_��>҉>Tt=P̾��x��Ǻ�!`?�#�?p��?���?]�%>��]���ۿSz���z��T�d?���>�㢾�%?w��rsھ�ɏ�����׾����ß���K��˂��9w"���}�t�߽�]�=�!?Mv?�s?j{_?:����d�-Z�ػ��)Q���	�f���8���=��?��r����7��FC��7��=6[|���F���?5(?�&���>Jn���,�Ѿ��>�h���0�X3=�O�ZcT=7�V=��O���/����ض?�|�>�1�>�??<�T�|:���-�tD��'�)K�=O@�>Ҡ�>~��>4�B<�&X�� 1�x���_��l���	+>LjZ?B;=?X��?����Xg���i��޾|����޾��8<N�={��>�A��f��?�E��}N��a�!^�w ��

��W�=;�D?��>�i�+ɬ?��>N&e�]�<�Vƾ��Y���<>���>�%f?U��>�Σ>�����m�T�> �y?r�?+� >%�m��i��<ϐ�����<8?���=�i�>���>�����1�����8���t�q��Y{=��?�ł�<B��˻-����?�sE�����FD>D!�>D@ӾV�$�n��Y�>qB2?7Qn��>�	0��<���R��-�ɾ� ?j5?�bk���6��+j>3-?��?���>��v?ܬ�>nC����=��?�Mn?X8=?p*-?�9�>tU�=x��r��I�i�#��&�>/h>|��=��E>0�ͽ�"���սW(�=x�\=�S���Ķ����T��	=��=�A�>�οy�H����������y���
�������؜�����˾}���x(�
�"�j�o�1J(��w����$n�wC�?fP�?=2����ɾ���d�������p�>�E�a�)�ʾ�(�������� xh������^��v�q�o���$?�W����ǿ�O���q��s~?(T.?{?zZ�}v�dcE���*>��@=o���D�p̖�;�˿���Y[U?�"�>G������K@�>N�'>�R>��x>�2g��}����>=�t ?��6?���>�����ȿ��3Ja=���?�'@XA?�g(��i�!R=#��>S�	?Y8A>��0���^԰����>{.�?q�?�bV=zW���
��Fe?��<��F�$�ԻM!�=v�=H�=-Y��EI>篓>#��O|A��l۽��5>���>#(������]�Zֶ<Q]>x1Խ',��!�?�c��e���Qw\�	t�>A/?�4�>5�=�o?W*��ɿ�h���>?lD�?H�?Qz.?z�о���>&�ʾw�I?��*?�x[>����i�w�N>C��a�=�Y��Fj���>��>���=Ց�����|4!�ʴ�=��>{���Eſpm+�����=A<' =c����(=���F��{,�:ϧ�=��Q>��>��4>��e>�e?��p?v�>��=��<���C��s'p�fp\�<�E�W6�����K���z߾��˾f� ��S$�����о�3�LZy=b�Y�	 ���=��tg���-�[�"?��>R��U��4� խ�����}�T�@1����ݾSC�M3p�o�?�"J?ϊ���oj��'�>cp�	.ȼ��a?K�ʽu>��6Ⱦ*>�`���t�=�Ĝ>:��<���w0���L��f.?0�?wʻ�}��#�+>oaؽʐ=a|)?8��>,KU<�r�>��&?́�kIv���]>0�$>Mѡ>Da�>y�>օ��P���[!?��Y?�"��ɮ��Ɛ>���L�n�*Iq=VJ>��,�l	R��n`>��<<,��Yy����q�+�1=�'W?U��>C�)���e_�����Y�==+�x?a�?`,�>	|k?�B?��<�^��x�S�A��dw=1�W?$(i?'�>[����о�x��M�5?�e?b�N>^h����a�.�UR��#?��n?k_?�f���v}����\���o6?Y�v?�]�Թ���q�ie��!�>ł�>���>>@6��λ>��8?��'�^Ɣ��꿿�2�
ڞ?��@��?���;�� ��Vh=���>0��>"mC��n��4������ �=~��>~S��	�y�/��!�$��P:?Q��?���>��~�������=W���1��?|j�?#����=���(_~���K�0�D�>�_�<"����nҾ/=0���̾��	�n��Y�C��i�>��@�ɽd��>����c_���w{�w�ξL#;��
?��>15X�e��󓆿-󄿕U�P��+���[�>Э>)%��� ����{��`;�K��B7�>���yG�>�NT�?7������k�-<�͒>���>4�>���������ę?q��<οW������n�X?-Y�?]j�?6l?X	5<�&w�|���_,G?��s?�2Z?� &�{]��B8�rj?"����`�x�4��G���P>��3?Ȗ�>��,�1�=�l>�t�>1�>2�.��EĿ�h��xC��%�?�>�?S��Q	�>b2�?�+?�\����Jq��c3*��m?���A?�V5>7 ��!�#�Y�>��v���
?c�2?Jv������_?m�a�H�p�
�-�a�ƽyݡ>�0�~c\�eL�����aWe���vDy���?9^�?s�?ײ�#��5%?��>뜕�8Ǿ���<��>�'�>�,N>�E_�V�u>����:��j	>x��?�}�?�h?N���x���ZY>��}?��>/ф?L��=� �>v��=�7���h">_�=\�8�""?RM?e[�>
/�=A[9��1/�t(F���Q�r�BC�4�>�a?�L?��a>�巽Ȏ3�e� �=�Ͻ'0��L뼨f?�W�(�nn�d 6>�?>{>�HF��)ҾT?p���~ӿ]R��u۾�k?���>?W���ƽG� ���b?.x>���l㯿𽃿����\O�?Ii�?�l?��о�#x��M->BH�>4��>��N���l�#?{����>CE?l��DI������7|C>]ֿ?}@SM�?#sV��]?��f�Wt���F��):��wV>��L?u�־u��>�ϊ>(�=�+q������n�F��>�r�?ba�?*��>&vp?��z�R�U� ��;C��>��?y�>��s=����T�<>�=�>z�N�ɻ������x?�@��@E�s?�\����ؿ����{���o����X=���=�J>������=݉��9���!�;�/�=ۆ>�Gh>'�D>�K>�V>��1>*���W{�ǣ��.����JE��*����j4P�)����B���'�$����о�(���߽֩��>�"���魼�=�T?qqP?:
o?�O�>̭ǽ�=(>y����x,<���/W=�>��7?��G?A"?M�8=����8�a��[��<��g3���ؾ>:>�h�>n!�>���>�"���-.>�N>�q{>�%�=��<�W=��w:=G&Q>�ީ>W��>�>�>J�>>0>z���糿Ӿl�����?ָ<���?ͣ����6��ߛ����h=��4	�=��!?���=^ې��*п����yH?�h���bZT��JH�'?ykd?��{>�M��|qȼ	,�=�e�;)�A��a�=�z*�k\��	Z���Z>&� ?�h>3u>�f7��P<�}�V��U���$�>�8?�߶�^U-���z��\C�I*Ծ��N>&��>������Wp�� �{��c�<a�=�G8?�R?�$�<���^�i�Z瓾�Q>[�f>8�=$��=��E>P���k��ôP���r=��=�;y>�?sb,>�7�=�
�>��	rI��ǭ>HXB>��1>�??n?%?lI׼Nz����w���(���r>xe�> ��>�I
>��K�F��=<
�>=if>�{������$��y=���U>��{���`��e���n=���_v�=��=P���V:��.=�~?���(䈿��e���lD?S+?_ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�g�>Yu�nZ��\���u�פ#=[��>9H?�T��c�O�`>�w
?�?�^򾫩��	�ȿw{v�=��>��?���?A�m��@���@���>e��?�dY?�oi>f۾�YZ�썌>��@?�R?/�>Z:�g�'�s�?߶?���?��>�"�?�L�?�.=�>�f)�U���5����{��9S��Z�=����W��X���w�������~�<��>���=���>�p�;��>�G�=H���,�}����>Y�?���v�v>���>�e?�7>0��-*���������=,�8?J�?�׾�	��?�����=��g�g�>']C?0�ཉ���T�>6�n?��?��M?��f>+=�B��0ÿYH��z�ƼN	L>j�>��>b?>��>~᫾����>Wk[>kf���E�wv���ɼ��>�U/?��>�0>ˏ?%].?琑>�g}>�-�������N����>o"�>�A?PIh?�K?�6����辕�u�����l���>��?�?7т>�!��ь�DU���u�<����\�?YCo?vN,�ф$?i��?�P?�?bil>�䩽<Fþ&�V�n��>SV?}��?U�sh�G��=\cZ?9���,�>Jk���Bˡ>C�b�\Qa��D�>Q��?ρb?��۽����ϸھ�ד���<Ǔ�<I�=����g�>�l>��\�@={��=�&�=f��� ڽЖǼФ�<�X�=ج�=>���a�8��7?��}�1[��znA<<�~��+���>Bה>ĳ�5�i?+v�4�d�0L��'˞�}8�"!�?� �?��?�3o�Ǝs��3E?�?d=?H�s>�7������Ӿ茶�Ō��yѾz��=$�)>+pc�H �6Ե��#��2so�B�}�
_3�5+?���>S�?C?ù(>�	�>>�����1�ߣо������c��&��h?��� �_��p���~s�u9��bϾy!q�y��>�ږ�р�>J?=jf>re{>}�>���ϓ�>�3V>�^>�M�>Ꚅ>��_>���=/8�<�	�=5R?c~��Π'�U�辒��L=B?P�d?)�>wHi��t��Vz���?~�?���?{5v>xch�g+�7�?��>����*
?�6=�?���p�<�����*�V����I����>�ս*�9�- M���e�c
?��?��	>̾Еս��u�>#-�?B�(?����N��e���^��Y��\y��7�uЂ���#��9c�ұ���U���c�����:�=d�?�"�?Ť�Z������Go��i3��;V>ߎ�>$!W>n��>)��=��߾U/"�v2r�0J8��s��%?Q�v?�~{>��4?�7?V2A?�b<?~��>�"�>dZ��I��>t)<3X�>�1?v�<?�#R?"T?�n�>��?��>�P���F��0`%?��$?v�?Բ�>g�>�MV�������&Z)=DJQ��}9�V�&;%*9�'o<�=��	</w8>D�?�"��7��`��Ϙk>�6?���>�W�>�ꌾ��}�3�H=���>��
?�y�>�a���bq���
�m��>:��?�&��.�<"�%>j��=j�]��0���=Q�ؼu��=�v���7���N<ȳ=+�= PF��c��O:'����;__�<v�>��?S��>/=�>|>��Ч �%���]�=�Y>�S>�>Dپ{|���#��+�g�	\y>�v�?Iz�?"�f=��=���=<w��LZ����'����<ܞ?HG#?�VT?k��?��=?�g#?/�>�-��N���\�����ǫ?�x$?	p�>�r��Y�&��z�7�t(?�?��Q�𷇽As@��,����x��>N�.�Vt��L��/�J�o�=Ӭ���Q�Q�?�??u��:*�dz���抿����IJ?��>�l�>%��>�>���r�c�מ�>�?��Z?|�>nhW?��v?�M?XV>��>�'��Uږ�
��=���=]�J?D�?�?%�~?���>V6�=H���ڷ
��������;��I~E�Omf>O�>��>���>���=�)���4���e�;�=?��>���>̨>�f�>�L~>�U��R[?�u�>W>߾�u�شt���S����e�k?L�?�G/?;{�hM���D�	�;��>߮?��?*,?-��u�v=|��=p!O��o����9>F8*>g�>�u�=��>���>��+>���>+>�=
���#f��2㽖�?�b?�`�=ƿ��r�N#y�  ����<��86T��흽|�d���=�k����h���� a�p�������b�������tt��?�2�=�,�=.6�=E��<��޼_i�<<�=X"�<ǡ�<ս��`�<5h;��C:�6���J��}�:t�"=�<�vܾ�gj?�R,?��?�R?>4>JD>A=UO�=P]���F?a/&=L�9������ֽ��O���P�P8��m��"�{�������=�Tս�,L=И�=+��="/=@2�<�AҼ��>��=���=�v>[+>ʼ�=�>.L>퍁>�=�?�-��"��B��޽�=Y? D<> ��>-�+�ZCQ?�C��k��ϥ�����}u?VH�?S�?��>a,�3r�>�V���:>>��=]�>��>Bix���M�qo>���[�*�J@���ҟ���?��@�h8?�����ϿҒ>J�6>P>�Q�d0�JU� ]�j)\�uc!?�v;�J̾���>��=��ᾇ�Ǿ�(J=��:>�p=���Ǩ[�I�=��dNC=��f=z��>�aC><ۼ=�~��=��D=8�=�kP>�l5�1�-�G�)�?�1=?��=�#b>5�'>��>��?t_0?:Qd?y4�>��m��Ͼ;���F�>��=�K�>���=�}B>���>�7?N�D?��K?���>��=��>��>g�,���m�)g徏Χ��<X��?�ˆ?�Ѹ>�R<;�A����a>��&Ž�q?:P1?�k?��>�lpѿ�U����21�57��@��>���"k���=�Z=�oM��f�>�}>�a�>Hӊ>Э�>tG�=Aq�>��>�ƀ=2n���5>�>�
D=t�=��i�֣����>#ü�\���4�=�[㽦� �]D�=��=�l�x�ں:v�=�O�>�\�=y��>Hod<c������=R�W�rA;�S|>!����G�j�h�b؃�)��71��x>TV<>�v�"Z��k�?�d>-�@>���?�m?sԫ=�s=�:���� �*�ޒ���=�'k>볽C��C�i��H�	����>	�>���>�ik>{+��>���j=~�d4����>=���V�����p��S��c��o�i��B��7E?*���K�=�O}?k�I?%z�?aY�>"���Y�վ�/>8��E�=���7�m��e��w�?��&?��>̿�n�D�
̾
L���5�>q�I�"{P�4���]C0�b������(�>r���|Pо��2�zY�������}B�6=r�ǅ�>�O?�ͮ?cb�x0����N��������?�Ng?
�>v?|\?�S���p�~P��8y�=��n?���?>J�?�h>$�=$�f��X�>���>�+�?�[�?�v?1L0�=3�>U��:}�F>	v ��>��K>Xx�=��=��?W�?2�?ڇ�p��^B�p�Ǿ�L�+�~��*�=�ŕ>��~>Ȝq>f>>*"\=��=��o>��>��x>AW>���>�U�>^��*D���_*?:��=��>\�$?�BX>OT�=UX��'������=��~��q��B������[�=��=��=����>ο�N�?ȓ�>vZ���?��4|��k>���=��׽"?5U>(��>��@>�\�=@��=�f>v�f==�ξ�$>=����$��F�X�R�ՠþZ-�>�ɜ�X����Q��f@������&�C#h����Ho?�Eɍ<�3�?H���ti�\�'����Y?{I�>6?7?�y�p�Jn>M��>��>&��������J���)۾�]�?Z�?x9c>c�>��W?�?��1��3�RuZ���u��(A��e��`�H�������;�
����4�_?��x?�yA?�o�<8z>���?K�%��ڏ��*�>V/��%;��<=�*�>�&��}�`���Ӿ��þ/��<F>͑o?�#�?@[?xNV�17��*!>).?Y�[?��n?�l?Q?���|c?<�&>$uJ?%�>?9�=?^�k?���>uG9=��=R7�>��>��ӽj᣾��=�v6>Yq=7�6=HWj=�]<�]�=���=�3�-Z�<y|=&���Kh��!F�=.�6���==�X>���>L�]?0<�>@��>��7?X��1b8������/?�p9=	���P���բ���>��j?y��?�YZ?&d>��A�1C��>�J�>�F&>�[>
i�>�Yｦ�E���=�s>�`>���=��L�����j�	��n�����<�T>;��>�#|>j����'>����3z�S�d>��Q�
�����S���G���1���v��3�>8�K?��?1��=�I龅O��YPf��6)?$\<?�IM?��?n�=��۾��9�b�J�sK�+�>�R�<���8�������:���:ŗs>	F��ʠ��Vb>���zU޾�fn�<J�Y���L=q��AU=�*��!־>�����=1
>q����!����|Ӫ��J?�j=r���U�(^��_>琘>˼�>�w:��v��p@�Xì�4��=Ϛ�>��:>�(��g
ﾞG�rD��6�>�.E?�_? ��?)���M�r��B�m���C���&���'?ȷ�>��?��<>�â=������d��~F��t�>@��>�I�
nH�"����B����#����>��?��$>C?3�S?�C?l�`?a_)?��?֏>?�����?&?_��?Z��=s[ս�T���8�>)F�*��>�d)?pNC��~�>R?��?]�&?�cQ?��?%:>� �83@�!��>�6�>��W�ob���P`>��J?/x�>�BY?\̃?P9>>o5�f٢�{<�����=��>��2?�<#?��?,B�>���>ܩ���C�=p��>�c?A0�?�o?=C�=��?�J2>���>��=×�>d��>�?�TO?Z�s?�J?��>v��<V8��!��{*s��|O�O�;�G<k�y=ӳ�DWt��o�$��<{\�;	W��P��G��O�D�q����E�;��>)�Y>�y���>>��;����#N>�䬼"�����Ҿi��:�;=�b>V?a��>��e�d}�����>3��>�'/���0?�$�>�@?�?>�x��+��-w��*r>Lu@?<>�<�����ﭿC{�����IW?��'?��f�m'�}�P?B�v?�ˑ��_k��3=�.$D���q;?�P�>�"���>U�}?蚍?4ת>[���f�v����#f�0¾Z��=�T�>�G��xd���>(J?��>[��>?T>�|��������
?J�~?0M�?}�?�� >�%n�bcؿ�����c��v]?a�>|թ�~%?��]��7ξ-b���=���v�R��D媾�ɒ������(�$���Kn�����=7?-r?�Ks?T^?"`���a�Y6[���~�`LP�����$�o�B�XC��B�)�k��6�5������=�q�b@���?�{*?��?�lh�>������P�ϾJT�=h���?�I��=k���29=P�%=��7h������?��>ɭ�>�$:?�c��d:��L,�-�6�	&�X@*>��>�ۓ>���>�fR��>*�e��������ki��F$��:v>�ic?�K?��n?�� �f;1�(���|!�B�3����,C>��	>��>	�Y��r��&�|>� �r�h���g����	��{=٩2?y�>G��>�A�?b�?��	��%����w��1��.�<�[�>E�h?���>6K�>@4н�� �߅�>.+j?R�>p�>D���$��b}�*�߽�K�>`��>� ?+>��U��3g�m	��G�����-��X�=@``?���Y\��^�>�@S?D�S=�Z�:�^�>泈���4�j��?��� >��?�ʨ=��>DRҾ؎��bz�~����N)?�O?)ᒾ��*�<~>"?.s�>�1�>41�?+�>�jþ�<�ڰ?�^?�>J?/TA?�F�>dk=�6��_JȽ��&�Ԩ,=~��>��Z>�	m=h��=����p\��r�1�D=\}�=2ϼb���<�f�� �K<6�<n4>�ֿ�7�������������y���PT���-���?"���&��%����ڽ��>z���$�u����-S����?���?"�s�����L����㗿�=���?�锾����鍍����S���%��-J�`�9�%�W�2 f�j�W�C�'?����׽ǿӰ���:ܾA! ?�A ?�y?��c�"���8��� >'B�<�+����뾢����ο�����^?���>��-��~��>?��>��X>�Hq>���>螾}+�<��?<�-?��>�r��ɿE����Ǥ<���?/�@d}A?��(���t+V=���>_�	?��?>3F1�J�E��<G�>f;�?k��?�M=r�W�:9
��we?��<�F�E޻�D�=Bl�=y=��~�J>U�>m��wLA�(ܽ��4>�݅>kq"�����^�c"�<�]>��ս��NՄ?�{\�#f���/��T��mV>��T?�+�>D;�=�,?�7H�K}Ͽ�\�F+a?41�?��?��(?�ܿ�Eۚ>��ܾ�M?�C6?x��>;c&�_�t���=7�(ڤ���㾀&V�q��=b��>�>S�,�s���O��/����=r����ſB�7�I��G�<A�k=)�����_��c��Ԡ��N��^���ӽ"�>F�=5~?>���>�T>�ߘ>�X?�?��	?��>oGO��U��<��F�H=/ld�0�"�ȾH��V���� �cY�$h�;����!���վp=�S!�=�2R������� ��b���F�$�.?[V$>��ʾ��M��,<wʾ�����R������5̾u�1��n��ʟ?��A?g􅿼�V����X�����y�W?�j����ެ����=�m���M=��>$K�=����3�fyS�/?=� ?pi��I����3>�k��ͺ<#�+?'?�Χ<�}�>i�%?��%�4�󽄌U>��9>���>�O�>d
�=Ѱ��d�0A?�V?C�򽳤��K��>h�Ǿ���e=>�%-������Y>7�;b�������K1<��q(=�{U?J�>&(����I��4f���=�)u?P�?�Ԥ>Zdr?rE?{T=@���ŦT����=��R?�i?7�>ǅ@�2�Ⱦ����a�8?�ah?�A>�c�B��L�2�?J�R�?��p?��?k�c�)�y�s�����.E1?��v?�i^��o��!����V��/�>�D�>���>)�9�e�>o�>?t.#��F�����`Y4��Ş?g�@#��?d�9<��#��=hC?[g�>��O�r/ƾ�����{���r=E7�>a���4av�(���\,���8?���?���>�|�����5��=�ٕ��Z�?��?L����mg<4���l��n��Q�<�ɫ=t�)I"����l�7��ƾƼ
�|���0Ͽ����>Z@xQ��)�>�F8�6⿕SϿ���ZоQq�v�?���>��Ƚ������j�_Ou���G��H����\�>J�����SD���)��+S�B|н�lV?������>	jվ
���
��#\#���?y��>��?�{���^_��R�?S~6��Kտ����r۾�M�?���?�D?�)B?ra�̆��
�����=�e?�<�?4!�?wQZ�h���n�̼ �j?�_��hU`�ڎ4�pHE� U>�"3?�B�>U�-��|=~>���>Tg>�#/�k�Ŀ�ٶ�M���W��?؉�?�o�-��>r��?rs+?�i�8���[����*�-�+��<A?�2>���?�!�E0=�\Ғ�ȼ
?]~0?�z�H.�u?鳀��\���^=�Cҋ�N�>'N+=W��<�{�=V%��B��K)���u����?w�
@6��?O%���J�G�j?���>W�����I��X!?e�>\�=�>�k��=J�:������>�D�?W@?��>������%L5>�$x?"�>4��?��=K�>;�>�*��K�Ƽp.->��>)�=%?��M?�>���=�8�X�)���B�'S��C�,�B��ʁ>j`?O?k/f>�!��!�弃�$�D۽�@-�)�Ѽ4�6�3N���ܽ/�$>��7>�T>�'��už��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji���?�p��3��߶y�iM
�!\�E��=�]@? ���ф>x)�>:�=�c{��%����o�*�>;��?+��?̎�>��n?�r��1A���<(k�>Wvm?�=?��<lx澋y=>���>�l�R���] � 1s?b�
@�@�^?�����׿�2������¾�'�=L�->�">)R'���R<�,=�چ:��<C��=�9�>Ӽ[>�n>G�A>�V>�~F>�����$��3��q���MDB�Y������(���a��R�O:��I��i���Y�	�C�+��3�G���b�; �=��W?��Q?��k?�?)����,>����\-\=����[�=	��>�/? -E?rM%?��=>���'�c����9����I�����>�J^>��>�K�>��>D���&8>1A>-w�>�>y�	="�v;=}�<DaD>z��>�,�>���>�C<>e�>Fϴ��1��y�h��
w��̽2�?f���H�J��1���9��⦷��h�=bb.?K|>���?пV����2H?;����)���+���>��0?�cW?��>����T�:>D����j��`>�+ �Hl���)�5%Q>�l?��f>u>�3��F8�D�P�p����4|>�6?�\��g�9���u���H���ݾ�]M>'��>�AK�4���ܖ�4	��i�c{=�U:?ˍ??ɲ������v��V��Q2R>�K\>ɢ=1/�=��L>$ d��ǽ��G�ئ,=��=9^>�Q?�",>�-�=��>�K���uP��$�>CbB><G,> �??%?�}�M����ȃ�}*.�yTw>a�>"�>*�>�[J�+�=�}�>�<b>Q.�be���|�|�?��1W>��|��,_�M�t�y,y=����-�=���=l� ��<�WD&==k�?Y����]��}��K=\em?��,?к�>
��rd��b���m�g��?X@@6ܮ?�<�MBI���9?)'�?��ὲ�>H�?�"�>Ou����' !?!������Z2-�G>r1�?�s�?9�Ҽy���R���^�=b�\?*W*�Qh�>Yx��Z�������u��#=D��>�8H?�V��U�O�>��v
?�?�^�ߩ����ȿ7|v����>U�?���?\�m��A���@����>:��?�gY?poi>�g۾]`Z����>ϻ@?�R?�>�9��'�y�?�޶?ѯ�?��K>�?2+r?;2�>�uG��/�m����w���ƛ<h%<q��>X
�=��ľ`�L�����Vl��g�c��+��HP>)1=�7�>P�齹ڸ����=�R��,���G��ب>�X�>�9X>�˨>/�?���>m��>�X{<�q��r	{��풾6O=?�`�?}ើU
��Ւ1>�N>�����v$?�yU?5
*>�gz�}|�>�ih?_I?��C?��>I��o���Zӿ~���7λ��">F8$?�B�>:���X=0J�������<>��>���<����غ�����G�>z7?�>�>�W1>\<?�'?��/>�#�>�G����2�b
�>�c�>�J-?w-�?�?���_8�4��$~��n|M�_8>�d?��?�d�>[Ї�}ж�߂��l<�w��fe?��g?P���C/?G`�?;�H?ʈD?iW�>4܃��;����z�>��!?���W�A�XB&�����^?�=?��>_!��$?ֽ��ؼ���h�����?�\?e+&?:���a�þM��<�$�rY��m <�D�;�>�W>����ʴ='>`�=�hm�BD6��-e<�W�=)��>���=X7������*?VD:I|x�䎻=3mr��6D�%Vc>�"E>)���\?��1�S��0_��@흿��Z�e�?��?�e�?�ڞ��Gf��09?^��?e�?�(�>�r���־EU�F���{�9�
�4�	>7!�>e���ᾞ���f�������ĽȽ��>��t>�e?�?��<{{Y>y��M�[������ �%rq���*�5�&��;!�&��;��\���<�:�����^���ܗ>X��<�Nu>��!?�!>��V>�>UwM���>�VP>�[�>�?�>���=[>	�I=�Hb����a^?�c� ��ƾ�_��ތO?�?jI�>X���������H?�%�?O�?Ӓ�>�Y}���&�q�#?���>s��VD@?�e�=)N�<TYT=���vϜ��m���l�22�>���?�J�#Ro�������>��-?X�ͽlUƾl����=���?�"?g�2�,GY�ٟn���Q���O��\*�gua�X
��wk$�\�k�GP���������aX*���%=t+/?���?ح��>]�#����o���>��ȋ>��>#��>�_�>�R>B{	��X3���]���*��恾��>j�{?ܨ�>[:T?��??��B?7sQ?%H>��>RS���Q?�I�=T�>�?H�+?lS?!�?�]?�*?�q >>�.�<����uྈ�?M�?�?��?W!?��ھe���=�*=b�?��/��l�=������>v��=./�>~W?���8�����k>Z|7? y�>(��>���/2�����<��>�
?�E�>F  �V~r��g��U�>z��?��=�)>���=����̺�I�=�����=LL��q�;�~<���=��=>�t�Gl����:䴆;[*�<�:�>7�!?j��>��>/Ǥ� ��"x(�Ǡ�=)��>`i�>>�@>Z��PS~�2�����g�)��>35�?q(�?H��<��x=kN�=�Χ���k��{��ʾ@)�=���>��>bM?�4�?��5?h?~}�=W_�Uݒ�ۀ�����%?�,?�b�>���spʾ訿�\3���?�J?�8a����D)�)�¾�ս��>]K/�N"~����K�C��&�������*��?���?A�C���6�lb�/�������{C?w�>�T�>���>	�)�+�g�����;>���>	*R?p#�>w�O?�;{?M�[?�mT>_�8�t0���љ�Y�2�2�!>[@?/��?��?�y?,p�>��>H�)�/�2W��-�����݂�V3W=
Z>��>�+�>d�>"��=��ǽ�Q����>��\�=��b>���>W��>��>��w>���<�]<?���>	7¾V�"�5/���Ъ�#�{���M?�X�?�#�>���x:��!R�°	�u�I>���?c��?�=?,ة�O�=[�@���!�����>v��>�I>4�->���>�j�>��>��>-}ؽ?)��`&�C(;<�?�\M?$Yz�w�ſߘq��Gq�E����;l<����e�Q1����[���=ۘ�����쩾
�[���������n0��n���f�{���>�.�=��=px�=��<F�Ƽ��<08J=���<R�=/zo�B$j<H�8��л�������%Z<*�H=�X��\E��xRS?��`? �C?X�O?���>���>W�̾���>}�p>Q�0?QW�>󉚼����#����)��mq�9Q���ɾHv�P�;b�=�[�=��=��[>��t>�����V�<j�=���=�s��vL ���=��s=�<t�=W��=>N>inw?E������.�Q���	�
9?Q�>ׇ�=d����>?X'>���׸���
�� �?��?Ç�?��?�J[����>o�����ǽ���=�V��s�A>���=0zG����>�Z@>���F��j#���=�?D@P�@?�����RпP�A>�48>�)>0S�G0��aQ��}j�:�[���?fW=��2ξ�u�>�#�=K��4ľ��(=g2>�j<=���\\�gq�=���1=a�u=z��>�%G>���= ֱ��{�=�rX= ��=��H>y�⻯�F���5�g%6=DH�=�T\>��>���>�?1�.?&Ub?��>�o�a�Ѿ�Z���`�>��=�)�>��k=�=>��>s�6?v�E??FL?�ĳ>O��=W�>�O�>7�,�@�n�q�r�����<��?4^�?��>1�Q<Bw@�>_��R?��iʽP�?e�1?�}?�>�>C8��z⿁su�s}=���;��>�FH=�Ծ>#5>�R�=�s!>��>���><L�>�ʐ>��>:�,>�<�>-u�>��=|����5>0�ѽ	=��;Cf�<��<�$�N�;-�=���:��=�?�'=u�<��=.g�����=�=92�>�e!>���>f@�=�7ξ:��=<�����K�魴=����@N���j��Ѓ���+���2�ܚ5>X�`>�������%�>B�C>B�y>U��?%�^?CK%>�%��d	��=��%zJ��^5�kݐ=��=�R_��I=���f��N�@��i0�>2��>�O�>k>6�(��D@��%v=c6���7����>G���/w:������n�N+��(����Ej�
D�;�B?�����=l{?P�I?,ŏ?@[�>�ا���پ.&,>�|��}="�&�z�9L��V�?`�%??��>[���E�×Ͼ�,m�A��>��2�<�Fک���@��2>(�澞��>�ӈ�Q𞾍�B��넿흑��X��+!��ƙ>��[?��?������a���+���ھp�d�>ˌ?s�l>0P ?y�>Y=�Vg��˾��|>KKn?�4�?"��?"8>Uh�=���e�>S;	?־�?ķ�?��s?��?�t�>�0�;)� >�U���"�=��>�D�=&@�=�h?W~
?��
?V�����	�ܼ������]����<<�=dz�>d�>2�r>
>�=��f=F �=�\>~ܞ>��>9�d>0�>�7�>�����3��
	?�[<>V�>�6?�M.>/w�<z�^�l$?�â�����A�-�/�d�ǽ>E!���N��+�=��߽	2�>R]����?ߴ�>�;��7?���`��H��>����bM�Ow�>�~>r�4>��>p�>Uˆ>W��>\��>UD��*>���������Z�7fh�ܾ(��>R��� !��j��{���X_��a���`��>s�
k}�4�?��(=V̒?��ͽS�Y��%�w/�	�>�6�>�P?����cP�<+�(>���>�~d>�������i���l5ž���?)i�?�4�>Y��>�&.?�?gᲾ�	�4�T��6a�G�%��G���6R������@i�K��P���q�^?�T?3a?s�>P5~>Nt?��0�m����>2l<���/�~�l=SH�>Uk������;�ݵ��#���o�="�|?���?>��>W���ˆ���>��m?*�p?�u{?�B7?��u?�L ���>c��>��?��	?���>�+�>��R>�}G>��=j�R�Y�=i|��6�q�@</D0�6�\<��~=��p=DV�<���;� �:yM��4 ���;���<�7�<o�=�3j=Hc�=T�,=��>,�V?���>�%�>;�? �/��:P�咾KU?��=1�i����pǾ�C���<�{?{��?��k?Es>TH�RB���G>��>�K�=X=7>{Q�>Յ�� w���=��p>�R�=��=��M�f�Z�G���8�?�c�\>y��>ٽz>����#>"������Va>�WP� �ʾ<nf��J�83�������>2�H?�2?#>={�۾_ޝ��cf���'?�5?4�L?�r�?_�_=W��D�9�-�I�Y���Ś>]Ώ��(�va�� ���>'8�����\`>|T���a��^�`>V��!ݾ�,l���I�X��B=��J=/d�#|־)/~����=á>¾��!��G��\Ӫ���H?d�h=p�����O�b����M>���>T�>�� �Ϸm�9s?�ꏬ��ڕ=� �>�$9>ҡ��N��OG��O�%9�>�LE?S_?Wk�?���>�r�5�B�+���MY���,ȼ=�?�y�>j?"B>W�=đ��q�m�d�G�N(�>��>�����G��1���)��S�$����>0?Y�>��?��R?��
?�`?�*?:D?J#�>{���#踾�A&?+��?��=G�ԽD�T�t 9�HF�z��>��)?^�B����>"�?��?��&?�Q?��?��>­ ��C@�ɔ�>�Y�>��W��b��"�_>q�J?嚳>�=Y?�ԃ?��=>*�5�ꢾש�&U�=�>��2?6#?7�?���>��>c���j�=���>�^e?�y�?L�n?���=�F?��->�~�>Lv�=�v�>Օ�>�?j�N?@�p?M�G?��>�r�<m���ӹ���w��;��u���[<�v�=�*�0�����$�e�=k Y<J߭�$�#�KyڼD�J�Ώ�IFF<{�>�2>,彾q�{=I���s"q�u��=|68���i�ž�-����=K�>	�?ɟ�>���7b�(i�>we�>v�4���P?*4�>�j"?Q �>(ec�	�	��h�ʸ�>�]U?w��=���}���f7{���=D�Q?s)?D�|��)�^\?�l?�R׾�n�hI��pM]�O�����?��>O�^����>:%�?�}M?u{�>����l����a��5�o��;� =]��>.?�g�)���H>5�-?́�>���=<+>���b���6����>
�?2��?+Fz?�ރ=�{��~ҿ�M����{fO?Mn�>.%����"?�ۤ�G��������� 徃ի��٠�e�i��n���=�H֓�tr��}h�=v�?�{?�Vv?~�H?*���^��+L�E�q��\,�W�5�z�G��	L�C�I���a���f���x�V�P��=?���0==���?��*?=(�`B�>>j���l��"B����=>Ķ����
�O��=)�y���$=���=�`�m�4�T1����"?���>#�>��9?�8S�yM7��,��q7�����؞ >���>��>4j�>���<i�#���ͽ����p��t����v>q�c?�uK? }n?G�1�s���~!��/�;���K�B>+g>��>+]W�����.&�>�,8s�e�:k��|�	��c�=��2?�/�>���>�>�?/�?18	�+⮾H x��j1�
��<�T�>�i?^��>��>��Ͻ{!�k��>�el?���>0�>�`��;� ��|�������>��>Iw�>Z�>�6�t[�(��������<�A��=�lm?hx���"H�/�>�@H?LW�;��=MZ�>�'���j�q:���4���>4?Tȴ=`�H>�����B��|z��3���O)?+K?�璾ä*�:~>�%"?*��>�*�>�0�?*�><pþ�XB�d�?��^?kAJ?qTA?�I�>��=�����6Ƚ@�&�_�,=A��>��Z>?m=c�=ܾ�u\�3x���D=x�=��μ�O���<�����J<���<��3>�Vۿ�:K��yپk��I�) 
�&F��],��#p���	����2!��Z%x�+���'�'�V�q�c�����Cl�a�?�,�?�쓾/������ˉ���}���d�>k�o�G�}�n��,��r�����ྛ���W!��O���h�pbe�Q�'?�����ǿ򰡿�:ܾ7! ?�A ?:�y?��8�"���8��� >lC�<�+����뾪����οD�����^?���>��^/��~��>�>&�X>�Hq>����螾1�<��??�-?+��>~�r�1�ɿh������<���?,�@�|A?�(�_��V=+��>0�	?��?>�C1�7I�����P�>;�?5��?��M=��W��
��{e?b�<b�F��ݻ�!�=wA�=�C=�����J>�X�>���eA�Wܽ3�4>}څ>%\"����+z^����<��]>��ս�<��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�����{���&V�}��=[��>c�>,������O��I��U��=����6ƿ)+$�'��)��<�%;vx�0��䫽c�t��w��ho������|=ȯ�=SnL>���>,l\>�Y>�BW?j�k??;�>g#>(�?#��Ӝ̾����Qy���_y���E�%Ŧ��8��"߾Tk��u�:��ž5`M�]K3=�.L������B%��`�&\��,5?���=�ݼ��S�V�fپ�亾7��񦳽ӷ���J)�\c���?(?�����W��	�U��\����[?5����b	�؆̾�_=�f���x=��>X��=��ξX2��N�{_1??qZ��,=���!>��
�X=@�*?i?�Y�<���>Q�#?g3�x����L>F7>��>�%�>��>�Y��k�ڽ?�?E�S?����[���a�>������~���|=�e>ط2�BI�7u[>Lm�<�r���X�:፽C<�<� e?S�>Ɏ�{�}ۡ�W\��������U?/��>�r�>�m?'�"?-�輯��פr�%�(����<"�%?�mp?P>���=
'Ͼ]5���L?m9l?�q]�f��� ��mB��[��B?��?ٽ!?-��=�@��wȳ�� ��_?�/w?9c\������[���`�利>���>M��>L�7�䳻>4�@?N�$���'^��eS6�Ν?�Q@4y�?��z;�%�{��=�?*n�>�P��ž	�������kE=�I�>���qu��[���0�8?�w�?g��>I⁾���U��=�ٕ��Z�?}�?���FFg<U���l��n��~�<�Ϋ=���E"������7���ƾ��
�쪜�3࿼ڥ�>CZ@�U�b*�>D8�X6�TϿ%���[оgSq�y�?5��>��Ƚ����9�j��Pu�L�G�"�H�������>ΰ��d=��8־�G��#0��}j�I??Y���de>��̾�!�e�ľ$���C>�>��>7ʱ>�������+�?'�5�+4�,��Q��(7]?�|�?��d?�)?������v���6-�<0`c?<ˑ?�p?���ξ��/=%�j?�_��tU`��4�sHE��U>�"3?�B�>P�-�~�|=�>���>!g>�#/�v�Ŀ�ٶ�/���Y��?މ�?�o���>n��?ns+?�i�8���[����*���+��<A?�2>���D�!�=0=�NҒ���
?R~0? {�f.���N?���Uݐ��a���1�~�>u�����dl���c�t@��bĤ�ش� ƛ?�3@��?�h����@���X?���>=��G&̾S��==?xy	?p��>x�#��N>� �g���>kp�?��@3%?2���T��ښL>�n�?>E�>���?�8�=�>a��=�R��,�o�8�=)��=
�P�]>�>��f?NU�>~��="�A|-�of�4:������'��"r>�Rn?�Sz?� V>ML���=>����\=6t���� �Y}ۼ�=��>�Щ>�s]>��e�����?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��4a~�)��7�
��=��7?/0�Z�z>���>��=�nv�ͻ��V�s�>�B�?�{�?���>�l?d�o�0�B���1=M�>��k?�s?�o�d���B>��?������L��f?��
@ou@5�^?"C����y�<6[�Q�gqJ��:��{=�Uܽ못-�=����f�;�P!=�6>/>��;>�R8>>��=UN5>$��;��Կ��������k�q�C��#^���a=����蒽 �%�vc�wT��i��e�������f�:�I���V�P<ǖ�=�fu?=�p?��?�??�s<=���>p���>�K��'>f�?��,?�<?�)?���=<س��u�T<��
�о�*1�u?��>�>�>��?�T�>�� �&�^>�ř>��>���=��>(aS��Խ(��>�B�>� ?Z,�>�@<>j>�д��3��;�h�
w�'-̽� �?��� �J��3���H�������Y�=�i.?N�>^��D>п��8H?�	���0�,�+��>��0?�eW?��>����	U�<>4���j��>����ol���)��Q>�q?�n`>K�s>4�7�7���N��!��Cx>f05?�뺾α;���u�C�H���ܾ�8O>��>*��I��������=l�I�=1&9?�?��������sv��:����U>��_>�=2�=p�H>�g��7ƽwYF��t=���=)Y>��"?��#>#>�׵>F^�d��t�?p$�>���>�-�?4�V?�5���Ͼ�*��x�e �>1N?M��>ټ����F��N�=1��>�08>#s��H�ƽs��Y����=��½)qľ��"�����*D\>?�M=z7;�Q�J����<�9s?��������,�3��=�]Q?�
?s�?\q_��"=�:����G����?tp	@C��?�M��~E��/?6q�?/Q�:\ >�*?���>����L%��-?�?�澖�Aփ<�׷?m��?�w�=�Z�������&=JEq?g=�^h�>Tx�~Z�������u��#=.��>�8H?�V��e�O�E>��v
?�?�^�ީ����ȿ8|v����>Z�?���?R�m��A���@����>9��?�gY?Xoi>�g۾l`Z����>ջ@?�R?�>�9���'�k�?�޶?Я�?1J>��?�(s?o��>��u�/7/�O��b^��`nz=
}W;�o�>��>�.���QF����������j����c>��"=��>�t�?���׵=[�������
j����>��n>\H>�n�>�� ?Qx�>T'�>č=���O{���W����J?,֐?�'�\e���<M v=�"[���>f�0?		��eʾǽ�>��U?8|?�2]?�3�>���`��%����S��Wr<z>�v?�O�>�3��3^>q�پ��*���>�}�>h6���q˾h�g���!:L��>i%?���>��L=�!?U�#?�i>]ݯ>��D��,���F���>'��>�c?ߢ~?5�?����/j3����
���O[��L>��y?S�?��>N1��5���Q6��$*7������9�?�e?�t�d�?|k�?�@?�sA?�h>+��O�۾fM��EՂ>��!?g�m�A�O&�m��}?�O?n��>�;����ս
Eּ���v~����?�'\?�>&?^��-a�@�¾7�<j�"�)U�I��;��D���>]�>爈���=�>,Ұ=�Lm��G6�)%g<uw�=A��>Z�=�47�R���t~/?�h���vi�!��=��w�m�M�|ڤ>k�^>����k?�Խ�w�㪿���[���z�?X/�?��?�z���ib�C�:?�r�?�Q	?��>1���YѾ	Ⱦ�Ep�뗍�xG��&�=�f�>�c?������d��<���G��R���U�C����>�̲>��?r�?��C>�}�>�����B2��G��e�b;]��l�Z.�t?&��\���_b�g_~�	�Ǿ j�0�>��8>�>�G?��W>�<]>��>K�<�֌>�;>��h>Ԧ�>`�M>c�;>�}�=>C������)B?H��t9�5P��[ʾ9?��r?��>I��������
��:?�Ϊ?���?,�>�U��\w#�,�!?� �>疳�c'3?c�=iӽ��������ꣾ�2þ� ~�OL{>�b���,=�.�R�5㯾���>�Y?l"*�3pھU)�1����g=p�?��(?��)�eQ���o�U�W��}R���"�g'i�Y���4�$��o�M����3���	��Ju'��^0= �*?	R�?U��!������k��>�"Re>Qz�>IY�>T"�>U�F>68
��2�ڐ]��]&��������>�W{?{Z�>�I?U"<?��P?#vL?��>j��>b}���z�>���;	�>AU�>x�9?I�-?)0?�s?	H+?%hb>+���
���QؾP?c�?�C?t/?��?�ㅾm1ýR����a�ʭy�''��ԫ�=�ɿ<�'׽��s�ɒV=��T>�h?6����8�����/k>�B7?$�>1��>?����������<��>��
?�F�>�����r�������>`��?}��g�=P�)>���=b+���l���=M�ɼj��=qL���0=�[�,<ښ�=�Y�=�X1�7B5:g��:�� ;MH�<�]?���>���>��C>l����:�������>Z��>��>�\�>y�&�ύ�O�����o����>�8�?J�?�|ĽY�}>�7��
����:�T� �����
8=���>�3�>�d?��?��*?s ?��]=ekA������n�������?e!,?P��>u��h�ʾ��ŉ3���?F[?v<a�R���;)�p�¾��Խ
�>�[/�G/~����dD�������(��/��?���?�A��6��x�Կ���[����C?!"�>�X�>��>'�)�\�g�=%�,2;>!��>(R?�#�>��O?Q<{?�[?�hT>��8�1���ә��93���!>�@?��?��?y?�t�>F�>߻)�V�HU��������߂��W=�	Z>8��>�(�>��>I��=��ǽwY���>�kc�=ʋb>I��>��>��>��w>(B�< e>?}h�>w돾���d����ξx���+r?ڢ�?u�+?�Y>b,���R��G�K=�=s�?��?�2??=���ƩD>������K��i��>��>ό�>�S>�F�����>�*?9N�>��6��n��0��隽)�?�2?���<ƈ���xU�W0��X���,B>�eE�>á�\�f��#��]��l�����C���p�� /��f[�Zױ�r#��TB�OǾV]�>�o=l�>��G>Z�%�1V;!�G;ƽ��~>��<���:�+C ��S�9��߽d;�=��=�=�=��=&��Gu?�_?�4:?� M?��>�$d>���2��>�]P���?1B�>-���㞾+i&�4{c��5���W�cuƾ�CM�=ש����=g֨��>%fa>\E{=�e��g�=XhA=���=�7���@L<8�J=v�*=�-�=�@�=g�=M�>�1s?�������zV������6?q�>T��=�&ľ�:?�_>����pܸ�zb��d�?���?��?O��>(S�aK�>�-����ս�n`=Hf��C>\��=�@�&l�>]�8>������������?��@��>?5����Ͽ-%J>��3>�>��R�.�0�ؾX�hc�i\��� ?%�;��k̾�>e=�=O�޾�Nž��1=҈3>�V=����\�*Ŗ=<z�zP7=�w=E�>d�B>��=�+��Uu�=.BO=��=��N>&æ�3�6�ӷ.��H9=��=A�`> �#>8�>�r?��-??�]?~��>�^l�a�Ѿ�ټ�4�>�b�=�s�>�==�j1>m�>�4? :G?jrM?}��>�tj=;��>�W�>B�*�Eo�[[��S�����<y�?�׆?�þ>�y =մM�@>��?��ʽ��?�3?(!?iŏ>pT�ݠ࿭W&�S�.�6����\<7��*=zr�acU� ����q�Ϯ�:�=<w�>n��>Xߟ>�>y>�9>��N>�"�>۩>Qy�<�k�=_���1�<e
����=۪��K��<'�ż����D�+��,�+Ȧ��l�;��;�$_<���;��=���>��> o�>(��= ��mu.>�����0M��W�=w���&B�C d���}�2�.��R7���A>K�X>�>���,��	�?�X>�@>���?$�t?�#>C����Ծ���&�d��!T��=�=*>~�<��6;��_`���M�)�Ҿ���>���>#�>��k>5�+���>�@�s=u�ᾄ�5�14�>�挾������p���������i�$<��0D?�I���|�=�}?��I?�
�?��>������ؾ�0>xU����=�A��r��Ȕ���?��&?w��>�Q�m�D���������j�>�F���U]����z�d��U�=��ξȻ�>��ľb�M
C� ����̓�n�7�6�]��>	J?��?�]ƾ�#���yX�Ѐ��� ��n�>��}?��>W��>]�>��h�zg��r� �5>��g?H'�?�q�?���=m�r=�4�� &�>6�?�ۙ??�?#�h?������>~Ǻٴ!>[���,>Yi >�I=u�>��?��>d��>~�=:)�1;��^پ`2���*=O��=Z;y>�I!>��%>m^=tV�=��=>{^�>H?�>x`�>	�S>���>bk�>�s��y��'�>;s.>���>�6#?ʤ�=�j�!�2�)?��_��ͫI��;3� ��=�O���"����F��=H'�}��>o¿��?�};>�`=�־1?^⾣�e���>�=(�ټky�>��I>�6f>�_>|�>�S�>�h�>���>�JӾv>>��eb!�3+C���R�}�Ѿsz>ԝ��&�����x��O;I��h��]f�7
j�4.��@9=���<�G�?���3�k���)������?�Y�>�6?wҌ����e�>���>�č>rJ������#Ǎ�Nbᾇ�?z��?=5>C��>��<?��>�֎�����\��o��_����f�q#e����b�n��pھ;k���V?��c?��]?E��=���>�b�?����ﾊ�Y>>�@����nz�>c� ?i�J��\C�~����l���y�ۂ>cO�?<�?E�?hb��-9�z2�>ϟW?&Cf?��?�_g?E1?@���?bT>�U�>�?��?��>�>.�>]�<u������=�[����R(�������#��o� =o�+n@=��<��(=��߼�'��PD�g�-�y�I����9�F��uܻ ��<ٰ�>�)\? ��>��>pN4?��&�z�5�ګ�;�/?8�n=��z�~݋��e��������=
mj?)R�? Z?�b>�V?��C� �>`Z�>q�">�nV>�ܯ>����4D�D)�=��>ta>r�=K�G��?���	�����|��<�>>��>��{>\2�� '>�_���z��Fd>f�Q�|���T���G�I�1���u����>��K?w�?ŗ�=���tF���af��n)?�2<?�SM?�	�?jŒ=y?ܾ+�9�G�J��9�K�>Y"�<�B	��������F�:�^ :�Js>3[���㢾I�c>�����ᾋ�n�0>I������O=���D=M���վKB{�_�=��>��¾L[!�������]eJ?�Y�=�I���[_�����>8�>ƃ�>� 5� �u��y@�b��:��=���>у7>�tǼ����:H�3��SX�>S E?�s_?=��?jx��$�s��7C�l>��:��������-?:�>��?H}=>ʌ�=�k���t��d���F��V�>x��>�e���G��Z�����qL$��Q�>�B?� >�?�S?�V?�k`?Y�)?q@?O͎>����O/��?B&?���?��=�Խ��T���8��F� �>�)?̼B�o��>^�?�?+�&?��Q?<�?��>�� �E@����>JZ�>E�W��a���_>�J?V��><Y?�ԃ?�=>��5�!좾թ�iT�=#>��2?Z5#? �?e��>���>L���?
�=П�>�c?�0�?�o?�|�=[�?(=2>,��>2��=z��>*��>�?�WO?n�s?�J?���>��<j5���6��xEs�0�O�*�;M�H<��y=���2t�I�Z��<��;�i���P����K�D���8��;�S�>�ks>ᕾ;1>=žd����@>	��j'�����@�:���=�j�>�?���>%#��i�=���>�C�>8��J(?6�?
?U�;��b�w۾�vK�B�>Y�A?�x�=�l�!��� �u��)g=.�m?�^?�W������%_?�.~?�þ�n.���������˾8�K?��>*�ܾ���>'V�?C�?H�?Z*��ꗇ��9��'~h��������=M��>8�ξ�*���~f>ԒU?A3�>2*�>�o�=fJ���~����'�%?��v?,v�?�ى?�$�=�F�;�ֿ�뾻g���U?�/�>q�44?N.�6ԾmXO��񥾥�˾R���ծ���ׄ��������� �f3z=~O? b?U}?'oZ?H���䁿�k�c�x� �=��������ϨD�q�T�RC���]�Cu�������X�}� >ͼ~���A��=�?N�'?�;0��L�>c�������̾��@><枾��c�=�ۊ���?=�HZ=�ii�װ/�Q����?��>v��>ܿ<?P�[��>��D2���7�p���'Z2>� �>o��> *�>�9-�����ǾӃ���Ͻ�5v>�yc?�K?Z�n?�]�&*1����q�!�D�/��a����B>�>^��>��W�����8&��V>���r�����}��g�	��~=��2?�*�>���>�M�?�?�|	��d���fx� �1����<0�>�i?�@�>��>Kн� ���>(k?C�><��>�ㄾan$���{��ɽ���>��>��>ިe>F5���]�ۡ�������4����=�f?�˄�v�Y�N�>�Q?z��<��8<6r�>����L�#��O�%0"�5�>��?�=�=��;>��Ⱦ����y��ň�MK)?��?�����*��l~>r�!?�H�>"�>o9�?��>�!þI5:D�?g�^?XJ?2A?;�>�=w����[ɽ�g'�+/=3�>4[>�2j=�+�=�����\�ǋ�PRH=�=�Լ�4���n�;�A���Y<��=5>t�ֿ۷9�l�־�+��L��d���+����,�������V��]��cVY�}�7����@K��\9x��2��g�x��f�|��?���?��n�꾁�T��ľxb?����2�ڽJN���gO��e�~�����L�7��T�Jt���F�v�?�4���ǿ���Ѿ��!?��?��w?�
��"��9�� <>1�==غܼ�����˧ʿW۩�3Kf?�Z�>�o���n���/�>�>:id>v�F>��z�������%=J�?�4?˪�>7!{���Ŀ�ȷ��p�<]H�?�@}A?E�(���HV=A��>�	?��?>XS1�I�_����T�>r<�?���?O{M=9�W�-�	��e?�}<��F���ݻ��==�=CM=�����J>�U�>���9TA��?ܽ0�4>�څ>�"�ޫ�΄^�@��<R�]>_�ս�7���ք?�\�jf�>�/��R��zu>�T?�+�>�ՠ=&�,?aMH�wϿX�\��Ea?�6�?;��?��(?�_�>��ܾ�xM?�U6?��>�v&���t����=��伱���D�㾢.V��f�=���>�>&�,�T����O�"ܖ�X��=J�bd���G$�9���f�<^�ϭĽ�P9�i"�n�������E�@�̽<v�=ʫ�=�dN>=�|>�1`>4�B>kSV?�|p?�>u��=b~�(ٍ���;�To=@:���&�����w��l����۾��y�����*���k��ʭC�k`�= �M��唿 O'�J�X�̳<��9%?�">Tپ��R�#p�;�{���(��:C���y��u߾T7�h�`���?��K?� ��� p�q���BE=��_��i?\b���d��$�����=k��:$��<I4>Y�@;��پS�?�:o@�\�/?�8%?�������94>n"��=~�'?N�?t��<�ի>:�*?T��޽JdR>ş4>94�>���>O��=W@���+ �wY?��X?es�������>Q�˾	倾�0=|�>���Y�$���N>f������W���E�(��T=S(W?䛍>U�)���d���C��Q==�x?5�?q3�>}k?��B?��<j��L�S���kw=��W?�'i?�>�|��hо�����5?a�e?��N>�ch���� �.��U�u%?��n?�`?ܘ���v}����g��{m6?)�v?��^�ʚ�������R��G�>� �>���>=9�H�> >?��%���������ܿ3�ﬞ?�@(��?G�<��im�=�"?T��>u�P���ƾ8S������u~e=���>�Ω�yw����*)��8:?<#�?���>���������=ؕ��Z�?;�?����̬f<��Hl��q��Fw�<�Ы=�"��a"�T��R�7�w�ƾ��
�Ǩ���˿���>VY@�L��*�>�:8�^5�8SϿ0��m^оcPq�m�? �>��ȽD�����j��Ou���G�~�H�����L�>Y�>5���ё���{�Ax;�T��.2�>�����>)�S��u���ş���1<�В>���>��>|�������r��?���$οg��������X?�g�?}�?r{?��K<�v���{�x���G?7[s?BZ?O�#���\�}�8�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�rn?�U���T���><�� ���>��E�`|��!�置Y���s陿�n��w��?"@���?�&����9��lK?|�>�f�����t<.=���>��>����l0>%t�<Sa��n>V5�?d�?%/?�*���貿c>7t?`�>�w�?��>>�K ?�+>{'���.8=���=��B>졁���	?�a?} �>A�>�-V�1*'���9�!L@������qJ�e�;>ےf?�sT?HAq>�ׄ��T�;��+��>+��$�u���"P�Yv��}�s�Ԍ?>��+>�=�Y�d(��y�?FY��ܿ�<���%�a;?��);��?�ܾ�&�;��=�Fs?�s>j��mf��� ����\��?�@vx?�����ý8y�>�ӭ>)�z>�*t����<�K=�Cs>z�W?1���
���
Ec��r>-�?ߐ@e�?�<{�K�
?>8��ϒ�K�r�e����}�-x��gL?�ʾ���>!i?_��=�D�����:�r��Q�>�ɳ?W��?,��>��m?'���������=��>DO?�  ?��=UC�Μ�=��>��J�����;��'�z? r@��@AQ?m���P_ѿ���s����?���B�=�o�=m~>F�!����<�Ϳ<�n+����<��>���>�rM>�|s>z/>B*>��>>���W �8ã��|����S�5�"�D7�*琾)��5���3���ľ򫰾�h�Ҁ�n�z�&KT����,l�M�=ŠW?,�R?Z�n?f2?@|���(>TQ��/m0=6��B٘=$J�>�f2?��J?��'?AZ�=n����b������������E��>�/T>��>i��>��>ʈ�R�>>b�D>�3�>��=5�=�h���7=^�T>���>���>�=�>��:>}P>����V����h�d�v�̽�ڢ?9A���J��1���	�������=�=��-?�u>A���:пM���CKH?en����m-�H�>1?GW?	F>��U�S���>q���
j��< >K �/�m�|))��O>ʕ?��f>u>��3�H\8���P��`����|>h-6?�嶾�M9���u���H�^Xݾ�=M>ν�>D/D��r�R�����]pi�*{=u:?�?凳�0̰���u�3;��iR>"\>]�=�f�=�eM>
�b���ƽ�G���.=l��==�^>�d?K,>���=�>�.��0>S���>�C>5�*>hZ@?�t%?,\�����ᄾ�/��.w>��>T�>��>�J�[c�=���>�0b>b���U��d)��qA��AU>��~�	|^��p�y=�◽"��=ծ�=�2��>=�J$=l&�?�����?z��o��xY���,]?c9?6�R=\��%M9�,��������?��@�j�?��پdqM��<?.L�?N�J�_6^>K?���>dh˾�����-?g;�>��ul��"��q�?�O�?�>�ꂄ�(�^��h�=h�?�W
�C֧> }�^��M*��"�U�܋�=��>�LH?�N辁���k�R�X�?*F	?�~��%��XοMPl� �>1D�?�͕?b�q�G؝��!�C?��?��'?��{>�L��'2ڽ(��>�E?@3?���>���������	?ӯ�?,��?��W>�4�?;�w?.�?� �<H+A�����ԅ�9[���;=t��>���=r�ɾ9�R�_���t��DJN�q���I>��<�]�>����E���f�=���~���������>SF�>�dp>gș>��?:N�>�8�>h�Y�0V��$x����!�I?�L�?	紾Ve��Vm<�X�=#E���?(H?���Yo־���>�Z�?	Ul?��g?�
>SM%�9o��"ʿ�o��-o��|�U>��>��>Wơ���=>�[���*�<��>�խ>���=����Κ��-h��~�>�1?+��>��I>�0?Y�!?�|>��>c�(�������F�;��>��>3�?�|?;�%?��]��t,��A���+��QW����=L�`? �?��>�5��8˪�1����<�=�=j�n?��h?DR�����>ZP�?f^G?��`?q�>6x���x�0:a��K�>��!?)��n�A�>(&����?�z?_��>�����Vֽ�-޼b���3��6�?l�[?6&?���6a��¾w��<�o+��?F�Z~<BTT�f{>��>�⇽�ص=�>���=��l��P5�k
u<Cռ=�y�>p!�=�M7�rю���.?=��;Ԛ���G>	 ��)sq���5>���>Od7���?��#>�oV�����(��ޠ��k�?���?�s�?�~:�7^�b�#?P*u?�(?6� ?�ʙ��g����~[�/3���=�.�>���=�w��&���`ݘ�O�����޻��V��>�h�>�G?��?�}�>35�>f��:#��'�1>�*�`��y��0�����B
���ݾ��C�)|���¾Z�:�Fс>/�Z���>�8?��h>�c�>���>����ɓ>@ =>ￚ>i��>�c'>O9�=J:=�w��EԽ�S?t�Ⱦ0&��I辳c��`�D?/�i?�L�>�q�n7����	p?Y��?��?3͈>�d���*��?��>A�����?X�h=��;H1=ƻ�X������`'����>6�½��7�i�K�������?�k?��_�#X˾�;�Ѕ��{o=�M�?��(?_�)���Q��o��W��S�rV�)h��m��	�$�D�p�6돿�]���!��@�(��_*=��*?��?r���)��b%k�`?�sqf>��>7%�>�ܾ>܅I>��	�ٸ1��]�*M'������J�>�W{?��>�;a?�fA?��E?�qJ?6�<>�>y ���.?AF@�#D�>ׄ#?��4??�)? i�>�?#�>>����#-�* ?�A/?�?cj�>���>1о��:�����F/=�V��{����=9a캹�ý"A�L0=�*q>͞?����J8�������n>��7?���>�@�>fZ��fJ���P�<?��>
?E�>o)��K�q�~'����>�)�?����=N�)>9��=����H:@��=!�����=}���֖6�"[+<_��=L�=��F������0]:�BT;Q�<��?��?�>���>����5-��{���58>�9;>�	�>*@�>^�̾�������g�#e�>��??��e���=|��<V�ؾ "о|�S�ھ����*'�>�0?�r7?�?��O?b ?3>y9"��+����L4���!�>w!,?��>�����ʾ��щ3�ܝ?g[?�<a����;)�ڐ¾��Խݱ>�[/�e/~����<D�r���L��5��?�?'A�X�6��x�ڿ���[��x�C?"�>Y�>��>W�)��g�q%��1;>���>jR?($�>.�O?�={?��[?�}T>��8��0��[љ���5���!>�@?���?�?�
y?�h�>e�>��)�v��O�����;�Gゾ"�V=(Z>7��>9�>J�>���=a�ǽ56��E�>�ׁ�=L�b>���>���>���>(}w>��<�=?���>6L��O��`,*���¾d�>zE�?k��?��m?H	;>_�c��D�k>-��K:>�#�?���?��o?����Kg>�;=)`��9:�َ�>ʧ_>%�?�:->�+���
?�`.?���>�����-'���!��Y�;���>��4?�p'�\�Ͽ��u�xU��Κ���<�&y��1g���<�x����D�<�+�����bA��w@��˂��o�������"���3n��?�I�<��ּN^=���<W�<�5�=y"P=�=���=Zv�KkZ=�z���iͼHJ��̗<��=O��<���<�ƾTVu?7aG?tI*?�YM?b�>[#I>?z��K^�>_dV�n�	?�+K>d�Q����7��㡾
����ؾ	Ҿ��b��1��n�=	���>�VB>\��=��%<0`�=�X_=�=�=�xR��b=QC�=p_�=1(�=i��=�� >�=fw?�I��<Ϥ��5O�l�;�79?�K=3�>e����x?�'>�牿"u���w���y?�D�?է�??��l���>u��v��|$'�]�V����<yɐ>pA���N>@<�=ecN�����^�V����?�V
@*�V?U���\����>��7><,>��R�i1��M\�0ib��6Z�Ô!?:E;�H̾��>c��=�%߾͓ƾ�v.=�z6>�8a=�y�DK\��Ù=��z�l�;=�l=\��>�D>��=�믽�#�=�eI=x��=��O>b
��,7��,�~�3=��=��b>��%>8��>_�?1?x�c?�u�>+u��\Ѿ����0�>�:�=�5�>�tS=C�5>C�>�t6?��E?�M?]��>�Ē=?»>�^�>�c*�� n�_5徸Ȧ�Y'�<�?�,�?�>�sb<
#F�����=�5ͽ��?��2?�	?��>���ƿ�AL�m!���< �	>�,�=�<�R��]W�}>ս<Oo=�ƼR��><�>t��>�:�=��>O��<��>P}>�w��$=`�<W�
�8h����=c�<��E=W��=�֙=5_=I. ���ϼ�~��G��<;��=�BC��^>s�>}Ä>U�?�׫=%D��'�x=ۘb�49X����=d(���>���f��|����.��;��ф>�
>��[����G*�>]n�>��>K|�?:}Y?`�I=.)����'��Ę�b���uh��#>��=�d���F���W�O�G����h��>{ߎ>��>|�l>�
,��$?���w=⾼c5���>{������-�C:q��?��^���i��Ѻ�D?F�����=w!~?�I?��?���>� ���ؾ�.0>�H����=���%q�al����?�'?��>��?�D�t@̾�!��Z�>#I�4P�����I�0���	�����> �����о3)3�e��a����B�N,r���>��O?F�?b�;Q���RO�w��͘���l?�g?�+�>�N?*9?�H��ex�@v���e�=�n?.��?f=�?V>$��=�V�����>��?���?Y��?�s?��>���>�n;<>�ߛ���=?e>�[�=k��=yz?� 
?+�
?�'��/�	� �(A�(`�`�=��=�z�>���>`Cq>��=e�h=jݥ=��]>/ў>׏>{�d>s[�>U��>dV��[@���?��#>}8�>a5X?���>9<=��Ν��ƞȽCጾ�>Ͻ���W؝���<S��~��u'��>�q̿��?�^�>�$�K?��!�a�)����>�޿=���=N�>ؚ�=�kp>���>�:�>+#m>N�g> �=�7ﾕ�Z>m�{GX�8���&�aϿ��<�>V=����z����ꁽ�䨽������TO����v�E\����=!��?O������G� �3.F=AM ?��`>�??�Œ��*i�2%>'}?.\�>�g��Y���t������B�k?"�?��P>�K>��Y?��"?(A����m���]��rV�.���b�s4L�P�����}�Q*[?�&l?Μ5?'�>R`�>Y��?iGӾږ�1dm=�}t�M�*��u�>���>��7�H唾1��(#ؾa�T�A{>G1�?��?�\??�׽*� ��+j=_Wo?��T?�̒?�9?�-d?�w	���?���>���>�?��>��?e8�>���=��������<S�g�7Ű����k�1�������Q>��=�f�6���=���<��8������=i;�[�ՠ-<�>J<(�"=c�w===�>�\?��>�F�>ֵ8?&�/�.S9�I��ʉ&?M�D=��|�g����-������tn�=�f?^Ӫ?_�X?�]d>�UC���;�о>n�>��5>�X>?��>�"�WQ��܏=�>%p>�Ʋ=I=_�(�~���
�����<�< �>|��>g��=�����>�1��{�ݽ���>0�O��n̾���(�h��0�������>�JR?�m?:�"�,���z����,_?�?�eE?C2�?Z!p�[����"��;�l
=VX�>t.��VG�u���T����)����@�4>w���K��<On>2�����R�x��WW����v�=��	���<y�
�+�ɾΚl�=h >,>�VϾt��`��ԇ��i�Q?���=� z���W�$Ɲ��8>"+E>_��>����b�n���=��a���ĕ=��>��->����\���[�M��e޾y>�>[QE?0W_?k�?"��As�
�B�����Bc��Oȼ�?_x�>�g?SB>��=�����s�d�yG���>C��>G��D�G��;��S0���$�#��>�9?�>��?O�R?g�
?D�`?�*?1E?�&�>s��d����=&?�y�?�+�=��Խ%^U�k�8�KF����>��)?rIC��_�>xU?h�?A�&?��Q?��?��>�� �%@����>[�>��W��m���S`>f�J?���>nY?{�?�A>>�k5�Bޢ��ʩ�27�=\�>/�2?�;#?J�?�Y�>K��>�>���=��>�]c?_�?�#p?�~�=^?ύ4>u��>LΘ=H�>.��>M�?��N?0�s?V�J?�4�>�܈<U����Z���.p�F�@����;�FH<�wz=�/�H>w�U�����<k��;Z_��]�}�X���r�F��ǌ��}<K��>�g>�Қ�2�*>��ʾ�Li�?Ad>2���V����"��p�d�z�=;�>�c?J��>"^)�6MF=B��>���>��%�_2.?�s?�(?F�W=��e�U边�i��_�>0C?���=�gi�X���>�LX<�6m?CzY?��a�M?����]?��v?���L�S���7���*���J?1�?��Ⱦ-?�>���?4{�?\��>x������79��U�F�o}����+����>�c��	�$�̋">3�>�y�>���=Sh;��Ѿ�d����*�8>g�?^��?�R?�,|>U9|�]r��_���P�O?ϕ�>���F'?ߥ��w律����W���׾���j}��fܗ�#n��d�佗8����	��=�R?�`?�{?܂k?g�$�i��g�}�~�'�C�j�����AC�-[@���I�f�Z�D�$�о����=�}��+A� s�?I�'?=3����>�Y���v�;�8=>,������(��=�x���!K=	
l=Ayh��I0�p ��J�?y�>*��>a3>?on]��?�S�2���7������/>=��>��>�8�>~ث���(�Mgٽ�ƾ���!˽�	w>7�c?�.K?3�m?�b �yY1�F~��� �,�1������JB>��>>�>ʞU�j��L�&�h�>�(Xs��l�-Đ��}	��	�='�2?��>�ƚ>�<�?�?��	�7����vy�
~1�h�B<���>ci?��>u��>$@ս�V!��e�>
�l?�|�>_�>攀������~��N�����>��>�?��>�(齅I\��ѐ�Ï��:?� >�o?-E����Y�@�>L?d�<�=�<+��>QO���� �f�ﾞ�6��Y�=pb?��=MX:>̒ɾf"���w����G)?,M?�����*�AT~>Z'"?2��>:#�>�%�?e
�>>�þ~�q�x�?e�^?�;J?�NA?� �>�-=����CȽ��&���,=my�>��Z>g�m=���=���h\�.����E=�g�=t�μn���<������K<ۦ�<��3>-ݿ�<;�^���5�$�G��!,�Ɠ��즽�����=6�Y����݀�^G�^I�|���v�I�Q���F�S�����?v#�?��=�Ϝ��ݡ�F��}&��K	?�}���x鮾d9���O7��7u����.��d1�~�`�'H�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >^C�<�,����뾭����οA�����^?���>��/��p��>ݥ�>�X>�Hq>����螾{1�<��?7�-?��>Ŏr�1�ɿb����¤<���?0�@}A?��(�S��tV=���>��	?��?>�P1��H������T�>P<�?F��?uM=��W�e�	�Q~e?=x<��F���ݻ��=�=�=0K=����J>�U�>��JWA��Aܽ��4>�ׅ>f�"�J���^���<�]>��ս F��4Մ?2{\��f���/��T��U>��T?+�>�9�=��,?\7H�b}Ͽ�\��*a?�0�?���?*�(?Yۿ��ؚ>w�ܾ��M?YD6?���>�d&��t���=^7�Ȃ������&V�D��=w��>Ņ>��,�݋� �O��K�����=j �Rlƿ��&��%!�S=I`�
���!�Hu�O,��C����`�b����K�==�=�P>>v>fPV>!�,>��Y?��w?�d�>�T�=E� �@/��W���j;;��~���F��z���G��H������I���w�&��)���7=�#l�='�Q�=���� �#�b���F��.?�@$>��ʾZ�M�H�,<Kʾw}��yT��"Ǧ��$̾ڛ1��!n��Ο?h�A?gǅ�x�V����CR��]��g�W?�q����������=/��3s=��>�K�=_���93��IS��t0?�Z?`z��PV��H*>l� �5>=a�+?6�?k�Z<�&�>fI%?��*��_�ob[>Ō3>yޣ>��>�:	>U��'۽R�?��T?�����ڐ>Ps����z�%�`=��>dE5������[>5Ӓ<�茾��U�oD��X:�<��]?���>��$�-#��H���ҽ�b(�#6w?�L.?���=�w~?�m�?/M�>߄�1悿#�H�F�L@?o��?؀�=�}��?�Ǿk���!Z?�br?�Ӄ����t�7�4��@����>���?��?%��=os�� ������r1?��v?�p^��p��1����V�L2�>YP�>���>��9��v�>��>?�#��I�����XU4����?��@���?��:<8�%x�=\5?:^�>3�O��9ƾ2f�������!q=��>w���bv�����D,�b�8?̟�?���>S��������=�ٕ��Z�?��?����,Ag<F���l��n����<xΫ=���G"�1����7���ƾx�
�����g࿼���>>Z@V轜*�>�C8�U6��SϿ,���[о�Sq�d�?'��>7�Ƚ����:�j��Pu�_�G�!�H�����D��>;�>���������H}��9:��ɻ��r�>��ܼ	�>��[�����j쟾^E<E՗>�i�>�>Rt��y4���V�?����!$Ϳ�]��&��5_W?i��?}��?�h#?g�c<��v�;{�{�	���E?�>r?��Y?~�GX�9=N� �j?�]��2U`�*�4�BGE��U>a!3?�C�>��-�_�|=>��>�m>�#/���Ŀ�ٶ�G�����?��?�o���>
��?�r+?�h��7��#[����*��.�P<A?G2>G�����!�A/=��ђ��
?�}0?�|�@/���h?���$���Z�L�Lw���Q�>���Ipb;�""�'G���#q�'���{���?re@��?�����[R��M?�d�>#�{��ي��;�=�=��>�/�>�W�X�i>Z�G�,�:�Z>��?q#�?���>k����ʽ�p��>�+�?(f�>j�?7>���>��>����齌D>d?�<4���v��>�F?��>�my>����I�e�C��ގ�_T�ZD���N>�cq?�ft?��8>.�ʽ�`�=��E�w��Dz��F@�@n���)��ɏ�嶀>�`�>�v�>�����x���?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��S�>i������W勿3�̾�GD��D��t?[����>��>���` ���?��b�G�q�>2�?Q �?��>��?�r���凿��J�>>�w?P�?C >�'��>�s�>e$��G��b8����r?c@(e@I�i?b���e�T���e�Ӿ�鸾��=5M�=mS>�HC��\=}�=�W��;*��Lc+>�W�> x>*��>{�9>��>>'�0>w���ڗ%�҈�������\6��*����A,V�������࿾����xȄ�S�L���i�&��d+�c��=MTw?\�e?�,t?�d?�s½i��=vb�f�?=O��x��=���>_�1?��;?5
?]�D=8z���z�� ��S.��~V��@�>�c>K.�>-?���>6%%�?�>$i>��>��U>DO�=�iw��V ��Y�>(�>�*?���>�><>��>�δ�1��/�h�a�v�U�˽s��?	�����J��2��6?��Z����x�=�`.?W~>a��o=пg��� /H?�����&�y�+��>a�0?RaW?w�>�����T�BJ>3��r�j�Vi>2 �orl���)�$#Q>?h?�[>�{>�z7��89���E����D��>�`/?�¾NZ�+	w�'J�lHԾf\^>Ӟ�>�߁;��#�/���0�x���c�K�<��:?��?F���������^����*O>��X>}��=s��=+/>y�n�0���6-���=k��=E;W>Ҁ?q.,>X"�=��>{6��y,Y� �>��I>X	>k6>?�"?U�:�:�ս�ɐ�Z/��nn>:z�>J�>F�>��T�+��=F��>]7�>����XY�V��t�f�/%1>����kށ�/y��m�M=�dý�u�=��=����2�5�M=�?8���(�������e���^?�1"?K�>&R��lA��r���M�:��?�%@�R�?�d�/\_��!?��?@��Bϩ>�8?~��>����2���uE?�C]��Z���1��=�h̹?�M�?ҿ��]v�;:v�~v=�+?�!�gh�>x�yZ�������u���#=��>�8H?MV����O��>�!w
??�^�橤���ȿ<|v����>]�?���?S�m��A���@�ɂ�>4��?cgY?�oi>�g۾d`Z�{��>��@?�R?��>�9���'�]�?�޶?ѯ�?vI>���?��s?i�>2x�XY/��6��敌���=cwZ;�e�>`_>����(gF�ؓ��h��P�j�\��\�a>;�$=��>�E�4���=�=�싽qH��g�f����>:,q>��I>�Q�>�� ?/b�>ܥ�>�i=�r���ှ�����K?�?][�i�m����<t�=6~`��H?�v3?����
UϾ�x�>l~\?���?�8Z?O~�>�4��|��t����ߴ�p��<*�N>A��>���>�#���uM>�4վ�E��`�>Gd�>���.)ܾ����2Z��'�>w�!?A�>͚�=ϸ*?�	/?�D>	g�>|�O����iN��:�>���>�"?�r�?��+?�P����@��K��a����:�dO�>E�l?�!?>ģ���u����=�W�=�Qq�!y?�#�?	3��j-?���?,c?�S?8�;n����B�轎�>��?�����0L��+���s�ԩ?Z-?0��>m)�S7?����GS#��uݾ�?4Q?2?���q_�¾Xb<D��{�<q�|�ǽW�C>
�>+(��J�=�5�=t3>3hZ��4���=�><b�>Y(�=��$�u0ɽ�U(?kQ̼x����Y>}-��{�t���z>(��>[����?2�>��`��%��z뗿�����l^?��?]*�?�.����P��(?'XV?�Q?�	?U����>�1�ھ�B꾚�侚X>�Z� >Dd�>l@;�Y����� ���R���� ?�X�>��w>�$�>�w?��x>Z�>3����-��
���&���b�����N$��� ����K׾��i���>�g�;�-��U>�>�ꥪ>��
?�Ւ>$�>�G�>ɡ轴Ɩ>a�>[�j>.ƹ>�$C>4�L>r��=K���&,0�{�S?��¾�'�� �0!ƾ�J?R�p?ɑ�>ڧ������P����?�?�?�;�>E?f��D-���?�A�>�ԙ�nv?�؞=���<��w=6�žǌ!�Ll潙�Y� -�>���P*�UK�"��Z��>{K?�J6�F�˾�H�������p=�J�?�+'?�*��VR�#�p�iV���R�,��gi�ǫ���F$��Dp����L������
4)�&;2=W�*?�:�?E��p���Ϩ�_ai��6?�]�g>�=�>�	�>��>|�G>*�	�r3�0�]��i&�Ї��Ġ�>��|?0`�>	�I?�3<?*�P?�lL?"Ύ>�Q�>"���?��>�z�;W!�>Ey�>fl9?'�-?5�/?'?�'+?��b>����s���(پ��?IS?M�?�?=�?[Å��2½�Y��wg��Dz�Ɣ�����=O�<�5ٽ�#u�,X=٪T>G'?����8��n��TKm>+M7?E��>%��>�R���s��{��<��>}0?���>�, ��9r��=�(3�>䛂?cF��{=�(>�H�=������9K�=���O��=�ŏ���9�6��;2�=��=T�&�1���:�gy;�M�<R��>�?���>Z�?�7����C�{[A�_��=�u'���>+�S>4�!���4����KW���d>���?�^�?�D>H�:>�}>�*��$䌾3��������=�k�>?B�>�4?���?|Qa?]�?�S`>��A�(L��Wq�~F����?� ,?=��>����ʾG�6�3�͝?YZ?x<a���z;)�|�¾��Խf�>�Z/�*.~�v��GD�@��P��J�����?6��?�)A�*�6��z������Z��
�C?l"�>#X�>�>�)���g�'$��4;>p��>�R?��>0P?rj{?�[?�U>�;8�����ҙ�)�=� >��??��?�َ?�x?���>�>��)���߾�����}�B��I���^�U=$�X>��>�0�>�g�>�6�=�Ľ�T���J?���=��a>1��>�'�>)��>l�y>ݩ�<s�??���>��q�S�}/��΅�:�(�-7|?�s�?B�?�8-��=@�89���W��>�θ?p��?ȋC?u�� �$>�U��{����/��g>����?p��>"֌=��6?saH?Ľ>�+0�fD��ކ��a[��/;?=�M?�^��ſ�Eq�6�o�8R����G<�œ�\If�:���[�y��=ט�F� ����[��g���ד���������|��O�>~��=���=�
�=�@�</pǼD�<S|L=A��<j�=�4r�f�n<q[8�,x��o���5X\���H<s�C=��ӻB㋾�hY?�[M?�=?2�A?�b�>�>rM���^�>�mɻ ?�w�>!!!=�)o��$r�crǾ�Ӓ�ظ������k_�Iþn��=84�x~�=C�F>?5>��T=���=�Q�=���=Y̒�M�I=���=��=�D&=�R�=@�>K��=-�n?&��e(���
{�
<��,?@HA�X�>��!A?wuM=�j��@hο����?P��?���?/��>�R��'��>U��?�����=��ɽb�c>4�>�����#�>��=G��=���q�n��E�?b��?�k?5��"�6#�>�'7>$/>?�R��1��Z�
�`�r�W�bF!?�f;��̾���>�7�="�޾��ž�/=�6>�X=a���\��=�}�l�;=�mh=l��>��D>�d�=JA�����=1�E=�V�=^O>㜗�2��&���7=JR�=�eb>��$>���>6�	?��,?w\?O�>-�`�KҾ���� �>���<:�>�X(:�)>ۨ�>o!D?8JX?��B?��>���=!
�>��>��(�P�{�>ƾ{	��{��<�h�?��?�F�>ڑ�<�r>������6�'�׽�a?�2?Iv
?wz>��@�g�P��7��������=��>8���s�3����=p���oy<����=j�>e��>�˰>�e>B�6>k(>^��>�R>δ�=�;~�`3z��F�����g�=�u �.�=M��=���=Q6X�n(���ܖ�Jr
�ۄ*�5�=H{��>T0�>7>%#�>�c =�����>�=��d��Q��(>b���<��.a�u�(s��<�&Mr>a��>m�2������
?g�=> {d>p�?Yt?���=�`q�+!��.���[6���{���<k=j%��!���K�>;��=��%��>pԎ>��>]�l>e,�E'?���v=(�ᾰ\5��'�>�P����mi��3q��,�����h�=�����D?�C��|��=~?��I?0�?|��>������ؾ8�/>T�����=��.Yq��ړ��?�'?͕�>���E�D�j ھ)���A�>��U�2��ؐ�=\^�� �=��A�>0�������[�*�����9�)O>������>�8t?�`�?m2���>��]C��踾e!U=O�>���?Џ>�Y�>���>�Y��������]�>�?��?vs�?t�>���=3����>5S	?J��?��?�^s?�@�?��>?��;�� >.s���m�=X�>���=_��=Y<?�g
?6~
?�*����	�K����"^��<M'�=�F�>I2�>�r>���=Hre=H��=e\>���>)Q�>)Nd>k�>~`�>`w���k��y��>�[�=�Zz>Y�@?KK�>���8�w���m3Ƚ�萾�H���s$�\��=ֽ&�S��r<��2�>��ƿ,,�?-��>
�-�8�>�)$�n�W���p>�\O>Wn=?�>��4=Sڢ=��>�E�>Ӝ�>�_�>�XE>�7�g&>�����;2��H��\b�sK�l�>/ة��������0ʽs�/�/ַ��.���u�`��b�L�e�&=Y��?��<��X�I���߶=�K?xM@>p�-?�ʆ��'�=��=�j�>�P>[�)��폿�Q|�7���? �?��g>�+c>�SF?R�&?��Ѿ�5�q�P�Z�q��30��r��_�N�����w�������=��?�wT?�%(?���=�?�>�i?l������=I�4����@D9>�J?ȣƾ�~˾!�ݾh���7A.��[�>���?	*d?��?u����6���3>��a?�iZ?�L�?pU?��8?�k"�-�?���>�
?P)?��>)!�>ue�=t�L����=͹i��B<�
�p����*ѽd�����<�9�=���=���<�+����=��1���έR���h<�k==�d�;�4=��=[�=ö�>�]?��>+͉>R�5?����7�签�,?x�<=(r��*Ջ�ǥ��W��*>E�i?v(�?�?[?d�c>ZlC���;�1*>�X�>Ȥ&>��W>Hx�>�% �;�H�F��=�9>��>�ѣ=�\�澂�7��y)���	�<�k!>���>6�d>����>�������>��e��m���N�X�f�em'�?�����>�wP?�X?�|ټ߱̾�Kͻ/��Az>?%?34?'Е?�������ND�;��%����x>a�w#��q���+��f�
�������=�j���㢾I�c>�����ᾋ�n�0>I������O=���D=M���վKB{�_�=��>��¾L[!�������]eJ?�Y�=�I���[_�����>8�>ƃ�>� 5� �u��y@�b��:��=���>у7>�tǼ����:H�3��SX�>S E?�s_?=��?jx��$�s��7C�l>��:��������-?:�>��?H}=>ʌ�=�k���t��d���F��V�>x��>�e���G��Z�����qL$��Q�>�B?� >�?�S?�V?�k`?Y�)?q@?O͎>����O/��?B&?���?��=�Խ��T���8��F� �>�)?̼B�o��>^�?�?+�&?��Q?<�?��>�� �E@����>JZ�>E�W��a���_>�J?V��><Y?�ԃ?�=>��5�!좾թ�iT�=#>��2?Z5#? �?e��>���>L���?
�=П�>�c?�0�?�o?�|�=[�?(=2>,��>2��=z��>*��>�?�WO?n�s?�J?���>��<j5���6��xEs�0�O�*�;M�H<��y=���2t�I�Z��<��;�i���P����K�D���8��;�S�>�ks>ᕾ;1>=žd����@>	��j'�����@�:���=�j�>�?���>%#��i�=���>�C�>8��J(?6�?
?U�;��b�w۾�vK�B�>Y�A?�x�=�l�!��� �u��)g=.�m?�^?�W������%_?�.~?�þ�n.���������˾8�K?��>*�ܾ���>'V�?C�?H�?Z*��ꗇ��9��'~h��������=M��>8�ξ�*���~f>ԒU?A3�>2*�>�o�=fJ���~����'�%?��v?,v�?�ى?�$�=�F�;�ֿ�뾻g���U?�/�>q�44?N.�6ԾmXO��񥾥�˾R���ծ���ׄ��������� �f3z=~O? b?U}?'oZ?H���䁿�k�c�x� �=��������ϨD�q�T�RC���]�Cu�������X�}� >ͼ~���A��=�?N�'?�;0��L�>c�������̾��@><枾��c�=�ۊ���?=�HZ=�ii�װ/�Q����?��>v��>ܿ<?P�[��>��D2���7�p���'Z2>� �>o��> *�>�9-�����ǾӃ���Ͻ�5v>�yc?�K?Z�n?�]�&*1����q�!�D�/��a����B>�>^��>��W�����8&��V>���r�����}��g�	��~=��2?�*�>���>�M�?�?�|	��d���fx� �1����<0�>�i?�@�>��>Kн� ���>(k?C�><��>�ㄾan$���{��ɽ���>��>��>ިe>F5���]�ۡ�������4����=�f?�˄�v�Y�N�>�Q?z��<��8<6r�>����L�#��O�%0"�5�>��?�=�=��;>��Ⱦ����y��ň�MK)?��?�����*��l~>r�!?�H�>"�>o9�?��>�!þI5:D�?g�^?XJ?2A?;�>�=w����[ɽ�g'�+/=3�>4[>�2j=�+�=�����\�ǋ�PRH=�=�Լ�4���n�;�A���Y<��=5>t�ֿ۷9�l�־�+��L��d���+����,�������V��]��cVY�}�7����@K��\9x��2��g�x��f�|��?���?��n�꾁�T��ľxb?����2�ڽJN���gO��e�~�����L�7��T�Jt���F�v�?�4���ǿ���Ѿ��!?��?��w?�
��"��9�� <>1�==غܼ�����˧ʿW۩�3Kf?�Z�>�o���n���/�>�>:id>v�F>��z�������%=J�?�4?˪�>7!{���Ŀ�ȷ��p�<]H�?�@}A?E�(���HV=A��>�	?��?>XS1�I�_����T�>r<�?���?O{M=9�W�-�	��e?�}<��F���ݻ��==�=CM=�����J>�U�>���9TA��?ܽ0�4>�څ>�"�ޫ�΄^�@��<R�]>_�ս�7���ք?�\�jf�>�/��R��zu>�T?�+�>�ՠ=&�,?aMH�wϿX�\��Ea?�6�?;��?��(?�_�>��ܾ�xM?�U6?��>�v&���t����=��伱���D�㾢.V��f�=���>�>&�,�T����O�"ܖ�X��=J�bd���G$�9���f�<^�ϭĽ�P9�i"�n�������E�@�̽<v�=ʫ�=�dN>=�|>�1`>4�B>kSV?�|p?�>u��=b~�(ٍ���;�To=@:���&�����w��l����۾��y�����*���k��ʭC�k`�= �M��唿 O'�J�X�̳<��9%?�">Tپ��R�#p�;�{���(��:C���y��u߾T7�h�`���?��K?� ��� p�q���BE=��_��i?\b���d��$�����=k��:$��<I4>Y�@;��پS�?�:o@�\�/?�8%?�������94>n"��=~�'?N�?t��<�ի>:�*?T��޽JdR>ş4>94�>���>O��=W@���+ �wY?��X?es�������>Q�˾	倾�0=|�>���Y�$���N>f������W���E�(��T=S(W?䛍>U�)���d���C��Q==�x?5�?q3�>}k?��B?��<j��L�S���kw=��W?�'i?�>�|��hо�����5?a�e?��N>�ch���� �.��U�u%?��n?�`?ܘ���v}����g��{m6?)�v?��^�ʚ�������R��G�>� �>���>=9�H�> >?��%���������ܿ3�ﬞ?�@(��?G�<��im�=�"?T��>u�P���ƾ8S������u~e=���>�Ω�yw����*)��8:?<#�?���>���������=ؕ��Z�?;�?����̬f<��Hl��q��Fw�<�Ы=�"��a"�T��R�7�w�ƾ��
�Ǩ���˿���>VY@�L��*�>�:8�^5�8SϿ0��m^оcPq�m�? �>��ȽD�����j��Ou���G�~�H�����L�>Y�>5���ё���{�Ax;�T��.2�>�����>)�S��u���ş���1<�В>���>��>|�������r��?���$οg��������X?�g�?}�?r{?��K<�v���{�x���G?7[s?BZ?O�#���\�}�8�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�rn?�U���T���><�� ���>��E�`|��!�置Y���s陿�n��w��?"@���?�&����9��lK?|�>�f�����t<.=���>��>����l0>%t�<Sa��n>V5�?d�?%/?�*���貿c>7t?`�>�w�?��>>�K ?�+>{'���.8=���=��B>졁���	?�a?} �>A�>�-V�1*'���9�!L@������qJ�e�;>ےf?�sT?HAq>�ׄ��T�;��+��>+��$�u���"P�Yv��}�s�Ԍ?>��+>�=�Y�d(��y�?FY��ܿ�<���%�a;?��);��?�ܾ�&�;��=�Fs?�s>j��mf��� ����\��?�@vx?�����ý8y�>�ӭ>)�z>�*t����<�K=�Cs>z�W?1���
���
Ec��r>-�?ߐ@e�?�<{�K�
?>8��ϒ�K�r�e����}�-x��gL?�ʾ���>!i?_��=�D�����:�r��Q�>�ɳ?W��?,��>��m?'���������=��>DO?�  ?��=UC�Μ�=��>��J�����;��'�z? r@��@AQ?m���P_ѿ���s����?���B�=�o�=m~>F�!����<�Ϳ<�n+����<��>���>�rM>�|s>z/>B*>��>>���W �8ã��|����S�5�"�D7�*琾)��5���3���ľ򫰾�h�Ҁ�n�z�&KT����,l�M�=ŠW?,�R?Z�n?f2?@|���(>TQ��/m0=6��B٘=$J�>�f2?��J?��'?AZ�=n����b������������E��>�/T>��>i��>��>ʈ�R�>>b�D>�3�>��=5�=�h���7=^�T>���>���>�=�>��:>}P>����V����h�d�v�̽�ڢ?9A���J��1���	�������=�=��-?�u>A���:пM���CKH?en����m-�H�>1?GW?	F>��U�S���>q���
j��< >K �/�m�|))��O>ʕ?��f>u>��3�H\8���P��`����|>h-6?�嶾�M9���u���H�^Xݾ�=M>ν�>D/D��r�R�����]pi�*{=u:?�?凳�0̰���u�3;��iR>"\>]�=�f�=�eM>
�b���ƽ�G���.=l��==�^>�d?K,>���=�>�.��0>S���>�C>5�*>hZ@?�t%?,\�����ᄾ�/��.w>��>T�>��>�J�[c�=���>�0b>b���U��d)��qA��AU>��~�	|^��p�y=�◽"��=ծ�=�2��>=�J$=l&�?�����?z��o��xY���,]?c9?6�R=\��%M9�,��������?��@�j�?��پdqM��<?.L�?N�J�_6^>K?���>dh˾�����-?g;�>��ul��"��q�?�O�?�>�ꂄ�(�^��h�=h�?�W
�C֧> }�^��M*��"�U�܋�=��>�LH?�N辁���k�R�X�?*F	?�~��%��XοMPl� �>1D�?�͕?b�q�G؝��!�C?��?��'?��{>�L��'2ڽ(��>�E?@3?���>���������	?ӯ�?,��?��W>�4�?;�w?.�?� �<H+A�����ԅ�9[���;=t��>���=r�ɾ9�R�_���t��DJN�q���I>��<�]�>����E���f�=���~���������>SF�>�dp>gș>��?:N�>�8�>h�Y�0V��$x����!�I?�L�?	紾Ve��Vm<�X�=#E���?(H?���Yo־���>�Z�?	Ul?��g?�
>SM%�9o��"ʿ�o��-o��|�U>��>��>Wơ���=>�[���*�<��>�խ>���=����Κ��-h��~�>�1?+��>��I>�0?Y�!?�|>��>c�(�������F�;��>��>3�?�|?;�%?��]��t,��A���+��QW����=L�`? �?��>�5��8˪�1����<�=�=j�n?��h?DR�����>ZP�?f^G?��`?q�>6x���x�0:a��K�>��!?)��n�A�>(&����?�z?_��>�����Vֽ�-޼b���3��6�?l�[?6&?���6a��¾w��<�o+��?F�Z~<BTT�f{>��>�⇽�ص=�>���=��l��P5�k
u<Cռ=�y�>p!�=�M7�rю���.?=��;Ԛ���G>	 ��)sq���5>���>Od7���?��#>�oV�����(��ޠ��k�?���?�s�?�~:�7^�b�#?P*u?�(?6� ?�ʙ��g����~[�/3���=�.�>���=�w��&���`ݘ�O�����޻��V��>�h�>�G?��?�}�>35�>f��:#��'�1>�*�`��y��0�����B
���ݾ��C�)|���¾Z�:�Fс>/�Z���>�8?��h>�c�>���>����ɓ>@ =>ￚ>i��>�c'>O9�=J:=�w��EԽ�S?t�Ⱦ0&��I辳c��`�D?/�i?�L�>�q�n7����	p?Y��?��?3͈>�d���*��?��>A�����?X�h=��;H1=ƻ�X������`'����>6�½��7�i�K�������?�k?��_�#X˾�;�Ѕ��{o=�M�?��(?_�)���Q��o��W��S�rV�)h��m��	�$�D�p�6돿�]���!��@�(��_*=��*?��?r���)��b%k�`?�sqf>��>7%�>�ܾ>܅I>��	�ٸ1��]�*M'������J�>�W{?��>�;a?�fA?��E?�qJ?6�<>�>y ���.?AF@�#D�>ׄ#?��4??�)? i�>�?#�>>����#-�* ?�A/?�?cj�>���>1о��:�����F/=�V��{����=9a캹�ý"A�L0=�*q>͞?����J8�������n>��7?���>�@�>fZ��fJ���P�<?��>
?E�>o)��K�q�~'����>�)�?����=N�)>9��=����H:@��=!�����=}���֖6�"[+<_��=L�=��F������0]:�BT;Q�<��?��?�>���>����5-��{���58>�9;>�	�>*@�>^�̾�������g�#e�>��??��e���=|��<V�ؾ "о|�S�ھ����*'�>�0?�r7?�?��O?b ?3>y9"��+����L4���!�>w!,?��>�����ʾ��щ3�ܝ?g[?�<a����;)�ڐ¾��Խݱ>�[/�e/~����<D�r���L��5��?�?'A�X�6��x�ڿ���[��x�C?"�>Y�>��>W�)��g�q%��1;>���>jR?($�>.�O?�={?��[?�}T>��8��0��[љ���5���!>�@?���?�?�
y?�h�>e�>��)�v��O�����;�Gゾ"�V=(Z>7��>9�>J�>���=a�ǽ56��E�>�ׁ�=L�b>���>���>���>(}w>��<�=?���>6L��O��`,*���¾d�>zE�?k��?��m?H	;>_�c��D�k>-��K:>�#�?���?��o?����Kg>�;=)`��9:�َ�>ʧ_>%�?�:->�+���
?�`.?���>�����-'���!��Y�;���>��4?�p'�\�Ͽ��u�xU��Κ���<�&y��1g���<�x����D�<�+�����bA��w@��˂��o�������"���3n��?�I�<��ּN^=���<W�<�5�=y"P=�=���=Zv�KkZ=�z���iͼHJ��̗<��=O��<���<�ƾTVu?7aG?tI*?�YM?b�>[#I>?z��K^�>_dV�n�	?�+K>d�Q����7��㡾
����ؾ	Ҿ��b��1��n�=	���>�VB>\��=��%<0`�=�X_=�=�=�xR��b=QC�=p_�=1(�=i��=�� >�=fw?�I��<Ϥ��5O�l�;�79?�K=3�>e����x?�'>�牿"u���w���y?�D�?է�??��l���>u��v��|$'�]�V����<yɐ>pA���N>@<�=ecN�����^�V����?�V
@*�V?U���\����>��7><,>��R�i1��M\�0ib��6Z�Ô!?:E;�H̾��>c��=�%߾͓ƾ�v.=�z6>�8a=�y�DK\��Ù=��z�l�;=�l=\��>�D>��=�믽�#�=�eI=x��=��O>b
��,7��,�~�3=��=��b>��%>8��>_�?1?x�c?�u�>+u��\Ѿ����0�>�:�=�5�>�tS=C�5>C�>�t6?��E?�M?]��>�Ē=?»>�^�>�c*�� n�_5徸Ȧ�Y'�<�?�,�?�>�sb<
#F�����=�5ͽ��?��2?�	?��>���ƿ�AL�m!���< �	>�,�=�<�R��]W�}>ս<Oo=�ƼR��><�>t��>�:�=��>O��<��>P}>�w��$=`�<W�
�8h����=c�<��E=W��=�֙=5_=I. ���ϼ�~��G��<;��=�BC��^>s�>}Ä>U�?�׫=%D��'�x=ۘb�49X����=d(���>���f��|����.��;��ф>�
>��[����G*�>]n�>��>K|�?:}Y?`�I=.)����'��Ę�b���uh��#>��=�d���F���W�O�G����h��>{ߎ>��>|�l>�
,��$?���w=⾼c5���>{������-�C:q��?��^���i��Ѻ�D?F�����=w!~?�I?��?���>� ���ؾ�.0>�H����=���%q�al����?�'?��>��?�D�t@̾�!��Z�>#I�4P�����I�0���	�����> �����о3)3�e��a����B�N,r���>��O?F�?b�;Q���RO�w��͘���l?�g?�+�>�N?*9?�H��ex�@v���e�=�n?.��?f=�?V>$��=�V�����>��?���?Y��?�s?��>���>�n;<>�ߛ���=?e>�[�=k��=yz?� 
?+�
?�'��/�	� �(A�(`�`�=��=�z�>���>`Cq>��=e�h=jݥ=��]>/ў>׏>{�d>s[�>U��>dV��[@���?��#>}8�>a5X?���>9<=��Ν��ƞȽCጾ�>Ͻ���W؝���<S��~��u'��>�q̿��?�^�>�$�K?��!�a�)����>�޿=���=N�>ؚ�=�kp>���>�:�>+#m>N�g> �=�7ﾕ�Z>m�{GX�8���&�aϿ��<�>V=����z����ꁽ�䨽������TO����v�E\����=!��?O������G� �3.F=AM ?��`>�??�Œ��*i�2%>'}?.\�>�g��Y���t������B�k?"�?��P>�K>��Y?��"?(A����m���]��rV�.���b�s4L�P�����}�Q*[?�&l?Μ5?'�>R`�>Y��?iGӾږ�1dm=�}t�M�*��u�>���>��7�H唾1��(#ؾa�T�A{>G1�?��?�\??�׽*� ��+j=_Wo?��T?�̒?�9?�-d?�w	���?���>���>�?��>��?e8�>���=��������<S�g�7Ű����k�1�������Q>��=�f�6���=���<��8������=i;�[�ՠ-<�>J<(�"=c�w===�>�\?��>�F�>ֵ8?&�/�.S9�I��ʉ&?M�D=��|�g����-������tn�=�f?^Ӫ?_�X?�]d>�UC���;�о>n�>��5>�X>?��>�"�WQ��܏=�>%p>�Ʋ=I=_�(�~���
�����<�< �>|��>g��=�����>�1��{�ݽ���>0�O��n̾���(�h��0�������>�JR?�m?:�"�,���z����,_?�?�eE?C2�?Z!p�[����"��;�l
=VX�>t.��VG�u���T����)����@�4>w���ˠ�jb>l��fz޾"�n���I����UN=�u��U=��v�վ��~����=�C
>����� ����٪�'J?Suj=�l���dU�W�����>EŘ>��>_:��<w�xy@�����8�=)��>�M;>������nG��)�p|�>��E?V�]?�̄?:����^s�|WB�����C&��c�G�[D?���>�	?�:>��=����^���d�fE��^�>�J�>*��~J�����<��q�$���>/?A�>P�? R?K7?��a?��)?P3?f�>H���]����X&?.��?�|�=S�ݽ�X���7��)F���>��)?�B��ɓ>�?� ?�5'?�Q?N\?I>�0��A���>�?�>g�V��Q��,�[>�gI?9��>�9X?Tу?�9?>6k5�q����歽���=1�(>��2?]	"?^\?�*�>Q��>���Z��>b�>�n�?@�x?1�z?�wؼ 7>�R�>���>��>�U�>���>75�>%�'?��\?�6S?�u�>�3N=��S�K�]�ɤ�<�C�=�mTM<�hM�$��=�����=�L�;��(������Ͻ�RJ�]u���=Gg�>��s>��`�0>\žs(��~�@>�ˤ��O��*犾\�:���=*z�>)�?��>�5#��c�=ӝ�>NJ�>����G(?�??��';��b�A۾��K����>�B?�0�=t�l�K����v��/f=��m?W�^?a�W�2����V?�tn?��ƾ�S!���Ͼ�Q�hK��`O?�?W���?>���?Ĺ�?���>I��&Jv�H����i�yӾ�,�=ú�>��k�����=Qo??=�>�f�>t�>�	��3���o����?S�?-��?@E�?� ��>D��ֿ�]Ѿ~{��9(6?vG�>v����7? ��<i|�2:��ݰ�s�v୾W��yp���f�4�
�x̾��~�M��=~I�>峃?��~?Q�H?ж �M0}�'�[�tQ��ܲI��E��=K�?�K��4P���\�1	��������;�L,�9�K>��~��A�х�?[�'?//����>�J��e��[F;��B>�~�����=�l��R�@= p[=~<h��8.�r ��6 ?��>5u�>%�<?Q�[�t>���1���7�.?����4>6��>+��>��>(��:�-�B���ɾ���N�ѽe�u>�Yc?��K?9�n?W� �w1��T��ݙ!��^,����X`C>\4>z�>��W�~�/�%��,>���r�G��֔���	�Oc�=�2?+�>�n�>^�?�?~�	������&x��%1�䚃<B��>�'i?ؠ�>I�>eMѽ�� �I��>p�l?��>�I?@x&�cR1�r�i�9�ʽ�T?�y�>�*?p�>�M��?�h��%��*���B�2#&>�Y�?�g�񉾮J>�OY?nJc=Q�"���?4��: 4����8�=���>�z?�=���=菵��������Nz��D(?�p?:���ZJ)��E~>C�?w��>p��>Z��?�Ρ>sÿ��)��^?�e[?�7F?�NA?<�>��=��ӽ}�ʽ�+��?-=죇>�d>��=={��=Hs"�W�5�%���}=l��=�i��"Խ�]E�;�,��:=��=X5>ҋ�]�L�~��R��4Eھ�\�7K��Ƒ񻈣,�(��48ʾpE���`�!�ͽ��<��X�����.��n�����?t��?8{/�u����#���̃�W��-#?�@ ������ξ�OU�>���Siʾ�a��'���P����u���?�~w��vͿ뗿5��,��>�/*?���?{! � �*�֣'��e�=m5"=��%���������Ͽ����b?:��>���h�����>*\^>	�2>l�X>cu��'վ���>Z?Y(?�Y�>}ߊ�l�ǿ M����=v�?DZ@KrA?��(��O�t�U=�%�>��	?H3@>�y1��\�����n0�>hA�?��?�QN=�W�'�	��ue?`�<k�F��
ۻ��=�1�=�=���A�J>B+�>6����A�a۽�~4>��>�"�(��.w^�<}p]>4�սѯ���Մ?�|\�`f�Ԩ/�JV��oi>��T?8&�>�&�=�,?�;H��|Ͽ�\��1a?P1�?��?Q�(?�ۿ���>��ܾA�M?'D6?���>Ag&�5�t����=���$��t��*#V���=���>�v>��,������O��^��i��=����ƿ#�T���$�<@Ɓ�?F���[�ʂ���N���g����W��Rҽ
�=��=��Z>*�>�k>8�U>a;`?>�o?�`|>� >�.½���ddپhɏ=����� ��z���������YMྟ,ξr��`q�������D��ێ=��]�	\��N*��i��F��A<?J�5>���R���0��ž�ѝ�� <��ڽU�ľ��=��v�+��?DcU?Z{��(�E�}"�&_߽�&���t?��[���_�����a=�]��*w�<��>��=w�mT>��K��0?C?{����C���P+>x���_=��*?��?�#�<��>�L$?*�=p�D>X>s�6>�s�>���>�W>X̮� ���?6�T?����ޝ����>>g���\y�fHU=R
>�=1�����>X>�l<Tt��5�)���E��<(W?���>�)� �Pa��D��H==ֱx?�?�.�>�zk?�B?Lˤ<�h����S���lew=a�W?k*i?��>\����	о+���^�5?H�e?>�N>`h�N���.��T��%?��n?T_?z{���v}�~������n6?C�x?0�b���c��/?�mt�>���>���>N�;���>fjD?���y���,���E.�g�?�0@O��?��;�9���f=p�>Z�>�?)���ǾM��1�ƾE�G=P�>�i���k{�P�b��u0=?{�?	I�>�V�����}�=����:�?	�?�����o<��Z)l�H������<���=����#&��.���7�1�ƾ�
�D朾�F��K��>�T@h����>��8�U3��EϿ���\`оq�p�c�?��>�ɽ)ԣ���j�Du��eG�8�H�+C���M�>��>���o���H�{��q;��$����>2��	�>y�S��&��������5<��>���>��>[,��%轾8ř?dc��@οI�����N�X?5h�?�n�?�p?~�9<��v�(�{����2.G?��s?QZ?r%��=]���7��j?g_���U`�Ȏ4�~HE��U>�"3?�C�>z�-�l�|=�>;��>+g>�#/�m�Ŀ�ٶ�e���<��?��?qo꾔��>���?9s+?�i��7��v\����*�ά*��<A?�2>����U�!�20=�5Ғ�Ƽ
?�~0?ay�=.�khw?����̀�3^]�����\�>��K��.뽄�8��F����|��褿v���}��?��@���?Z�ν3�@�_�D?��>m��c?����TYb�q��>j�*>�X8����>��A���l�+����Q�?^q @�F?%l���.��U��=+?�r�>��?��=o.�>՟�=����y�;�ʯ">�=Y6��g?~N?`:�>d+�=6�<���.���E��Q�@���C��j�>rTa?��L?.7`>*^��v/�b� �P(Ͻ	/���ҼPD?��`-�g@�V$4>�D<>`�>,3G�AӾl�?��ِ׿e1���I`��	?�w[>(c?���l�W�9�a=s�M? R�>d;�+������d6��e�?J#�? ?�9�E�=.��=�>�b�>�mm�ۉ�a�#���J>��7?G�Ž���ke��K�>E��?� @��?w�c�fu?���<����S���K��ܴ��؞:��w?w-�_QK>:�?xj�=���5ʟ���S�v\�>���?�>�?��?b)�?L߈�j�'�	���?�&�?1�>�C)�h�޾({�=#?����w����Ѿ�uj?{3@�J@��Z?�Z��¾߿�T����������п=���=OK>2J ��U�=���=���<J"�<��>��>���>��>A�v>�VD>�t�=�!��H#��4��ᷚ���4��;����'V�%B���<���_��k���(��dXV����t������罊��Nb�=w�X?�P?��j?M��>�����\>�����t=�h����=:�>d0?3\I?�+'?�= 䚾�b�_������)���Oc�>�H>�V�>��>u�>-Q;�hE>�2>���>��>Z��<�ѕ�u�%<cMX>�`�>o��>� �>�]	>�,>Ϲ��ު���e�ˎ���y��Z�?�Ԝ�md\�\j��3����=���=U)??U�=����mӿ˭�tcT?ĚZ� /-�Ǐ�Y�=�:?'�m?��>�O������YW>��[#G��@�=>)��ە�Ht9�Ӷ:>��(?�_>��R>n�2�Ck2�w�N�����y�>��-?�˶}�c+o��A�0Q޾M_S>�F�>Kͪ:��������~��<^��U=n9??t5?����!����}�5����HW>(�P>���<'|�=;f(>ʽ٥���R����<�m�=�{�>��?$�1>G��=uǤ>_��h�T��J�> a@>�3>b!@?#h%?n%	��"������-2�X�w>���>g�~>{�>�VI���=�w�>�e>�#��x����
��B���U>��}�w�Z�aCj��v=Sڜ��f�=��=�y��*?;�^'=�]�?�L��)����.���ľ�h?���>/ʗ<�k����d�Q븿�/����?�B@��?m��*�Z���?�͝?�[��z�>Ӷ
?3�>������)U?$g��rĽڕ����R����?܎�?F�_��ǁ�5�c��>o,?@���/�>U��e�������u�W�=���>�gH?����sO��G=�/X
?�?>r����ɿ+wv����>��?��?��m�a��@�?�>0��?=�X?�1i>��ھM�Y�9��>�@?�Q?c�>!��'��&?��?���?G�;>�p�?5%X?Κ?��1�@A�e*���.}�-�>T�.> C�>P�|>����\�H����)��\dI������>�{�=b{�>P9��ž��=<���W%��L�E�(��>�>R�=���>?�?��>�de>I0Ͻ�Jq������ɾ�/<?�]�?2	��w�a��<���d�B��
\?N?=)�>���`	�=�de?Mv?��k?�C>�<��_����ʦ��=���>��>���>�sD�8S>�G����V={�>L��>�5&��G�T�����⽺C�>g ?F��>I> �? )?�|b>�U�>UI:�����B���>�(�>P�?(|?��?����w4�Z���sѤ���Q���>0Tn?I�?E�>�����-�����;�ƹ�ý�n�?�G\?s���A�>#_�?��E?o]K?eqp>8�����z�ý"�'>�p?�Y#�H�@��� �܃���?�7?�W�>I���j�7�	����
����c?��[?VO$? ��?�b�:Ѿ�<g���	*={�<��R���>_�>��y����=A>ʘ�=��\�׹J�����Q@�=�T�>�H�=�1�y�.=,?ʾG�{ۃ���=��r�?xD�~�>�IL>����^?pl=��{�����x��,	U�� �?���?Zk�?Q��>�h��$=?�?S	?p"�>�J���}޾/�ྱPw�~x��w�`�>���>��l���I���י���F��X�Ž�C�۾�>�B>�&�>�?I��>F\�>$�о��8��X�I��Y�:�>#���'��Z��쾅S��v�d�V��������U>�߭=+G�>��?2ۗ> �>=��>��&�%��>8^>�|�>�{�>���>Ã�>��)>��|5��KR?V����'��辡����4B?!od?�/�>$i�S������O}?1��?�s�?+Lv>y{h��-+�.k?�8�>����r
?�g:=�D���<+W��-��'9��.��ױ�>�8׽�:��M��zf�^i
?�-?���j�̾K׽�~��m�q=���?�(?$*�@�O��rn��qX���S��k5�ʬi������&�}q��X��6��������(��?0=O�)?Y��?�G ��fS��,5l�C�?��{\>#��>�J�>�Q�>*�A>'m
�G�1��^_�0�%����Y��>;�z?���>�WA?��;?k<a?A;A?���=%z�>9�;�`?�q=y��>V��>�>8?�g?�?��?�B?��V>��ӽ1z���P ��V?��2?#W�>�#?�Y$?�b�E���'�ܽ|�T<f#<��zp<=Ά=h�6>��K��V"��Dռ��U>�Q?�����8�ͷ��tk>��7?�}�>ڽ�>����4��+C�<��>ɭ
?-?�>����Tpr��]�I?�>���?���Gc=v�)>�8�=�j��W?ٺN7�=D:¼���=���,�;�L<�H�=*��=p�r�"B���
�:�o�;fJ�<9�>9�;?\X�>�:�>�c��p��H>x�ջ���>��>�b=��2��G��_T��6Ɂ���B>2��?���?<#E>��h=(BD>Le����[�6��1������=��?�5?:�J?c��?Z?:d(?%>�uо�Ap�=�W�5�~�QD?��?�}�>Yc#��4����p�E�?��?�Gm��)������þG���Y�=Y�2�:݋�b��}�@�Ӈ�=,��B�޽/��?���?G���R,�.O	�yF���3���UP?vn�>ke�>�y�>^)��2f�p�WF|>�?��]?�%�>P?Z{?�[[?zT>r�8�������������">�??��?Ҏ?��x?��>j>�h)�$
�z����r�f��]���o�W=c�Z>��>8�>W�>��=��Ƚ4���/>��ɣ=KFa>���>�ҥ>\��>T�w>P�<�G?G�>NF�� �0�w��#�P�}is?PP�?�G,?6s=<�V
D��������>��?K�?Z5(?8L\��f�=D��촾B�k����>�´>Ԕ�>O�=��L=�Y>�8�>.�>�h�����w9�V63�-�?B�E?R��=��ſզq���p�P���Re<����d����'C[��y�=H����i��ȩ��[�_���Fl��r�s����{����>�2�=�E�=US�=�8�< �ɼ낼<��J=l��<��=bsp���m<\�9�Yڻj_��4E"��Y<YOI=:�軄�ǾH/{?��G?��.?� B?&�m>�7>�wD���>٬b���?ەg>�� �������A�@��ʥ��^X׾/+о�b�zi����	>�$)��
>z3>z >Q3I<���=f:l=7�=��;��	=��=k��=e��=�L�=J�>�e>df�?�<��W����sb��҅<ֆ:??N9>WX>�����#?:ژ>�K|���̿�S����?��@� �?�?�=d�Q��> ׼�l"ؽ�	�;���lK�=z >����z�>i��=��H��{����=���??� @WN?V���l}߿1�W>��6>��>��R��0���\���Z� X��� ?�6;��Ͼ�H�>菹=߾�ž{!8=�]7>\�Y=l����\����=����wJ=��s=���>q9C>�'�=�������=Z'B=���=��O>v�ֻ0�B�n#�W�1=p��=��a>t�(>���>�?�^0?�Cd?�2�>�+n��%Ͼ�1���x�>���=i=�>>��=�mB>1��>"�7?f�D?��K?o�>.�=���>w��>W�,�(�m�1@�q٧�밭<���?�Ɔ?��>��U<gaA�-���k>��Ž,z?�_1?`l?4��>8~��޿ s���)��iѽi^ȼom�</R�g&ڽ����/����ӽ���=��>B�>瀧>�>�C�>��x>�k�>P
>�<�)S=$<�;<�vU�r��=���=��>vA����<�����f<<��i<$J�;�z�1��7�=�z�>s�=g�>��v=�����d>�X��b�U���=X�¾�mB���f��ru�ŵ,��	��B��=��#>_SĽ��o!�>�5>[Ն>u%�?�i?@>����X־�ܠ��W|���|�=��=��{��?=��^���N����l��>�ގ>�>l>�,�M?�-�w=n��g5���>p���S;�~M�>5q��<������ji�����D?E��4��=~?��I?W�?ɍ�>ޘ��ؾR20>`_��ߪ=���-q�Fr����?�'?#��>?쾠�D�ɾ����>Q�A��{S�������-��V�=��ɾ�S�>Ŀ��&4˾:x)�΀���<����Y�V>r�Vd�>��]?�}�?�D���[��2R������<���>5�\?BY�>#L?J/�>�&7��I�A뀾��=s�y?ގ�?^|�?- �=��=	��I��>�J?��?�?�0v?ҚM����>H�=��>빁����=�=>�z=%��=��?LR?b>	?熄�@,��:�ɤ�eJ��@8=�h=��>��\>܋�>.�=�`�=���=�Y>3�>s�>�`>@T�>�J�>o�����c�?�$�=S �>N�K?��>��?;,2�_��Z�r���A��I.��u��\k����=k"���G�%�!����>�8���.�?ޛF>s�$�\?OE��jF=�q>���=�;����> �%>J�y>y��>U��>-*>H�|>1�E>�վ��&>-%�\��D�h7b��ȳ�{~�>ۿ���0���P�E�9?���^����l�������M��Fy��'�?�#̽�n�l��VC����>N��>�:?�bԾ䏅�h�i>���>�]�>�D���ᕿ�f��I����o�?q�?�L><U�>��9?�B�>�驾��V�[�`��h����:��n�6�b��ٕ�6Ò�K�)�Zd���E<?�"K?u�:?7W�=�7D>�#r?�ᾈ�Q�|�->�U��|�2f>��?H�!�'@O�[���뢾l�!�Bi���&;?_�?ؓI? �$�=,Ž������u?|BL?�x?�?{G�?R����>�"�>%@?�2C?�H4?��>}��>Hg�=��>�n�=� 2���U�}\��\&�:D&���=�~"=<l�=��;Q������<K��F���S���'��<�ˈ���<=�=p�>3�j=�ϧ>{Xj?8��>�j>�%1?�����-�G'��k�T?,G�=�)7����|k��|� =�$l?~��?.PF? b�=��I����M>b��>\5>>SS>���>��R��N���T��X>��>w�=Vm��"��o�e\����=�_w>"'?�kS>(���,���(	�EӚ��vW>�����Ⱦ�~���L�W� �:�_�4��>�O?Xb
?n$��IpվD�|�s��I?�?�JL?��?NW��+���1�3�'�`����=]��>�%�=�@5�1���񷿓�T�zm
�֕�=����6�ž`�r>�Q'�s�˾L#i�$�b��틾۫>���j��B+���㾝ٌ��O>l��=� ���&��p��Y�����Z?_Q><���P�.�3Ѿ�ɋ=:��>~d�>z⮽-�C�|0�zM�����=�z�>y �=Su��������P��ݾ�8�>\DE?@W_?�g�?����r�>�B�V���`A��ެǼ��?[��>�m?.!B>��=���j���d��G�'�>���>g���G��1��M���$�A��>�4?��>d�?��R?��
?N�`?^
*?i:?$*�>i෽���@&?i��?@��=�Խ=�T�;9��F�Y�>j�)?!�B�.��>ă?��?��&?S�Q?+�?G�>G� �>F@�n��>S�>��W�]]����_>.�J?���>�DY?�Ճ?�>> �5�Y碾,����M�=>.�2?L2#?Ϫ?���>���>Hڡ��Ƅ=��>�zc?`^�?�o?���=N�?��0>rE�>��=��>d��>�U?�8N?[Br?��J?,��>���<Ku��~,ƽx����4�;�<,�w=��92��j��)^�<۰�;�����&�j+޼��?�4���A�Z<	�>�fr>K�����0>��ž,s��3�<>�Ǽ^͜�V����=�#�=�	>�� ?�͕>i�#���=�?�>���>����(?��?.	?�;��b��Nھ�N� �>�NA?8��=ql�?���3v�p�l=�m?`S^?��S��;���!Y?(�^?V��3��	߾�#p�bL��-yY?)�>%̮���?� R?��?��>�^X���w��r����z�	�����a=�>��ؾ�+B�\�>��?x�>ȿ?̳�=���Vj�i[���%?��?��?'�?�>�NL��쿫?��VҐ�X\?OT�>���t(?���׾�솾�|��ǧ�ȩ�JR��a��4���%�Z���muٽk�=�?4|p?�Cp?O�\?���g�ɱZ�Z#����P�!z�y��E�J�F���A��g�7��K��"���4l=�~�[G?����?b�$?ՙ(�V��>�?��l���u����16>�朾V@�r�=����1Y>=��b=vn���,��į�? ?�L�>
��>�8?�\��m<���0�k
8���ﾺ?(>�f�>	��>d!�>T�e;9�-��ٽ�ʼ�mLn���ڽ�?v>�vc?��K?ķn?�~��*1�s���=�!�>0��]��b�B>�]>v��>�W�+���=&�dX>���r�~��@x��8�	���~=Ϊ2?�)�>î�>�L�?�?с	� n���|x�8�1�@��<�)�>�i?�A�>B�>fн� �*�>�Dd?���>���>�ڥ�"  ��y��r�,��>�P�>��?e>����V��鍿����'8����={l?����x@4��>u19?��v<�<.)�>C2��"�3�[J�@ ��Ǥ=6@?].�=�G9>�'��	+�mZx�����G)?�;?Ӓ�N�*�Jz~>�."?�}�>� �>�3�?�>1Wþ�I�|�?��^?t(J?-LA?g>�>�F=U���P9Ƚ6�&���+=n��>e [>��l=�&�=���3�\���r�D=�N�=l�ϼ.U���<:ô���J<O��<� 4>J�/�M��d�Rc�{�ξ����:���n�ui���}�w�о�ȟ�H���h��$=S΁���S����f��KW�?;��?;�����7���Vo��)'���!?&Ύ�7+�;����f�g.������L�Ǿ�U6���X��쁿�j�zF'?(y��5�ǿz����yܾ$�?�b ?��y?�%���"���8�+ >ݒ�<Y��.�������ο�Y��)�^?���>�>�o/��0��>�T�>c&Y>��o>�⇾h�����<��?/�-?�o�>�Gs���ɿui��ᒧ<
��?i�@�qA?��(�\���V=\��>�	?��?>�1��%��尾�U�>�C�?^ �?+XN=��W��	�`pe?5+<��F�Dػ���=��=�=F��	�J>�D�>����9A��zܽA�4>]�>��!��b��}^�U�<�]>��ս����ք?4�\��f���/��J��	�>�T?a�>]�=�,?SH�wϿх\��aa?c:�?���?l�(?���0�>(�ܾ��M?QT6?�И>��&���t��9�=Ӥ漁9���侓=V�;��=B�>k+>�F,�y���P�L���Gd�=��K�ȿ"7*��,%�ԯi=_a=�JƼD������/fؽ#��P2i�c)�<S�=8|>�U>��>D c>a18>I(a?@r?��>��M>�L��%�����[�<�Ӆ���!��2��v!R�B篾��۾Ma;��l���>� ʾ�=���=DS������ ���c���C��d/?�K!>k�˾�M��y <�ʾ�ƨ��ׄ����S*;$�2��o���?|�B?�%��S�U�,p��u���J�W?Lz��%��&�����=2ͧ��R=AJ�>�&�=����4��R���/?I�?�ʼ�%���Qe'>K���c=9[,?5�?��.<Ͻ�>�$?�4'�����[>�x5>�I�>Q��>i��=�����aؽ�&?��U?D#��>���ђ>~u��2�w�B8r=g�>R�3��F�#Z>��<(ԋ��~�@K�����<D@W?�b�>�)�)��1Ȑ�]�!�т:=B�x?Z�?dɠ>��k?��B?p�<�|���T���
�/}=� X?Yi?�'>��}���Ͼ5æ�Ұ5?�xe?�hM>�Ji�`c꾞�.�(��=A?^�n?	y?C�����}��������&6?QVu?Al��`������r�U\�>���>��?S�;�׸�>#�5?�(��K��c�����5�ۘ?��@x�?��e=?�
����<R'?���>86�IF���Q��u���ș=���>漶�0i�a�/�S��~Q?��?�$�>Q���\�Š�=�ٕ��Z�?��?����Cg<S���l��n���<�Ϋ=�zF"�����7���ƾ��
�񪜾ῼ���>@Z@�U�s*�>�C8�U6�TϿ'��\оzSq���?Q��>��Ƚ����5�j��Pu�W�G�&�H�������>ʤ>��k鋾H����vN�-=ǽ��?6Z�=��>��G�Tݾy~���S1�?�>�	?�C�>z,�9�꼾␓?d��B���@m��r ���3?{�?࿊?�5?�ű>�U��������=�?۬N?KD_?��U������t�=%�j?�_��pU`��4�sHE��U>�"3?�B�>K�-���|=�>���>�f>�#/�y�Ŀ�ٶ����[��?��?�o���>p��?ys+?�i�8���[����*��,��<A?�2>���C�!�>0=�GҒ���
?P~0?#{�g.���k?����}�|�>?Q���_����>M�=����;��s]3���p���ͦ�����?Q@���?�5½�V3�n@>?�̃>�zB��a��Ά�]������>ݣ�>��j�)e�>��1�Rk^�u�r<T�?��?�$?�ǐ�傯�@��=�Ӂ?5c�>�҇?��>Ql�>�|�=���8a�;l_=>AR>5p���?��F?�1�>��=�M/�#��v<�t�G����E��9�>{�^?B�S?{>>{��7���!�)��z�� ��a�켞�*��i���Ͻ���=�8>�g.>#N�L���բ?F8�#ڿ�ߠ�0�/��6?�=p�?V'�������=��8?H�Y>��	��9�����b.�=%]�?f�?RA?V8���R���=Y?�0�>��W����S�a�.'y>�,?��e�o�����S����>w��?@\ì?��N���
?����犿Ζ���F�@#�wAX=*!=?o���p�>��>^�=��r�����j�w�@�>���?,K�?�'?@�h?!�n���4��Ɇ=���>}Kc?�3?}�9���Ӵ5>��>X������x� Pn?�C@��
@�D\?�����Կ�d��LF��d���>#��=5.1>{Q��S�=y� =�4�Ou=F�7>�ߗ>D%a>�	�>�lS>��:>Y->������#����0����7��������lN�`��I������F����̽�/����#��N�L�܀9��G�q劽q|�=J�Z?9hQ?:�m?Ԇ�> ����J'>�����8=��(�R��=�>81?8LH?�'?�=�=�����^� Ղ��ɮ� ����$�>]�e>5�>/��>��>0{��K>��L> �{>[�>>F�<�岺��i;0�J>���>�y�>���>�?">˅!>I��� ����Nh��ю��bs�p�??w��F�K�eZ���2��l�=�(?@��=د����ҿ�鮿�I?�����A��m�D��=UH,?P?^�!>ð���>���>�,�Z�\���=���v�x�B (��.E>x:?�_>�<v>�@4���7��JN����dw�>�4?�$���S=��u�ϤH��|ݾ��J>���>az���Z��,��E�~�Dd� �i=�;?�l?B���d���|�~��]����S>6IX>,�%=mp�=��M>U=u��u˽d�G�I(3=J�=2<`>�"?��->V�=|�>����qX�� �>p><>�_>��A?��"?�Y(����'����2���o>!��>���>�D>O|N�\�=���>Q_a>� 뼪���K��E@�BM>Ήc���d�%�|���S=���D��=N�=�����<�^Q%=�~?˅��pq�������g��~T?7? 	�x�;
�6�� ����~ �?��@�c�?y�վ��P��?2��?,�$�{Ry>eo?�g�>�����{z��n?qj{����_���E���?E��?���Ά���e�ۈx=�.?���m�>�uR�Fo����� �m���:��ʔ>Z�d?g�����V��<?�x�>-6���w����¿J"V���>s��?Z��?�����v���|{�:N?v��?}B ?�o>9Q�辽��>�%?�9B?fK�>�J �.��+7?\��?k�?��K>��?L�r?�
�>u눽�/��ٳ����zu=���;���>�\>꿾l�F�@`��R��)yj��N��&h>��%=�߸>�=�kF���Ӹ=s퇽�]����D��ҳ>�d>Y=M>�ě>4�?�s�>Ʒ�>_�=螞�`ԁ�=��v~B?��?�ľ]TM��7F�l3��k{��4?�� ?��'��%;�나>!�}?uig?��e?Z��>����v���0Ͽ�Ⱦ���=��H>�?6��>~5�c�>��+���M�>sU�>L:�x`�@끾��>�3�>�7H?�X?�b�=t�?Q�?��v>�^�>� K������DR��U�>E@�>�6?�[?G�?
���o�4��f�������P�&�=6�?[B?w�>�݋��2���wʽjPǽ�F
<L[?��a?_c����9?��w?G�E?��C?u�*>�[�6��Tɂ����>N�!?���A�1O&�L���?�F?g��>PK��7ֽ�׼W��\~���?#\?�5&?����&a��þ��<�"���M�gC�;��F��>�>����İ�=��>�۰=�Vm��X6���e<�y�=)��>�6�=T7�gq���l??Y�����Lt>=y��N���=��i>�d���-z?���=4�D��}��s����Eξ4j?s��?c�?Os�:�Y��J?��r?�/?���>�焾?^�(D��r�ٓ���Lܾ�HF> �>�#�=k���d���ғ�A^�tw�U:�\	�>���>��>�?��@>i��>�#ؾC"G�'H��fO&�c�b�Q�+���3�5������~��A�S�s���\���z{�j$�>��߽w}�>?w!?~@�=��>Q3�>��4��<z>��>9<J>>r.>���=j��=qٗ=Nto�$m2��IR?�����'���辘Ұ��4B?�md?|��>a�h�\�������r?@��?|x�?@�v>�nh��-+�Zl?�D�>�3���
?�Z:=��
�=l�<�n�����Ly��h�����>��ֽ]:�#M���f��O
?)'?����>y̾��׽X����o=M�?o�(?A�)���Q���o���W��S�}+��?h�3n����$���p�!돿�^��� ��ӝ(��i*=h�*?~�?����R��� k�P?��ef>��>�$�>�ݾ>�uI>C�	���1�t�]�fJ'�˷���O�>�X{?��=>�r?� E?|I[?��;?)��=xy�>O�����?-������>���>��*?&�?Գ�>\b?h�?2R>*�E�c�Zr��F8?��?:#?��?)�?y
��h���S=��(�?[��wx<���=��!���ph�K���w��>*V?����8�����k>x�7?	��>���>����,�� ��<2�>w�
?9G�>�  ��{r��c�KR�>$��?��|=��)>���=�����κ4J�=Ǟ����=j���u;�0R<�=1�=aYt�0����d�:G��;|Y�<^��>5Q?O��>]T�>#N��\�?�;����=\�}�'��>�;�ྋ?���(��K�N�G�;=so�?V��?D��=�0�=ym�=GV߾�L�!���0�J�<a�>�N?͊?u؎?,�L?±:?���>r� �p2��%v��ָ���(?�,?׍�>��Ԫʾ*�7�3�0�?�`?R=a�����:)���¾;ս��>L]/�;5~�	���$D�����8�� ������?绝?kpA�G�6�G��h����R����C?�#�>�e�>Z�>z�)�_�g�!#�5;>���>�R?&"�>��O?;{?�[?;qT>��8�!.���ҙ�H2��!>�@?{��?B�?$y??j�>��>�)��W��L����삾��V=pZ>���>�#�>s�>K��=fȽ�\��	�>�zg�=g�b>���>N��>��>��w>@a�<z^S?��D>|�l�uҾ��Z���`>"^�?���?��q?�ы��F��(�ܺ.��V�>��?��?ۦ?�x��ɯ">���ꆾ��]���>���>��>�`ȻmS=��>WU?f�?L�*�����vS�+,�2&?S�<?��>��ſ=q��p�9ؗ�F�u<瑾d������[�Z��=�����������[�dx��~���[��cМ��|����>〄=��=zO�=�<ü���<��J=Iۓ<�=�yn���r<��7���ػ�4���� ��'e<E K=!Y���߾ٕ�?�b?��&?�|J?�p>���>�"�b��>�5��0?���>�3==������$��w��1＾�xԾ�詾i�o�&
��o 8>wR��>ŗT>��=y0��.�=�a=��=U�k=�<=�O�=�I�=5C�=�=%��=���=V�{?��`��7�`��V=]G;?ײ>thA> ��Q1?i�>��w�cKÿ^����s?>��?��??f�?� �>- ��V
�X�<v86��b;>P�b>�և�ш�>1a�='p&�����I�ܽ�.�?	�@�4R?"���3ݿI�>"_7>�G>G�R���1��\�+%b���Y�qa!?�L;��L̾ԅ>7�=-;߾`�ƾ̮.=�=6>�`=}���N\�pz�={��4==��k=y��>yD>��=C����#�=��H=���=��O>�u����8���,�53==��=zb>�%>��>ݷ?X)?�iO?�j�>S ��A���8���_�>��<�O�>!;4�>�N�>��<?�K?GnL?�Q�>��r<���>���>_�!��V��X��FϾ�w=�ٕ?)��?Y��>�g];��@�CU�f\8���ҽ�?n�?�i�>�t�>u��Y�mZ-�Dc7�ci���t1=|��=貁���E��s����M�߻�e-�=��>���>,j�>��{>�*<>Ȑ$>J�>}p>]��}�=ly;�by�<Ӻ<��=��켙3t����/xʽ5��a|����<2Q���*;x��<��g���>b	�>$G>�w?& �;5�Ӿ-��=����ҏb���\>֩��]A��W�z�x��/�,�o���><�z>����i(��.��>VD�>ܒ�>��?WL?r�>feE���/���|����8�þ'n����L���l�-�|�D��hE��p޾���>]��>n<�>~�>L~,�6,@��>Z=J��w:8����>���"oC��M�L�q�s������b� ��;�uA?���ٔ�="}?��I?*��?��>~���ɥھ�C
>?x�"w~;l'�CYz��v���*?�1$?y��>��쾆�C�5оR�Ƚ�ܐ>�5��\U��c��E�(��KO=z˻�Q �>�줾�Oþ��1�[ă�vƐ��4J�l���)�>O<P?�!�?UG����s�6Z�M���<R��>ef?�?�>�?6?�h��̆�%ׅ�*�N=��j?@�?���?K9<>�=��6�>aT?���?/4�?�!h?���w9??{L=-G>^z#>��d>WD>��8�\m�=	��>uU?,��>Vu=L���+�.�
��1C��k�=b��<�[>#Ї>��>>j,�=�G >8�>@ϖ>l.N>��G>O�>��>9�@>������?�Z�<��>�Ge?�V�=���oƽ{#g�)���ZI��c�l`����̽=�H���Ѫ�v�7����>�ػ�:�?#T�=i�1��� ?�)6������_�>qx=�eL����>��R>m�,>�>!��>�\>]��>�=p�(�'>"h2����_L���q�]U\���>��{�d�����%�&lT��,��A��;���l��&c�%�;���?s7f�%�-��d���'��5?BM�=?�'?T�Z���v<h�S>'?=�{>������6|��ͦ��$�?Q}�?��B>?��>��@?���>SW��6�9�Sen�����$��On}�rG��܆�g8���4��_�=[T?s�]?��M?�H��=�`>;r?��(�+���L>#t{�����w>u�>������ʽ���$Ҿ�NA�$}>�}|?��?��0?0[�}E��v>	�D?5�0?T(�?�_0?a�%?n�޾�r6?;y==N��>QP�?�L=?��"?���>3�m>�'ؽ�=}�'��<m�޽�耾�\�I�<�G=�F�;�գ�!��;�2��[��컑H�#X2�# ����=r^R=��<�$R�s�/=�|�>"Z?���>�5�>m$.?��7��=�G��Ő?gW�=J<��Z������Gx����=�\?�%�?m+W?H�V>�PH���>���>�i>tU3>��s>2�>Q"��=�2����=	l
>>ɰ�=&�~�̹q�Z�ܮ��o=��(>��>�I>M2�E�#����`��^�>k;�gþ�R��*�m���"�a2�%'�>�9^?�J?7%+��P���ĕ<�!{��wS?��?Z?9j�?���/���p�#�%�V���$=��>/+j<,{8��8��OΦ�%�(����!<>�ؾ�Xm�n�r>A�?�ɿ���ꄿ��`�{-ܾ�)>X��wH���	�4�Ͼ�����h,>A�">=b�����������]6N?���=ɺ����1�^��͕=F.�>��>g;W�q_����J�����1�=67�>�.>U�������C�S�F,�>E?p_?�??G���ss�@�A�/��'����~׼�M?8�>��?C�:>�f�=G���{y�<d�M�E�!��>y��>�����G��e���d��e�$�)��>��?�b#>�*?�R?X�
?8�_?Y�(?�t?_�>�V��\���OE&?牃?,�=��ս�T���8�� F��)�>ׅ)?��B�Ќ�>�?��?��&?�yQ?�?1J>�� �_Y@���>T�>M�W��U���_>+�J?���>�-Y?-׃?T�=>9�5���sƩ�=��=�X>g�2? 1#?}�?��>���>夡�� �=-��>Wc?;�?��o?���=B�?.�1>���>S�=�g�>>f�>�?IO?��s?f�J?�z�>^4�<���q����lr�f�S�.��;��E<��y=,��t��c���<5�;�����ˀ�R��D��������;�X�>'�s>	ӕ��0>�ľ�\����@>]	�������9��P;��X�=��>��?݋�>��"�\Z�=�_�>���>���"[(?i ?-�?��;�b��۾vXK�r��>L�A?���=mm��s����u��Gd=��m?ހ^?AjV������]?��g?�D��r�J�W:׾ﻷ�,~�ܮm?�?&�ݽ>%�>a��?ߵ�?�'?ᯋ��c��f���nS�1�پ4��=�y�>��<cl��H�>�]?�د>f��>8�>"�	�lW���V��Q� ?y�?8�?�a�?���=�KM�`ѿ�*ھ�L?��>N��n�F?��L�������=����z̾=-���ؾ5	��X��|X���v������>1�
?�7n?Z�?��V?�����c��IW�=�b�U�k�
�Ұ�r\��:���:�o�h��Q߾�aþJ W���V>O�}��A�.�?��'?��.��[�>�#��)u��̾�M@>������Ö=�=����?=�~Y=h�%�.�9��`�?pҹ>�1�>��<?��[�%c=���1�`]7�����c�1>�8�>k�>�<�>�U��k�-��4�8Ⱦ����gǽM+v>!gc?ݣK?%�n?���'1�Nq����!�ٸ6��<��
`C>��
>���>��X�i ��o&��T>���r�����_��r�	���{=��2?�y�>> �>�h�?��?��	�կ���w��1�r�<��>��h?��> >��н`� ��P�>��[?GV?�?�*���R��3}�"���T�9�ʪ>O�?e5[<XJj��y�������.�R�7>"�2?T�i�	5T�_��=-�?�>�4"�*�6?�����r�Z��2ʟ����>|�A?r�=��k=?�N2��o�����K)?#Q?�ْ��*��>~>"?#��>]�>�/�?�$�>�nþ�z"�(�?�^?�2J?�MA?�3�>�>=
f��soȽ��&�$t-=	��>6�Z>�2m=���=����\��l�	�E= ��=��ϼG��3�	<������N<���<2	4>�ƿ33?��P��#����9
�֓������:�4��\���u����C����)�c��7�Z�����a����?���?|������3����[���	��>pJ!�N9�Mu����(�tl;)x��>׭��>���%�+,p�P�i�&?Sބ�ȿ�a���U���?�I?���?�.���,��3�0�>��Z<!m��d��T��sʿH����,W?f)�>�I���>ʼ���>�א>>А>e�E>�gb��N���"�=i3?P/?�� ?.I���ʿ����s=�n�?�S
@ wA?��(��쾅FV=!��>'�	?�?>7�1�G�����L�>"9�?�?� M=��W�P�	��ue?�<"�F�n�ܻf�=,|�=��=�����J>B�>���WA�jYܽ��4>�х>��"�û��^�p��<w�]>2�սά����?\�W�u�b�T�5���{�3M>CU?��>Bap=<x?��W�N�˿�J��x?�5�?2��?�=?�Iɾ�$�>�I㾞+W?ͬ.?���>��5�b;q��>pWǽyL�<0�<,^�:�
>�>�$>��1�T�.Jr�b�=�ߝ=v���D�ƿc�&������ݮ=݀�;�"�����M�4�C��O����[�>�r�I >�d>@�@>f�x>�v>��>˷U?�m?X �>�s�=�5!�*d���Ҿ��<�M��P�c��"u�gp��g�����Ѿ�X������_��WǾ��4��ܚ=\XX��ɉ�#,�`�`�ΡD�[�.?��2>ͼ㾣b>�n��;Q�Ҿ6����N��}���	��^�5���l� h�?�fH?�Ǐ��^C���� İ� Wҽ4�T?�d�	�G4��wu�=�Zj��(�<�*�>~��<�۾ۧ6���]���.?i�&?�r��W�>Xa8��=�'?�x? �C=Zb�>��)?r��8�˽)�E>�3E>���>b&�>10�=�+���o���$?��\?�S���Y�����>
ƾ�����K=�C>������.>���H���S�W=������E=�(W?t��>��)��}a������X==��x?��?%.�>o{k?��B?Kդ<+h��~�S����aw=�W?2*i?��>����	о[���D�5?�e?��N>�bh�!��<�.�]U��$?�n?4_?{~��)w}����p���n6?p�~?j�郞�y	�{3;ʻ>�Q�>ߙ?��=�؀�>"F<?�c���o���Ƽ���A�sI�?��@�2�?���h��f$?���>���>�w>��!��D���>Ҿ ��=�I�>�:¾�Qj���=�Ӯ��\�^?#ĕ?�@?�设)'���=�ؕ��Z�?��?����Og<����l��o��p�<DЫ=���G"������7�+�ƾ��
�˪��VϿ����>Z@�Q�*�>fE8�_6��SϿ����Zо^Sq�7�?��>K�Ƚ}���6�j��Ou���G���H�r����M�>��>����������{��q;�1(����>K���>1�S��&��U�����5<��>��>:��>p.���轾=ř?�b��@ο���ݝ��X?h�?�n�?�p?[�9<��v��{�����-G?��s?�Z?}r%��>]��7�"�j?�_��rU`��4�pHE��U>�"3?�B�>U�-��|=�>���>�f>�#/�w�Ŀ�ٶ�:���V��?��?�o�#��>t��?rs+?�i�8���[����*�N�+��<A?�2>'���H�!�@0=�ZҒ�Ǽ
?X~0?�z�].��n?k>a�H�g��G?�5b뼝n�>�'��a���ϽL:�� `�����L���e�?�@@ꃻ?s�׽��9��%9?�ȋ>�8ӽ����D<���=9"�>DŐ>6c��`ԙ>v�J�o�b��Ѫ=���?*��?�z?y�����5>�{?��>�C�?t��=�j�>?a�=�̶�}���
n >�w>�f%�p?�3O?��>�U�=X�<��,��,B�	�O�u����C��ǂ>-d?��L?�<f>9έ�2��"���ݽ�@/�����c7�������20>;^7>U>��B���ξ�+?���*ҿi���贄��[B?$�%>h$?���> ��0>��V?+�>9��C���wV���[w8���?VZ�?�F?<�����<:3>U?��>W��!�x�R��ݛ>L/?O�������x�n�z�]>��?v@�"�?��Y���?Z��R���Ei{������ܽ��=,ZE?����>	?���=�i�����d����>�~�? >�?f?�-d?5�{�%�2�'ғ=٩�>��S?�?~5���>Ҿ�">���>z��r쑿S	���g?2P@��@�a?@ê�7�׿m��kڳ�#����<>�?8>!��=�,r�
�=�x�=����=�#"><�>�c�>y�x>݄>�R>�h(>�$���B'��>�������&(����)����S�:$���tý��$�sʾ�|��v=�9>�Y����>6�\q���=�U?�S?(�n?>� ?�O���Y(>� �Aq==GJ��K�=�ߍ>��2?G�I?8�&?�x�=�Ӝ�}qc�7����맾����_�>WG>�T�>���>�*�>E.����G>�PF>-E�>y�>�_9=&��['=��J>0h�>���>s��>RE>Ŕ$>�.��q.���>s�����w��:��?������Q�aD��-u��Ż��	�=~�)??u�=(Ɏ��Vѿ@��צD?��e;
�MP\�C�=?/7?�oX?��X>�6ƾBK��0�>`b��YG�x��=La!�����&(��MP>�"?�ac>���>�Y/�q,@�Ţ!������>�?^aɾ�1]�����#H��v��A">��>���<{k*�wǕ���~������[=�[5?^�?�Tz��7����p�K���@�N>W�e>6��=��=RWp>��O��1@��Qz���.=P�=EY>��?M�,>�?�=9�>����'�F�k�>�-:>��,>�8>?Ys$?1}���?������y-�Nv>5<�>C�~>
m>DbI�Y̭=���>�Wf>����|�#l���@��R>������\���w��:p=f����=n6�=`Z���9��$M=��?�\��D���&. �-�"��L?%_?#،=0��;s;-�����(%˾���?�@�k�?�ݾ�ST�;}
?h+�?i2���S>�/�>a��>�7�&�x�B	?�U��T��A���P��E�?r�?;����ㆿ�"o���=�(?C�ھ��>��޽x���Kc�������=)��>��m?����g۽\Ӝ�f�?�C�> �������ʿ>�c�G�>5'�?�֒?��{�x/|��A�ۻ-?w��?�S?�<=>��ݾ��=LR�>�sD?g�O?��}>�_3�y[���+?n�?vۖ?r�H>+�?��t?�{ ?�+8��A2��
������!�y�XZ��[�>�+�=7᧾�GR�1���񍿪5k�����o>`�3=��>����;��3�m=C��m��*����>G�b>xeU>�߮>d�	?�̵>1ڀ>&<o����%������J?\�? e��1dr� $̽�Q��������#?�p?�=?�@�>oZ?|�?��G?\:�>��,�Ì��Ţ��̧��a^�=m�M>X�?��>�~^�3��>[B��O�=U��>���>��4�����
��]"����>i�K?���>l!D>�Z?��$?�8�>�P?�1a��P���F����>��r>�%?w}�?,&$?2+�4�J�����2��n	j�2�=˩f??�>��&��K�n�ۯt������B�?.�?2��=�-?�Ȋ?7V?��l?YKG>-�9<��߾������=1?!?�J��JA�@�&�%��?�Z?��>�P���6ܽ�J��������?6[?O
&?S�q2a�p�þ.��<�k4���S��M<�C3��d>7�>ҽ���<�=U$>4�=6�l�{�3��P<��=�>��=^6�+鑽�:,?1�F�Wʃ���=�r�uD���>�RL>B�����^?�^=���{����<z��U�!��?��?m�?O��l�h�'=?�??b�>DB���޾��Sw��]x��p�u�>3��>b�l�\�񏤿o���AE��ƽy���]�>,'�>���>�})?|F�>�U�>�5¾(�-��������R������+��j&����,о�4~�r>7�}���a����>��=%��>\?@�=[e�=Ӂ�>��<�w�>Z/�>t�u>�˗>��=���=d�8>�n=���MR?�����'����,ɰ��3B?ud?� �>�i�^�������x?���?Kw�?�}v>�ph�7++�Gg?OD�>f(��z
?C[:=F�"�<�d��R������kP�⮎>�!׽�:��M�>�f��]
?@'?�񍼳�̾Pz׽}���=��?��@?��$�}�X���_���O�{7d�%����b(�����p���|�	O���ފ��P��&!�R�='�%?��?�� ����!̾Z�u�7a>���>�
?A�>���>�ov>#����*��_���#�p��:��>�t?��>��X?��H?K?#�3?�gK<�>�i��c
(?��=��>{�?jp4?1�?;�>ԙ?�n ?K%>K�+��k	�3�㾞^<?� ?l;? ��>_��>�־+E�D���E=��ｆy�=A��<�^�b�����R�<'PK>!9?����{8��D���k>o�7?~R�>���> �� w����<$.�>9
?qʎ>x����=r� D����>�w�?M��M�=�*>+F�=�.��]������= ü���=�R����;�z<8��=\o�=ȟ��q���lX;Mˎ;���<�L�>�(?S(�>��O>�λ����f�U9Y>R.>��=m�)>��F�3������&#�5�>f�?���?�Y�=�	�=��j��F$�⁾��侺 X�hHw�ɵ>���>
se?_�?Pj!?>?��g<�$���Ȓ�QX��T���o��>� ,?���>�����ʾ%�O�3��?AZ?�<a�e���<)�d�¾5ս��>:[/�	.~�����D�����y���������?���?�A���6�y�z���[����C?!#�>�Y�>��>y�)���g��%�92;>���>R?��>b�O?�@{?��[?NsT>��8�K$���ә��\/�6)">�@?_��?��?�y?�]�>��>��)�OྸX���
��C�߂� �V=��Y>���>N)�>�ҩ>���=��ǽ�J����>�RT�=�b>���>���>��>�pw>r[�<�G? �>�����������߃�;�=���u?���?5d+?EN=����E��c��%8�>�i�?���?�I*?�vS�΄�=�׼�Զ���q�j�>_��>	�>�g�={�E=��>�?�>I��>�O�	b��R8���N��?�F?e��=7$ſ�1w�bg���iq��=9.����F��b����E����=	`���n����j�E�)���wk���ʵ�-+��J�P�%@�> �=�t�=�>��;������=퇤=�-�;���<~�S��Q=R[����^g��d'<�7,<��-=I��;Eѱ��>t?�W?�j*?�9?�-G>�oh>xd-�.�>�Zg=0�?銴>~�=[䨾۳T����9���O߾��޾Jj��3�����=x����=҃>��>�������=���=jCu=��8�!=k&�=��=�=�=C�=���=3>C�?.��
0����V���=�uH?�>A�2>��df?e7Y>�#h�(t��ǃ��j�?�7�?��?���>�q�u�>�~:���=�i��$N����>&t>�@��F��>��^=K0����|`��A��?M�
@�uI?9J������>��7>�:>	SR��1��T��^��DT�� ?�R;���̾E`�>3B�=����ƾ��-=��7>�P=Ef�P\����=�W��5C=�*|=�I�> G>E�=o���`f�={�J=o�=yO>I$���c;�k�;���(=u[�=k8b>y?$>4��>��?�a0?�Ud?_0�>un�Ͼ�?���D�>@��=�<�>l��=lYB>τ�>��7?�D?��K?���>yʉ=��>��>Ԙ,���m�[l徍̧��h�<���?̆?QӸ>�4R<E�A�����f>��Ž3s?�Q1?�j?��>%���ݿ2.��7���ҁ>��>:��;��۾8)>�/>2�S���i�3�t>i�>D�?͵u>�MA>��>���>�r�>(N&>V�	�ҿq>EB��<�����<%�>�x��h����cj=�Q�����l�U��\����%=������<�B=#Z�=���>&u>p�>Ú=̷��B�0>�̖���L���=:ߧ��$B�qTd��~�k�.�M55���@>��V>:O���(��&�?N�Y>3@><��?�u?�� >����վ���3�d��S�"��=d=>,�>��r;�:O`���M���Ҿ.��>�ߎ>��>�l>n,�#?�^�w=��c5���>�{�����)�:q� @�����Qi��AҺ��D?TF��ɜ�=�!~?5�I?)�?-��>���]�ؾ�80>�I��^�=��4'q�.j��M�?�'??��>t���D�oH̾���޷>y@I�-�O���K�0����Tͷ���>������оa$3��g��������B��Lr�N��>/�O?��?`:b��W��DUO�����(���q?�|g?8�>�J?�@?&���y�r��:v�=�n?Ƴ�?R=�?�>��=PT�����> �?�i�?�?�?��r?��E���>XR�:;d >�������=�>���=���=*�?0|	?!y	?񘚽vj	�N��:��b���=�k�=N+�>��>Io>���=��i=�n�=�GX>�T�>�M�>�-g>[�>�ی>��������?t��=n��>E�M?��>���M�� ���$������v��Ѡ�bo�<�ru�%u���4%����>T���"?�?��>#���q.?��Lӽ.�x>Q>a��;!��>c�=ޖ&>��>��>y*z>��>���>���j�+>?S&������^�v�P�b���ܾ�>�V��+ȓ�l��[��\��ܠ�� �Z2x���|�
5P�Ҍ��(��?���A�h7?��н��%?.��>D�E?"����x1�'k>�n�>	�>���X��҈�+�Ҿ^�?���?g�a>�C�>��`?݄?S�Q�/$M��+O�?Ml��y7�ȫ���,_����<���> �yc^��nn?��~?�V?I|�>��A>i�r?�J��#᜾]}�=�vh���6��p�>$�>�c��;%��#%4�]|���v7��yX>�Oh?=�?|�=?�,`�jɄ��
�>6t?�e1?d+?�?���?v��g�^?���>L�>уF?eU?� ?��V>Fp>��<��&��#�� ���ދ��G��e��:ڰ���0>�g*>ي��P��.*e=�Z�;�GýGֹ��<ci=�CK=mrm=���=�b>���>��^?g?��z>��?�r3���=�䏾(?���$���I>ȾƳ˾>	�U�	>�Rk?���?�ak?��>��5���:����=��s>��>�R>>�Ǌ>�;C�C�?��>uMS>t*$>�4g=iԩ���N�y6�p?����<�x>�?�s�>G�.��-C��Om��D�9�>L���QӾ�s���z��b�p$z�\�>Flp?�.*?=���f��fLc��kw��1?�3?��?E}�?hc���蘾ש!�J>L�M���s�>j�;TO�������� `!���˽|��=�P��Xm�n�r>A�?�ɿ���ꄿ��`�{-ܾ�)>X��wH���	�4�Ͼ�����h,>A�">=b�����������]6N?���=ɺ����1�^��͕=F.�>��>g;W�q_����J�����1�=67�>�.>U�������C�S�F,�>E?p_?�??G���ss�@�A�/��'����~׼�M?8�>��?C�:>�f�=G���{y�<d�M�E�!��>y��>�����G��e���d��e�$�)��>��?�b#>�*?�R?X�
?8�_?Y�(?�t?_�>�V��\���OE&?牃?,�=��ս�T���8�� F��)�>ׅ)?��B�Ќ�>�?��?��&?�yQ?�?1J>�� �_Y@���>T�>M�W��U���_>+�J?���>�-Y?-׃?T�=>9�5���sƩ�=��=�X>g�2? 1#?}�?��>���>夡�� �=-��>Wc?;�?��o?���=B�?.�1>���>S�=�g�>>f�>�?IO?��s?f�J?�z�>^4�<���q����lr�f�S�.��;��E<��y=,��t��c���<5�;�����ˀ�R��D��������;�X�>'�s>	ӕ��0>�ľ�\����@>]	�������9��P;��X�=��>��?݋�>��"�\Z�=�_�>���>���"[(?i ?-�?��;�b��۾vXK�r��>L�A?���=mm��s����u��Gd=��m?ހ^?AjV������]?��g?�D��r�J�W:׾ﻷ�,~�ܮm?�?&�ݽ>%�>a��?ߵ�?�'?ᯋ��c��f���nS�1�پ4��=�y�>��<cl��H�>�]?�د>f��>8�>"�	�lW���V��Q� ?y�?8�?�a�?���=�KM�`ѿ�*ھ�L?��>N��n�F?��L�������=����z̾=-���ؾ5	��X��|X���v������>1�
?�7n?Z�?��V?�����c��IW�=�b�U�k�
�Ұ�r\��:���:�o�h��Q߾�aþJ W���V>O�}��A�.�?��'?��.��[�>�#��)u��̾�M@>������Ö=�=����?=�~Y=h�%�.�9��`�?pҹ>�1�>��<?��[�%c=���1�`]7�����c�1>�8�>k�>�<�>�U��k�-��4�8Ⱦ����gǽM+v>!gc?ݣK?%�n?���'1�Nq����!�ٸ6��<��
`C>��
>���>��X�i ��o&��T>���r�����_��r�	���{=��2?�y�>> �>�h�?��?��	�կ���w��1�r�<��>��h?��> >��н`� ��P�>��[?GV?�?�*���R��3}�"���T�9�ʪ>O�?e5[<XJj��y�������.�R�7>"�2?T�i�	5T�_��=-�?�>�4"�*�6?�����r�Z��2ʟ����>|�A?r�=��k=?�N2��o�����K)?#Q?�ْ��*��>~>"?#��>]�>�/�?�$�>�nþ�z"�(�?�^?�2J?�MA?�3�>�>=
f��soȽ��&�$t-=	��>6�Z>�2m=���=����\��l�	�E= ��=��ϼG��3�	<������N<���<2	4>�ƿ33?��P��#����9
�֓������:�4��\���u����C����)�c��7�Z�����a����?���?|������3����[���	��>pJ!�N9�Mu����(�tl;)x��>׭��>���%�+,p�P�i�&?Sބ�ȿ�a���U���?�I?���?�.���,��3�0�>��Z<!m��d��T��sʿH����,W?f)�>�I���>ʼ���>�א>>А>e�E>�gb��N���"�=i3?P/?�� ?.I���ʿ����s=�n�?�S
@ wA?��(��쾅FV=!��>'�	?�?>7�1�G�����L�>"9�?�?� M=��W�P�	��ue?�<"�F�n�ܻf�=,|�=��=�����J>B�>���WA�jYܽ��4>�х>��"�û��^�p��<w�]>2�սά����?\�W�u�b�T�5���{�3M>CU?��>Bap=<x?��W�N�˿�J��x?�5�?2��?�=?�Iɾ�$�>�I㾞+W?ͬ.?���>��5�b;q��>pWǽyL�<0�<,^�:�
>�>�$>��1�T�.Jr�b�=�ߝ=v���D�ƿc�&������ݮ=݀�;�"�����M�4�C��O����[�>�r�I >�d>@�@>f�x>�v>��>˷U?�m?X �>�s�=�5!�*d���Ҿ��<�M��P�c��"u�gp��g�����Ѿ�X������_��WǾ��4��ܚ=\XX��ɉ�#,�`�`�ΡD�[�.?��2>ͼ㾣b>�n��;Q�Ҿ6����N��}���	��^�5���l� h�?�fH?�Ǐ��^C���� İ� Wҽ4�T?�d�	�G4��wu�=�Zj��(�<�*�>~��<�۾ۧ6���]���.?i�&?�r��W�>Xa8��=�'?�x? �C=Zb�>��)?r��8�˽)�E>�3E>���>b&�>10�=�+���o���$?��\?�S���Y�����>
ƾ�����K=�C>������.>���H���S�W=������E=�(W?t��>��)��}a������X==��x?��?%.�>o{k?��B?Kդ<+h��~�S����aw=�W?2*i?��>����	о[���D�5?�e?��N>�bh�!��<�.�]U��$?�n?4_?{~��)w}����p���n6?p�~?j�郞�y	�{3;ʻ>�Q�>ߙ?��=�؀�>"F<?�c���o���Ƽ���A�sI�?��@�2�?���h��f$?���>���>�w>��!��D���>Ҿ ��=�I�>�:¾�Qj���=�Ӯ��\�^?#ĕ?�@?�设)'���=�ؕ��Z�?��?����Og<����l��o��p�<DЫ=���G"������7�+�ƾ��
�˪��VϿ����>Z@�Q�*�>fE8�_6��SϿ����Zо^Sq�7�?��>K�Ƚ}���6�j��Ou���G���H�r����M�>��>����������{��q;�1(����>K���>1�S��&��U�����5<��>��>:��>p.���轾=ř?�b��@ο���ݝ��X?h�?�n�?�p?[�9<��v��{�����-G?��s?�Z?}r%��>]��7�"�j?�_��rU`��4�pHE��U>�"3?�B�>U�-��|=�>���>�f>�#/�w�Ŀ�ٶ�:���V��?��?�o�#��>t��?rs+?�i�8���[����*�N�+��<A?�2>'���H�!�@0=�ZҒ�Ǽ
?X~0?�z�].��n?k>a�H�g��G?�5b뼝n�>�'��a���ϽL:�� `�����L���e�?�@@ꃻ?s�׽��9��%9?�ȋ>�8ӽ����D<���=9"�>DŐ>6c��`ԙ>v�J�o�b��Ѫ=���?*��?�z?y�����5>�{?��>�C�?t��=�j�>?a�=�̶�}���
n >�w>�f%�p?�3O?��>�U�=X�<��,��,B�	�O�u����C��ǂ>-d?��L?�<f>9έ�2��"���ݽ�@/�����c7�������20>;^7>U>��B���ξ�+?���*ҿi���贄��[B?$�%>h$?���> ��0>��V?+�>9��C���wV���[w8���?VZ�?�F?<�����<:3>U?��>W��!�x�R��ݛ>L/?O�������x�n�z�]>��?v@�"�?��Y���?Z��R���Ei{������ܽ��=,ZE?����>	?���=�i�����d����>�~�? >�?f?�-d?5�{�%�2�'ғ=٩�>��S?�?~5���>Ҿ�">���>z��r쑿S	���g?2P@��@�a?@ê�7�׿m��kڳ�#����<>�?8>!��=�,r�
�=�x�=����=�#"><�>�c�>y�x>݄>�R>�h(>�$���B'��>�������&(����)����S�:$���tý��$�sʾ�|��v=�9>�Y����>6�\q���=�U?�S?(�n?>� ?�O���Y(>� �Aq==GJ��K�=�ߍ>��2?G�I?8�&?�x�=�Ӝ�}qc�7����맾����_�>WG>�T�>���>�*�>E.����G>�PF>-E�>y�>�_9=&��['=��J>0h�>���>s��>RE>Ŕ$>�.��q.���>s�����w��:��?������Q�aD��-u��Ż��	�=~�)??u�=(Ɏ��Vѿ@��צD?��e;
�MP\�C�=?/7?�oX?��X>�6ƾBK��0�>`b��YG�x��=La!�����&(��MP>�"?�ac>���>�Y/�q,@�Ţ!������>�?^aɾ�1]�����#H��v��A">��>���<{k*�wǕ���~������[=�[5?^�?�Tz��7����p�K���@�N>W�e>6��=��=RWp>��O��1@��Qz���.=P�=EY>��?M�,>�?�=9�>����'�F�k�>�-:>��,>�8>?Ys$?1}���?������y-�Nv>5<�>C�~>
m>DbI�Y̭=���>�Wf>����|�#l���@��R>������\���w��:p=f����=n6�=`Z���9��$M=��?�\��D���&. �-�"��L?%_?#،=0��;s;-�����(%˾���?�@�k�?�ݾ�ST�;}
?h+�?i2���S>�/�>a��>�7�&�x�B	?�U��T��A���P��E�?r�?;����ㆿ�"o���=�(?C�ھ��>��޽x���Kc�������=)��>��m?����g۽\Ӝ�f�?�C�> �������ʿ>�c�G�>5'�?�֒?��{�x/|��A�ۻ-?w��?�S?�<=>��ݾ��=LR�>�sD?g�O?��}>�_3�y[���+?n�?vۖ?r�H>+�?��t?�{ ?�+8��A2��
������!�y�XZ��[�>�+�=7᧾�GR�1���񍿪5k�����o>`�3=��>����;��3�m=C��m��*����>G�b>xeU>�߮>d�	?�̵>1ڀ>&<o����%������J?\�? e��1dr� $̽�Q��������#?�p?�=?�@�>oZ?|�?��G?\:�>��,�Ì��Ţ��̧��a^�=m�M>X�?��>�~^�3��>[B��O�=U��>���>��4�����
��]"����>i�K?���>l!D>�Z?��$?�8�>�P?�1a��P���F����>��r>�%?w}�?,&$?2+�4�J�����2��n	j�2�=˩f??�>��&��K�n�ۯt������B�?.�?2��=�-?�Ȋ?7V?��l?YKG>-�9<��߾������=1?!?�J��JA�@�&�%��?�Z?��>�P���6ܽ�J��������?6[?O
&?S�q2a�p�þ.��<�k4���S��M<�C3��d>7�>ҽ���<�=U$>4�=6�l�{�3��P<��=�>��=^6�+鑽�:,?1�F�Wʃ���=�r�uD���>�RL>B�����^?�^=���{����<z��U�!��?��?m�?O��l�h�'=?�??b�>DB���޾��Sw��]x��p�u�>3��>b�l�\�񏤿o���AE��ƽy���]�>,'�>���>�})?|F�>�U�>�5¾(�-��������R������+��j&����,о�4~�r>7�}���a����>��=%��>\?@�=[e�=Ӂ�>��<�w�>Z/�>t�u>�˗>��=���=d�8>�n=���MR?�����'����,ɰ��3B?ud?� �>�i�^�������x?���?Kw�?�}v>�ph�7++�Gg?OD�>f(��z
?C[:=F�"�<�d��R������kP�⮎>�!׽�:��M�>�f��]
?@'?�񍼳�̾Pz׽}���=��?��@?��$�}�X���_���O�{7d�%����b(�����p���|�	O���ފ��P��&!�R�='�%?��?�� ����!̾Z�u�7a>���>�
?A�>���>�ov>#����*��_���#�p��:��>�t?��>��X?��H?K?#�3?�gK<�>�i��c
(?��=��>{�?jp4?1�?;�>ԙ?�n ?K%>K�+��k	�3�㾞^<?� ?l;? ��>_��>�־+E�D���E=��ｆy�=A��<�^�b�����R�<'PK>!9?����{8��D���k>o�7?~R�>���> �� w����<$.�>9
?qʎ>x����=r� D����>�w�?M��M�=�*>+F�=�.��]������= ü���=�R����;�z<8��=\o�=ȟ��q���lX;Mˎ;���<�L�>�(?S(�>��O>�λ����f�U9Y>R.>��=m�)>��F�3������&#�5�>f�?���?�Y�=�	�=��j��F$�⁾��侺 X�hHw�ɵ>���>
se?_�?Pj!?>?��g<�$���Ȓ�QX��T���o��>� ,?���>�����ʾ%�O�3��?AZ?�<a�e���<)�d�¾5ս��>:[/�	.~�����D�����y���������?���?�A���6�y�z���[����C?!#�>�Y�>��>y�)���g��%�92;>���>R?��>b�O?�@{?��[?NsT>��8�K$���ә��\/�6)">�@?_��?��?�y?�]�>��>��)�OྸX���
��C�߂� �V=��Y>���>N)�>�ҩ>���=��ǽ�J����>�RT�=�b>���>���>��>�pw>r[�<�G? �>�����������߃�;�=���u?���?5d+?EN=����E��c��%8�>�i�?���?�I*?�vS�΄�=�׼�Զ���q�j�>_��>	�>�g�={�E=��>�?�>I��>�O�	b��R8���N��?�F?e��=7$ſ�1w�bg���iq��=9.����F��b����E����=	`���n����j�E�)���wk���ʵ�-+��J�P�%@�> �=�t�=�>��;������=퇤=�-�;���<~�S��Q=R[����^g��d'<�7,<��-=I��;Eѱ��>t?�W?�j*?�9?�-G>�oh>xd-�.�>�Zg=0�?銴>~�=[䨾۳T����9���O߾��޾Jj��3�����=x����=҃>��>�������=���=jCu=��8�!=k&�=��=�=�=C�=���=3>C�?.��
0����V���=�uH?�>A�2>��df?e7Y>�#h�(t��ǃ��j�?�7�?��?���>�q�u�>�~:���=�i��$N����>&t>�@��F��>��^=K0����|`��A��?M�
@�uI?9J������>��7>�:>	SR��1��T��^��DT�� ?�R;���̾E`�>3B�=����ƾ��-=��7>�P=Ef�P\����=�W��5C=�*|=�I�> G>E�=o���`f�={�J=o�=yO>I$���c;�k�;���(=u[�=k8b>y?$>4��>��?�a0?�Ud?_0�>un�Ͼ�?���D�>@��=�<�>l��=lYB>τ�>��7?�D?��K?���>yʉ=��>��>Ԙ,���m�[l徍̧��h�<���?̆?QӸ>�4R<E�A�����f>��Ž3s?�Q1?�j?��>%���ݿ2.��7���ҁ>��>:��;��۾8)>�/>2�S���i�3�t>i�>D�?͵u>�MA>��>���>�r�>(N&>V�	�ҿq>EB��<�����<%�>�x��h����cj=�Q�����l�U��\����%=������<�B=#Z�=���>&u>p�>Ú=̷��B�0>�̖���L���=:ߧ��$B�qTd��~�k�.�M55���@>��V>:O���(��&�?N�Y>3@><��?�u?�� >����վ���3�d��S�"��=d=>,�>��r;�:O`���M���Ҿ.��>�ߎ>��>�l>n,�#?�^�w=��c5���>�{�����)�:q� @�����Qi��AҺ��D?TF��ɜ�=�!~?5�I?)�?-��>���]�ؾ�80>�I��^�=��4'q�.j��M�?�'??��>t���D�oH̾���޷>y@I�-�O���K�0����Tͷ���>������оa$3��g��������B��Lr�N��>/�O?��?`:b��W��DUO�����(���q?�|g?8�>�J?�@?&���y�r��:v�=�n?Ƴ�?R=�?�>��=PT�����> �?�i�?�?�?��r?��E���>XR�:;d >�������=�>���=���=*�?0|	?!y	?񘚽vj	�N��:��b���=�k�=N+�>��>Io>���=��i=�n�=�GX>�T�>�M�>�-g>[�>�ی>��������?t��=n��>E�M?��>���M�� ���$������v��Ѡ�bo�<�ru�%u���4%����>T���"?�?��>#���q.?��Lӽ.�x>Q>a��;!��>c�=ޖ&>��>��>y*z>��>���>���j�+>?S&������^�v�P�b���ܾ�>�V��+ȓ�l��[��\��ܠ�� �Z2x���|�
5P�Ҍ��(��?���A�h7?��н��%?.��>D�E?"����x1�'k>�n�>	�>���X��҈�+�Ҿ^�?���?g�a>�C�>��`?݄?S�Q�/$M��+O�?Ml��y7�ȫ���,_����<���> �yc^��nn?��~?�V?I|�>��A>i�r?�J��#᜾]}�=�vh���6��p�>$�>�c��;%��#%4�]|���v7��yX>�Oh?=�?|�=?�,`�jɄ��
�>6t?�e1?d+?�?���?v��g�^?���>L�>уF?eU?� ?��V>Fp>��<��&��#�� ���ދ��G��e��:ڰ���0>�g*>ي��P��.*e=�Z�;�GýGֹ��<ci=�CK=mrm=���=�b>���>��^?g?��z>��?�r3���=�䏾(?���$���I>ȾƳ˾>	�U�	>�Rk?���?�ak?��>��5���:����=��s>��>�R>>�Ǌ>�;C�C�?��>uMS>t*$>�4g=iԩ���N�y6�p?����<�x>�?�s�>G�.��-C��Om��D�9�>L���QӾ�s���z��b�p$z�\�>Flp?�.*?=���f��fLc��kw��1?�3?��?E}�?hc���蘾ש!�J>L�M���s�>j�;TO�������� `!���˽|��=�P��Xm�n�r>A�?�ɿ���ꄿ��`�{-ܾ�)>X��wH���	�4�Ͼ�����h,>A�">=b�����������]6N?���=ɺ����1�^��͕=F.�>��>g;W�q_����J�����1�=67�>�.>U�������C�S�F,�>E?p_?�??G���ss�@�A�/��'����~׼�M?8�>��?C�:>�f�=G���{y�<d�M�E�!��>y��>�����G��e���d��e�$�)��>��?�b#>�*?�R?X�
?8�_?Y�(?�t?_�>�V��\���OE&?牃?,�=��ս�T���8�� F��)�>ׅ)?��B�Ќ�>�?��?��&?�yQ?�?1J>�� �_Y@���>T�>M�W��U���_>+�J?���>�-Y?-׃?T�=>9�5���sƩ�=��=�X>g�2? 1#?}�?��>���>夡�� �=-��>Wc?;�?��o?���=B�?.�1>���>S�=�g�>>f�>�?IO?��s?f�J?�z�>^4�<���q����lr�f�S�.��;��E<��y=,��t��c���<5�;�����ˀ�R��D��������;�X�>'�s>	ӕ��0>�ľ�\����@>]	�������9��P;��X�=��>��?݋�>��"�\Z�=�_�>���>���"[(?i ?-�?��;�b��۾vXK�r��>L�A?���=mm��s����u��Gd=��m?ހ^?AjV������]?��g?�D��r�J�W:׾ﻷ�,~�ܮm?�?&�ݽ>%�>a��?ߵ�?�'?ᯋ��c��f���nS�1�پ4��=�y�>��<cl��H�>�]?�د>f��>8�>"�	�lW���V��Q� ?y�?8�?�a�?���=�KM�`ѿ�*ھ�L?��>N��n�F?��L�������=����z̾=-���ؾ5	��X��|X���v������>1�
?�7n?Z�?��V?�����c��IW�=�b�U�k�
�Ұ�r\��:���:�o�h��Q߾�aþJ W���V>O�}��A�.�?��'?��.��[�>�#��)u��̾�M@>������Ö=�=����?=�~Y=h�%�.�9��`�?pҹ>�1�>��<?��[�%c=���1�`]7�����c�1>�8�>k�>�<�>�U��k�-��4�8Ⱦ����gǽM+v>!gc?ݣK?%�n?���'1�Nq����!�ٸ6��<��
`C>��
>���>��X�i ��o&��T>���r�����_��r�	���{=��2?�y�>> �>�h�?��?��	�կ���w��1�r�<��>��h?��> >��н`� ��P�>��[?GV?�?�*���R��3}�"���T�9�ʪ>O�?e5[<XJj��y�������.�R�7>"�2?T�i�	5T�_��=-�?�>�4"�*�6?�����r�Z��2ʟ����>|�A?r�=��k=?�N2��o�����K)?#Q?�ْ��*��>~>"?#��>]�>�/�?�$�>�nþ�z"�(�?�^?�2J?�MA?�3�>�>=
f��soȽ��&�$t-=	��>6�Z>�2m=���=����\��l�	�E= ��=��ϼG��3�	<������N<���<2	4>�ƿ33?��P��#����9
�֓������:�4��\���u����C����)�c��7�Z�����a����?���?|������3����[���	��>pJ!�N9�Mu����(�tl;)x��>׭��>���%�+,p�P�i�&?Sބ�ȿ�a���U���?�I?���?�.���,��3�0�>��Z<!m��d��T��sʿH����,W?f)�>�I���>ʼ���>�א>>А>e�E>�gb��N���"�=i3?P/?�� ?.I���ʿ����s=�n�?�S
@ wA?��(��쾅FV=!��>'�	?�?>7�1�G�����L�>"9�?�?� M=��W�P�	��ue?�<"�F�n�ܻf�=,|�=��=�����J>B�>���WA�jYܽ��4>�х>��"�û��^�p��<w�]>2�սά����?\�W�u�b�T�5���{�3M>CU?��>Bap=<x?��W�N�˿�J��x?�5�?2��?�=?�Iɾ�$�>�I㾞+W?ͬ.?���>��5�b;q��>pWǽyL�<0�<,^�:�
>�>�$>��1�T�.Jr�b�=�ߝ=v���D�ƿc�&������ݮ=݀�;�"�����M�4�C��O����[�>�r�I >�d>@�@>f�x>�v>��>˷U?�m?X �>�s�=�5!�*d���Ҿ��<�M��P�c��"u�gp��g�����Ѿ�X������_��WǾ��4��ܚ=\XX��ɉ�#,�`�`�ΡD�[�.?��2>ͼ㾣b>�n��;Q�Ҿ6����N��}���	��^�5���l� h�?�fH?�Ǐ��^C���� İ� Wҽ4�T?�d�	�G4��wu�=�Zj��(�<�*�>~��<�۾ۧ6���]���.?i�&?�r��W�>Xa8��=�'?�x? �C=Zb�>��)?r��8�˽)�E>�3E>���>b&�>10�=�+���o���$?��\?�S���Y�����>
ƾ�����K=�C>������.>���H���S�W=������E=�(W?t��>��)��}a������X==��x?��?%.�>o{k?��B?Kդ<+h��~�S����aw=�W?2*i?��>����	о[���D�5?�e?��N>�bh�!��<�.�]U��$?�n?4_?{~��)w}����p���n6?p�~?j�郞�y	�{3;ʻ>�Q�>ߙ?��=�؀�>"F<?�c���o���Ƽ���A�sI�?��@�2�?���h��f$?���>���>�w>��!��D���>Ҿ ��=�I�>�:¾�Qj���=�Ӯ��\�^?#ĕ?�@?�设)'���=�ؕ��Z�?��?����Og<����l��o��p�<DЫ=���G"������7�+�ƾ��
�˪��VϿ����>Z@�Q�*�>fE8�_6��SϿ����Zо^Sq�7�?��>K�Ƚ}���6�j��Ou���G���H�r����M�>��>����������{��q;�1(����>K���>1�S��&��U�����5<��>��>:��>p.���轾=ř?�b��@ο���ݝ��X?h�?�n�?�p?[�9<��v��{�����-G?��s?�Z?}r%��>]��7�"�j?�_��rU`��4�pHE��U>�"3?�B�>U�-��|=�>���>�f>�#/�w�Ŀ�ٶ�:���V��?��?�o�#��>t��?rs+?�i�8���[����*�N�+��<A?�2>'���H�!�@0=�ZҒ�Ǽ
?X~0?�z�].��n?k>a�H�g��G?�5b뼝n�>�'��a���ϽL:�� `�����L���e�?�@@ꃻ?s�׽��9��%9?�ȋ>�8ӽ����D<���=9"�>DŐ>6c��`ԙ>v�J�o�b��Ѫ=���?*��?�z?y�����5>�{?��>�C�?t��=�j�>?a�=�̶�}���
n >�w>�f%�p?�3O?��>�U�=X�<��,��,B�	�O�u����C��ǂ>-d?��L?�<f>9έ�2��"���ݽ�@/�����c7�������20>;^7>U>��B���ξ�+?���*ҿi���贄��[B?$�%>h$?���> ��0>��V?+�>9��C���wV���[w8���?VZ�?�F?<�����<:3>U?��>W��!�x�R��ݛ>L/?O�������x�n�z�]>��?v@�"�?��Y���?Z��R���Ei{������ܽ��=,ZE?����>	?���=�i�����d����>�~�? >�?f?�-d?5�{�%�2�'ғ=٩�>��S?�?~5���>Ҿ�">���>z��r쑿S	���g?2P@��@�a?@ê�7�׿m��kڳ�#����<>�?8>!��=�,r�
�=�x�=����=�#"><�>�c�>y�x>݄>�R>�h(>�$���B'��>�������&(����)����S�:$���tý��$�sʾ�|��v=�9>�Y����>6�\q���=�U?�S?(�n?>� ?�O���Y(>� �Aq==GJ��K�=�ߍ>��2?G�I?8�&?�x�=�Ӝ�}qc�7����맾����_�>WG>�T�>���>�*�>E.����G>�PF>-E�>y�>�_9=&��['=��J>0h�>���>s��>RE>Ŕ$>�.��q.���>s�����w��:��?������Q�aD��-u��Ż��	�=~�)??u�=(Ɏ��Vѿ@��צD?��e;
�MP\�C�=?/7?�oX?��X>�6ƾBK��0�>`b��YG�x��=La!�����&(��MP>�"?�ac>���>�Y/�q,@�Ţ!������>�?^aɾ�1]�����#H��v��A">��>���<{k*�wǕ���~������[=�[5?^�?�Tz��7����p�K���@�N>W�e>6��=��=RWp>��O��1@��Qz���.=P�=EY>��?M�,>�?�=9�>����'�F�k�>�-:>��,>�8>?Ys$?1}���?������y-�Nv>5<�>C�~>
m>DbI�Y̭=���>�Wf>����|�#l���@��R>������\���w��:p=f����=n6�=`Z���9��$M=��?�\��D���&. �-�"��L?%_?#،=0��;s;-�����(%˾���?�@�k�?�ݾ�ST�;}
?h+�?i2���S>�/�>a��>�7�&�x�B	?�U��T��A���P��E�?r�?;����ㆿ�"o���=�(?C�ھ��>��޽x���Kc�������=)��>��m?����g۽\Ӝ�f�?�C�> �������ʿ>�c�G�>5'�?�֒?��{�x/|��A�ۻ-?w��?�S?�<=>��ݾ��=LR�>�sD?g�O?��}>�_3�y[���+?n�?vۖ?r�H>+�?��t?�{ ?�+8��A2��
������!�y�XZ��[�>�+�=7᧾�GR�1���񍿪5k�����o>`�3=��>����;��3�m=C��m��*����>G�b>xeU>�߮>d�	?�̵>1ڀ>&<o����%������J?\�? e��1dr� $̽�Q��������#?�p?�=?�@�>oZ?|�?��G?\:�>��,�Ì��Ţ��̧��a^�=m�M>X�?��>�~^�3��>[B��O�=U��>���>��4�����
��]"����>i�K?���>l!D>�Z?��$?�8�>�P?�1a��P���F����>��r>�%?w}�?,&$?2+�4�J�����2��n	j�2�=˩f??�>��&��K�n�ۯt������B�?.�?2��=�-?�Ȋ?7V?��l?YKG>-�9<��߾������=1?!?�J��JA�@�&�%��?�Z?��>�P���6ܽ�J��������?6[?O
&?S�q2a�p�þ.��<�k4���S��M<�C3��d>7�>ҽ���<�=U$>4�=6�l�{�3��P<��=�>��=^6�+鑽�:,?1�F�Wʃ���=�r�uD���>�RL>B�����^?�^=���{����<z��U�!��?��?m�?O��l�h�'=?�??b�>DB���޾��Sw��]x��p�u�>3��>b�l�\�񏤿o���AE��ƽy���]�>,'�>���>�})?|F�>�U�>�5¾(�-��������R������+��j&����,о�4~�r>7�}���a����>��=%��>\?@�=[e�=Ӂ�>��<�w�>Z/�>t�u>�˗>��=���=d�8>�n=���MR?�����'����,ɰ��3B?ud?� �>�i�^�������x?���?Kw�?�}v>�ph�7++�Gg?OD�>f(��z
?C[:=F�"�<�d��R������kP�⮎>�!׽�:��M�>�f��]
?@'?�񍼳�̾Pz׽}���=��?��@?��$�}�X���_���O�{7d�%����b(�����p���|�	O���ފ��P��&!�R�='�%?��?�� ����!̾Z�u�7a>���>�
?A�>���>�ov>#����*��_���#�p��:��>�t?��>��X?��H?K?#�3?�gK<�>�i��c
(?��=��>{�?jp4?1�?;�>ԙ?�n ?K%>K�+��k	�3�㾞^<?� ?l;? ��>_��>�־+E�D���E=��ｆy�=A��<�^�b�����R�<'PK>!9?����{8��D���k>o�7?~R�>���> �� w����<$.�>9
?qʎ>x����=r� D����>�w�?M��M�=�*>+F�=�.��]������= ü���=�R����;�z<8��=\o�=ȟ��q���lX;Mˎ;���<�L�>�(?S(�>��O>�λ����f�U9Y>R.>��=m�)>��F�3������&#�5�>f�?���?�Y�=�	�=��j��F$�⁾��侺 X�hHw�ɵ>���>
se?_�?Pj!?>?��g<�$���Ȓ�QX��T���o��>� ,?���>�����ʾ%�O�3��?AZ?�<a�e���<)�d�¾5ս��>:[/�	.~�����D�����y���������?���?�A���6�y�z���[����C?!#�>�Y�>��>y�)���g��%�92;>���>R?��>b�O?�@{?��[?NsT>��8�K$���ә��\/�6)">�@?_��?��?�y?�]�>��>��)�OྸX���
��C�߂� �V=��Y>���>N)�>�ҩ>���=��ǽ�J����>�RT�=�b>���>���>��>�pw>r[�<�G? �>�����������߃�;�=���u?���?5d+?EN=����E��c��%8�>�i�?���?�I*?�vS�΄�=�׼�Զ���q�j�>_��>	�>�g�={�E=��>�?�>I��>�O�	b��R8���N��?�F?e��=7$ſ�1w�bg���iq��=9.����F��b����E����=	`���n����j�E�)���wk���ʵ�-+��J�P�%@�> �=�t�=�>��;������=퇤=�-�;���<~�S��Q=R[����^g��d'<�7,<��-=I��;Eѱ��>t?�W?�j*?�9?�-G>�oh>xd-�.�>�Zg=0�?銴>~�=[䨾۳T����9���O߾��޾Jj��3�����=x����=҃>��>�������=���=jCu=��8�!=k&�=��=�=�=C�=���=3>C�?.��
0����V���=�uH?�>A�2>��df?e7Y>�#h�(t��ǃ��j�?�7�?��?���>�q�u�>�~:���=�i��$N����>&t>�@��F��>��^=K0����|`��A��?M�
@�uI?9J������>��7>�:>	SR��1��T��^��DT�� ?�R;���̾E`�>3B�=����ƾ��-=��7>�P=Ef�P\����=�W��5C=�*|=�I�> G>E�=o���`f�={�J=o�=yO>I$���c;�k�;���(=u[�=k8b>y?$>4��>��?�a0?�Ud?_0�>un�Ͼ�?���D�>@��=�<�>l��=lYB>τ�>��7?�D?��K?���>yʉ=��>��>Ԙ,���m�[l徍̧��h�<���?̆?QӸ>�4R<E�A�����f>��Ž3s?�Q1?�j?��>%���ݿ2.��7���ҁ>��>:��;��۾8)>�/>2�S���i�3�t>i�>D�?͵u>�MA>��>���>�r�>(N&>V�	�ҿq>EB��<�����<%�>�x��h����cj=�Q�����l�U��\����%=������<�B=#Z�=���>&u>p�>Ú=̷��B�0>�̖���L���=:ߧ��$B�qTd��~�k�.�M55���@>��V>:O���(��&�?N�Y>3@><��?�u?�� >����վ���3�d��S�"��=d=>,�>��r;�:O`���M���Ҿ.��>�ߎ>��>�l>n,�#?�^�w=��c5���>�{�����)�:q� @�����Qi��AҺ��D?TF��ɜ�=�!~?5�I?)�?-��>���]�ؾ�80>�I��^�=��4'q�.j��M�?�'??��>t���D�oH̾���޷>y@I�-�O���K�0����Tͷ���>������оa$3��g��������B��Lr�N��>/�O?��?`:b��W��DUO�����(���q?�|g?8�>�J?�@?&���y�r��:v�=�n?Ƴ�?R=�?�>��=PT�����> �?�i�?�?�?��r?��E���>XR�:;d >�������=�>���=���=*�?0|	?!y	?񘚽vj	�N��:��b���=�k�=N+�>��>Io>���=��i=�n�=�GX>�T�>�M�>�-g>[�>�ی>��������?t��=n��>E�M?��>���M�� ���$������v��Ѡ�bo�<�ru�%u���4%����>T���"?�?��>#���q.?��Lӽ.�x>Q>a��;!��>c�=ޖ&>��>��>y*z>��>���>���j�+>?S&������^�v�P�b���ܾ�>�V��+ȓ�l��[��\��ܠ�� �Z2x���|�
5P�Ҍ��(��?���A�h7?��н��%?.��>D�E?"����x1�'k>�n�>	�>���X��҈�+�Ҿ^�?���?g�a>�C�>��`?݄?S�Q�/$M��+O�?Ml��y7�ȫ���,_����<���> �yc^��nn?��~?�V?I|�>��A>i�r?�J��#᜾]}�=�vh���6��p�>$�>�c��;%��#%4�]|���v7��yX>�Oh?=�?|�=?�,`�jɄ��
�>6t?�e1?d+?�?���?v��g�^?���>L�>уF?eU?� ?��V>Fp>��<��&��#�� ���ދ��G��e��:ڰ���0>�g*>ي��P��.*e=�Z�;�GýGֹ��<ci=�CK=mrm=���=�b>���>��^?g?��z>��?�r3���=�䏾(?���$���I>ȾƳ˾>	�U�	>�Rk?���?�ak?��>��5���:����=��s>��>�R>>�Ǌ>�;C�C�?��>uMS>t*$>�4g=iԩ���N�y6�p?����<�x>�?�s�>G�.��-C��Om��D�9�>L���QӾ�s���z��b�p$z�\�>Flp?�.*?=���f��fLc��kw��1?�3?��?E}�?hc���蘾ש!�J>L�M���s�>j�;TO�������� `!���˽|��=�P��۠�J\b>˹��l޾��n��J�w��8DM=7��@V=���־$0�ɗ�=q
>����� ����Ԫ��0J?��j=�v���XU�9s����>���>ޮ>��:���v�6�@�ͭ��[B�=l��>� ;>^S�����_~G��7��g�>�.T?��a?<΍?��ݾP�����N���ǡ�O�6>���>��e>y�?s�!>2I����6J2������10�+t�>o��>~�?�bvu������� ����D�>1�?�v�>A�9?Hzo?�%�>�)�?txY?��?3ߨ>�e#��|�"/.?��?3��<ק���a���nA���5��+?�2?R�-�Y�V>�
?�}"?��=?ŦP?�?��:=v �B:o��R�>lZ�>kS[�1ڸ��I�>��r?v��>�j?�E�?��=��-��ү�P�ڽb�l>Qxc>X�1?�+?�� ?���>��>�����
�=���>a�g?���?n?V��=�-?x(>�&�>M��=
Z�>�c�>	�?��L?�8q?C�G?6��>P�<mI��Ѻ�P�j�v3������;�{=8��sXX��=鼔�=�FD<�����/���
���d�f\<�_�>��s>�	����0>��ľ�O��?�@>Ӊ���O���ڊ�C�:�_޷=���>��?���>�X#�͸�=خ�>�H�>?��$7(?��?�?$";<�b�^�ھ�K���>�B?���=��l�h���8�u���g=j�m?D�^?��W�<&��Zc?J�g?��߾S�9� Y���^ᾆ�@?�
?nֽ��>9�v?��q?��?�96���\��y��`x�꘰����=��>�_,����U]�>�9H?�۫>'M�>�z�>�Z����d�b���3�>��?�?xx�?��K>Q�\������8_��SV?���>�Ӿ�L�?���������e|��@Ͼ����QD��۬��x������3`���Ɲ!=Ҕ?���?�Qu?��_?;����s��Ga�K{��kV�Z*���	�}�?��u=�i�9��v�ʹ�����\宾*B=�S��C��Y�?��?XQb��#?`"��̂��X��F^>�^���'��u뻊��:�<�[9=L�<��J3�����kO!?K��>�>�~E?��\��?�`q8�<�������=�>���>�&�>���;;2��,�ڡ�����ҽ>|>7�e?� P?(�q?��-:6�j|��#sD�洶�d�=���=륏> ^�2�P��,�|I�ķu�O�߆����5|g=�
5?%s[>ڳ�>�m�?
��>W0	�S)��տ��D�,�ۤp=zܹ>,�c?.4�>>n�>����ye�f��>s>n?�?ӕ�>4a���:.����r�E��R�>��[>���>���=�j\��Z\�{��ѣ��x�N�@�<�RW?��Q��r1�fp>��\?Iqܻ&�켘��>���=0�����Z������<5?�7^>�+>����*��"j���!��7/?��?����b@��ח>q3?<�>]��>�с?��u>�%q�xY�>=0?�d?H+K?_3?��>�ƽÌ��+���֓�,��=S��>���>�y,>l�<��[��j��������S>`�=����/�=�м��<~����>�aֿ�LG�Wp;�p�X�����[��0�$p��\f�?��w�����l�g�Eս��F�]Kv������n�H�?���?C]�����Y���Ȁ����-��>x&���&ݽ�y��ߟu��4��S���X��7�d�]��w�|4J�N�'?�����ǿ򰡿�:ܾ ! ?	B ?A�y?��3�"���8�� >D�<�-����뾶����ο%����^?���>��0��S��>ܥ�>Y�X>Iq>����螾�2�<��?I�-?8��>Ўr�#�ɿV����Ĥ<���?+�@}A?��(�=�쾓V=���>��	?��?>�S1�dH�����jU�>�<�?��?N�M=B�W���	��e?�b<��F���ݻd�=?�=�S=���y�J>�T�>���TA�Q>ܽ
�4>�څ>Ww"�֬���^�1}�<�]>k�ս�4���؄?�;\�z!f���/��|���>�T?Sf�>�J�=�-?MIH�,�Ͽ�]�$�`?�&�?���?�H)?�	��^��>��ܾ�:M?�X6?C�>E�&�R�t���=�A�5L��~�⾝�V���=���>R>�-�LU��IQ��H��Y%�=�����Ŀ�+�1<�jK�ǳؼRD<h�5�k̕��׼�����c�t�ν�N=�>c�h><ς>�@m>�RC>6R?�:y?Pu�>~�->��%������ľ��-��č�>�N3>��n\�;���_m�����6�	������*��I˾:!=���=c6R�'���F� ���b�ږF�G�.?;v$>��ʾ��M�er-<pʾg����󄼤䥽�.̾]�1��!n�y͟?c�A?�����V�*���Z�����O�W?�P�����묾C��=���#�=�#�>5��=��⾁ 3�(}S��}0?��?8%������,>h����%=q'+?$�?f�N<�c�><.&?/)%�[ܽ%^>Uw4>At�>pq�>� 	>�C��~V�]�?R#U?������W��>$4���z�`s^=N8>-�4��u�*�Y>T�<����/�N�BA���!�<�(W?כ�>��)�>�"a��U���Y==��x?Ԓ?�-�>p{k?�B?�ݤ<sg��'�S����aw=��W?�)i?3�>���6	о����:�5?ޣe?�N>�ch�9���.�BU��$?'�n?�^?�~���v}�^��g��o6?R�x?r(B��߫���	���k��>�>F?\/?�L����>�C?��nf����¿����|�?��
@c'@ �=�������<��?�S�>u+��󴋾��2��뢾5Ƚ��?7���A���uX�|����P? �?�?9����B���>W���%�?�Ԅ?��ľ{��<���iSR�}Z�Ba����=�덽 ��� ���7�r�ž����ݒ����\]m>9b@l�Z8�>F:���𿢑ɿŎ�eʖ�NN��Ϯ?5��>�kɽn�����h���a���8�ux+��v`��P�>��>��������O�{�v;��-����>Q	�p�>.�S�"��������5<t�>��>ư�>�Q��T뽾Rę?A]���@οK���$����X?�e�?�n�?�t?'&9<��v���{�t��!3G?(�s?�Z?�[%��?]�%8�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�d�|=�>���>g>�#/�y�Ŀ�ٶ�>���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�TҒ�¼
?W~0?{�f.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\� N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>gH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?=�>=�?� �=.�>�%�=����u-�ON#>D��=�$?���?��M?W��>p@�=�[8�H�.�?F��KR����C�vχ>�a?��L?��b>�y����2�"� �UOͽ)`1����IZ@�n#,���߽I5>Z�=>	>��D�+�Ҿ�Q$?��ྑ	����w^����?��?��?����@��뻽�ie?���>x$�?P��S���i����?�A@�T
?�-��B���(>8Y�>��>���uoɽG�J�!�S>ߗH?�$�<�z��	Z���[�>u�?�X@y��?>|�b�?e[�0b���$z�2 �Q|"�K�t>0�D?|��s>�R�>�!>��q�e#���f]�9ڸ>e��?%O�?
�?�)c?"eg�]q*��xm=rr�>�fc?!p�> �Z=!��{�8>iT?�� �w���w��C??�@.9@��_?�����ؿE�hD��A�߾�q=X��=�0�=�����=4潪/V=r�C<��>��>&1�>�Ƃ>{I>��;>��=���F�#�r��{I��U�5�����T��%�����r�`�۾ut��+a��B�2�}�Ľq�ݽ�k�	�-��������=�*P?Q�P?�eo?�.?�B@�h>`��.[�=[�%��O�=<�>�2?6M?��*?�Х=�|��ݡb�ǟ������؈��3�>�2G>�q�>1��>NN�>���<�k>�B?>2s>�>�/=�W�<,��=�S>�Ǭ>���>�-�>�F<>n�>�δ�42���h��w�̽#�?�~����J��1��9������ru�=|b.?}>���?п����1H?�����)��+�J�>8�0?bcW?�>`����T�9>K��æj��b>�( ��|l��)��)Q>l?��f>�u>�3�Cd8�$�P��z��+k|>�36?붾SJ9��u���H��fݾ];M>��>5;D�ek��������ui�Z�{=6y:?;�?�:���ް���u�r@��uRR>G?\>B�=�m�=�[M>mCc���ƽdH�>q.=g��=�^>�T?Һ+>b�=�ߣ>BR����O�c�>:�B>*>,>	@?�!%?�m��ڗ��}��.�-��w>iG�>���>S&>pBJ����=@e�>f�a>��)΃�r����?���W>9~�$�_�U<u�*�x=@З��B�=�;�=�k ��=�%=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿܚ�>�Iy�U���JW��2+��#;ʽ�� ?�h?%R��ӽmϛ�D=�>���>@��Ba����ԿU}�����>��?�x�?��D�����Z@��%�>#�?��?�3>�~�R��(��>�,c?�Mn?��>g���]%>�$�?�S�?�3�?-s>@��?yF�?�D�>T8O��5\������ȉ����<��	�Q@�����jV��䧿=ᆿf�m�Ѓ߾#�">,�<î�>ւ��D��м\�*���A�QZ�{1/>=�8>ӝ{<��=>�j?U�>��>��������ߺ��F��R?��?5�C����<���=[�#�§(?�K?�=	<�#���"�>��\?�`�?�g`?T4�>�����9�����������f>���>��?!uD>�`>��򾻩9�T�G>
��>��?>Y猾=���(��gS�>\ ?� ?Yӷ>�� ?Т#?��j>�<�>[fE�">����E�I��>���>{J?`�~?l�?����4T3����a硿��[�(�M>��x?�R?�Ε>􎏿n����3E��I�����U��?�vg?3当�?:/�?��??�A?:bf>Z�ؾ�ݭ��΀>v�!?����A�dM&�:��~?�O?��>~#��&�ս4ּm���z��� ?�(\?&A&?���+a���¾E*�<#�ؚU�1l�;�LD�'�>��>D������=q>wѰ=�Im��A6�}g<�v�=��>��=�/7�l��B,7?��0;�����z�����N(��̩>��D>x4'��`�?�l�s���)����a��o��O��?DF�?%?p�.>� r�G�3?�w?.X*?a!?�d��O���!�6�I�r���d"�K�>���>-e��%�?�����c0��[Ĕ��|��k���/ ?�{�>*d�>�4?�>�i�>��[�e�+��|����n��<.�uWU�s�:���_�����$II�(�þEa�����>�4��w�>�|?Q[>��>��>9��=,�>F�_>퉞>�]�>�R>p� >��>���=�3d��KR?��� �'��������3B?�qd?1�>�i�������ހ?���?Js�?>v>�~h��,+�n?�>�>i���p
?�W:=��BF�<xU��ڽ��2��5��>F׽� :�XM�nf�j
?�/?�����̾�:׽�]���:k=*L�?�O$?Y�)���U�`�i�<�S�E O��5e��
}�����$�6[m�Ƹ��Ȑ���샿ϱ*�p�"=�*.?ɟ�?�/����x骾�yi�x'7�zb�>e�>�f�>��>�/1>�
���0��*^��`/�$���M:�>�(?*�>-�>?$�"?�f9?�r?�b?d>��ȹ?�0ý�5�>��?jTW?�$??BH?�Y?��?kt�=T�i7����۾/�0?�1?�O
?}
�>��>h�n�	9���^�8m5>]󗾵lb�Vi�;ja��`������~>:��<8Y?���8�8�i���k>��7? �>���>����,����<��>`�
?�H�>���`|r�.b��R�>��?��\n=d�)>!�=ff����к�S�=����-�=�0���;�bu<2��=��=k�s��o��%z�:�0�;���< �>\�?���>��>�͆��&��e�A��=��W>��O>�>(ھL������Ɉh���w>�ۏ? ճ?�b=k�=Ne�=����SO¾M��㾾��<I�?�$?�S?ԉ�?=?�f#?�� >:q�W���>�����(?j!,?a��>7��Բʾ����3�ɝ?<[?x<a���� <)�;�¾~�Խf�>\/�v/~����aD��酻���e����?㿝?A�b�6�Yx�ÿ���[����C?�!�>Y�>��>�)�.�g�8%�!2;>���>)R?|��>�9N?K�z?J�[?��X>�6�O[������Z���@>n??��?�~�?]x?'j�>z�>۶)�<�߾&����p#����`��r�R=
#W>0
�>7 �>�'�>�o�=B�Ľ�I���?�ݾ�=��i>'��>�>Ƞ�>#~q>�͓<��G?C��>�]��F��E줾�Ń�

=�4�u?曐?ő+?/U=4���E�wG���J�>ho�?���?4*?��S���=7�ּTⶾ��q��%�>۹>�1�>�Ɠ=�xF=Qb>��>Ԡ�>)�(a��q8��QM���?�F?���=G�ſŵq�K�p��͗�F�a<ƒ�] e�|���*[�J��=�Ø����թ���[� ����h��gص��x��c�{����>�ņ= ��=�|�=T��<2�ʼ���<��J=���<Q�=��p�k{l<��8�pgѻ5ǈ��y��]<��H=�7���jʾB�|?&8I?��+?��C?��y>%=>��8��`�>�����?��V>�0I��G��q<�L>���F��UOؾk׾��c�����%>էF�>�2>���=NT�<���=�o=II�=<���
=���=�9�=��=���=e�>c�>`t}?�T����Z��.���T??w[�>��w>&�%��׃?mD>���ȿ/���`�?Й @��?6?L�M���>������>�k<<����Q
>�X<�A��-�7>{�?D0W�	a��q�����?E8�?��P?�ڏ�gڿK�>N�7>d)>��R�;�1���\���b��tZ��!?BI;�Q̾.�>��=N1߾<�ƾBZ.=Ǆ6>�Ob=i�fX\�wؙ=�{�<=��k=؉>,�C>�x�= �����=��I=���=U�O>	���ޔ7�N*,�&�3=��=?�b>&>��>��?�a0?�Zd?�N�>Q�m�uϾ�*��g��>X��=G�>V��='�B>��>�7?��D?��K?Wa�>�%�=^�>%�>c�,�ܟm��^�6����ʭ<���?�܆?pǸ>�cJ< �A���|5>�R�ý�y?�N1?�N?���>�	
�V�-8��(�W�=�F4�Ŭ5��)��U&���/�O�<OH=T(>n�>�8�>�>7uz>��>��=�V�>vKA>�����>�W����=�=CR>q��=g�s<�;�=�}6�����P��� �#��/N=���z�=��=g��=�N�>ȹ%=Ao�>��=���d�7>Oc���ZY������4�\��x������5�IW�p�>�
�=�8+�N���	?�&h>�Ca>���?��_?��>{�^��.E����f��=擽*��=W�j=[�� �a���h�r�/�@ �>��>��>�>0�l>s,��$?��w=~⾆`5��>}�����2"�8q��@�������i�/�ٺԟD?ZD��$��=~?�I?�ߏ?��>�q�ؾ80>�E���=)�3q�U����?f'?���>C�$�D� H̾n��ܷ>^CI�Y�O�����0���η����>�����о$3�Tg�������B�Tr���>R�O?F�?�4b�RY���UO�x��� ���u?�}g?��>�J?`@?v��qu�q���x�=��n?L��?N=�?�>o�=n��p��>Q�	? ��?�7�?,�q?1�=�
�>�� ;��!>�������=j[>���=�A�=�?k_	?�?	?O|����	�]����4]�m9�<���={��>>B:r>kK�=rEe=�{�=�Wa>1�>�א>e�f>nɡ>���>����]@���
?0�=��[>��7?'�V>�a|>9D��R�=4ڒ<m���]������'�A��}���2=�>|=�-��4�>�п���?�>�Z4���E?�+�F�=��>d��>ȴO����>��>{,�>���>�>|aq>�T>�b>R�㾙]>�������C�d�aF٠>�ڟ��lU���#�d���?h��|��Gr��|�A��*�=�P>Ē�?M�=!冿��2�ԂI����>\�?�6h?����-(��!&=���>��>�c�p�������7f��bo�?y��?��w>��>fv]?��?�`�\2���zj�Z�f���=��O_���H��*��a��M���;�B�G?.3n?e�7?5���8>f�?d����Eɠ>�@T��'B�HA����?iڞ�W�s��4;����7#���=��_?��b?}�?����> 5�}-$?w?���?;D?-q�>u��=zi?E��<{-9?@1,?�9?ÈI?"
?��Z>��>Y���3ʽ�T�*���A�ڽ���M���|?�6E,=O�o��b���=��0;fM�9��ݼ��{������w<���<u�==��=z��>��]?Z�>?��>��7?Y�h�8��Ю��(/?5�9=����L��DТ���n�> �j?h��?i_Z?"Kd>~�A���B��>�=�>p&>\>gV�>d��vE���=wP>�[>�ĥ=��M�aց���	�\���:�<�>��>�J|>�:����'>ࣣ�Smz���d>R��=��q�S�kH�� 2��yw�Z��>ۧK?a�?���=�t��N���hf��?)?�F<?>\M?(#�?¥�=i�۾��9��WJ��5���>���<y���¢�b=���-;�sQ�7�As>�,���D��zwr>�}�(#���q�G�c���=G1��u=���S־�
}� ��=B>���}�#��6���;���*P?���=�"��[oZ��>���4>��>���>_�Z�"����B��@��Y��=~��>�]9>Cܦ�������H��Y�|u�>A~D?m[`?�j�?���s���C�>A��O梾���p?{7�>�?�*>>C��=��������d��E����>Q�>����G�����������$��m�>�M?�>P�?�LR?��?�'`?��*?;�?���>
Դ�雸��>&?Q��?��=w�ԽT���8��F��>�)?y�B�N��>��?��?	�&?��Q?5�?3�> � ��L@���>vU�>U�W�\��*`>#�J?���>95Y?}؃?��=>��5�&梾���d]�=�	>��2?/#?��?͢�>���>������=:��> c?�1�?��o?�}�=�?�2>"��>�l�=ߦ�>��>�?�@O?��s?��J?fr�>/��<�>��wf��o�r���M����;̓H<��x=����t�=���!�<�5�;G��s����c��C� d���
�;�g�>�]s>4���/S2>�ľ�����@>4���㋜��犾�i:�HJ�=�5�>��?֫�>��"�a �=�^�>�-�>�����(?�?��?�9;X�b�5�۾l�L��ð>APA?Y��=4m�Ŷ����u��g=��m?��^?c�U� �����s?;�~?�R˾�v��*��CF���Z�)�?�?矗�pĤ>g�?�En?W?H��S�v�����A�L����r'>�j�>�5>���s�-��>�^b?(??������>¨����b۾OS&?0'�?���?��?��>����t1���>о����ν[?��?�Ȿ(�?�i=6��S���d�P���Ծ�%��h���	&��g7��B����!@�S ���=��?%p�?��p?a�c?����\@m�,9l�4dz��V���5��V�ղO��Bh�_�9�L�b���� �����R�v��=��U�0�K����?��,?� 5��h�>ob���Ӿʓ;W@�>��5�<s�=x{����=��=?�?`N��h��h� ?_��>��>֊R?�d�0�E�_'���%�uW�G'�=Ź�>��>� �>��=��@��+�f�A���b	��w�s>}z`?��K?�Tn?V\�²/��j���
!��n޼���,�L>�2>P�>R�O�$|��%�g+=��r�}�@Q��l���gj=�x/?��>v}�>(�?Lr	?�� ᰾l}���0��s<T��>�h?��>$�>.����!��J�>�HS?\�*?�s?���]� �N�r�U';�~x>�>�E=>���=q$޽Z�f�oX��ds��M+���L>�׊?��|��P��FA�>{FE?�{�=�3���4�>�R�<�t�� ���`ܾL�U>��*?v1M��I[>�%���(�A��#\Z��6)?"K?�w��q*�`>P
"?��>R�>}L�?�ԛ>�>þ �<9��?�^?P2J?�A?6��>�=�D��i�Ƚ�0'��t.=˞�>�iZ>]9m=��=.�ڂ\�9��K�F=�e�=�Ѽiչ�� <$��ZRF<���<�5><	ʿ��=�a����%�=�e��$D��c�[�#���.[�H:U�B�W��fR���㽢��;�J`��@y�r����޽�N�?���?^���{������Q�R��W�}�>Hז�O6w�J}Ⱦ���g���})��t�_(�Z7Z��V�6 (��V&?���8?ǿ�;��oo��r?�J%?�!y?C�����?9���>\G�<��Q�����]!Ͽ`���z^?(��>7[��o��}�>�(�>9�M>Ԯ\>�ل�v_��fB
=�k?jT-?a�>��}���ȿ�.��*E�<���?�@�}A?.�(����t�U=���>p�	?��?>KC1��F�&����X�>�;�?���?��M=��W�� 
�"{e?z�<��F��}߻w��=Qm�==`���pJ>A�>}��lA�jlܽ�4>��>*("����\o^�}��<V�]>R�ս�����?�4A�|9q�9� �~V����u>h?�Qe>����?k?�h=���s�q�з8?�.@��?�_;?�����v�>�ݾs�7?��7?)��>=SE�'������=�h=����,}��#��������>$G�=�,��� ��P���e<CY�=�� ��&ƿ�)%��*�N��<ZLx��mE�8gݽ�д��:z�����^<U�/.ѽʊ�=���=�L>�z�>4�E>��L>TdW?��m?�5�>B�=:!��>�������1��F��#���܇��������j�־�~	���];�a����<�Q��=�S������q"���a�u8>�M�-?I�>��̾A�K�e��;~Eɾ�S���=�j����Cξ��1�яi�o
�?��F?����YX�	��뼙œ��9W?1�<�������=�ɼ��<s �>c��=,��3	4�
�Q� 2?n�!?�¾�3��@V>�,�ğ�;��*?�[�>y�'<�ֶ>~~*?x���0ģ�~�d>�>[�>%��>?è=������K%?��b?����;9���GZ>��������O�9���=�[�<|}</�5>�lb=�����Y��R��)�q=�(W?~��>��)��ja��h���X==��x?��?.�>p{k?��B?�֤<h��w�S����aw=��W?&*i?��>O���	о;���E�5?գe?U�N>�bh�%��>�.�[U��$? �n?*_?�}��(w}�|��k���n6?_u?�O�ޒ�����(e��q�>&��>i��>_T:���>d??���*ܗ�"���<0����?�@��?��<�t����=���>�$�>Ǔ-�AI����;�PqϾ�2=@S�>y�$x�S)����=:?HZ�?:�?�K���*���$�=L���p�?Gۇ?�&��ư�;�b�j�9W �*�<�m�=����R-�e��<6��,ľ�H��k��Vm��␅>=�@�cڽ4��>��4�P�ῠ�Ͽ�J����о���??��>��j���p�i�ݚs��=D���D����F�>��>x𔽳
����{��p;�l�����>�H�$��>��S�&��ř���`5<��>%��>x��>OJ��rݽ��Ǚ?�D��?ο骞������X?�h�?�m�?�k?�+:<��v��{� ���'G? �s?nZ?<�%��O]���7�ӻj?(X���S`���4��JE��T>*"3?G�>��-�u}=�>؆�>�Y>C%/���Ŀsٶ�������?]��?Ol꾬��>_��?�t+?e��7���p����*���'�@=A?W2>y���m�!��5=��ے�1�
?q�0?�N�k'�]�_?*�a�M�p���-���ƽ�ۡ>��0�f\�CN������Xe����@y����?N^�?j�?ĵ�� #�e6%?�>j����8Ǿw�<���>�(�>*N>4H_���u>����:��h	>���?�~�?Rj?���������U>�}?ƍ�>�р?+ơ=3��>mw~>�@��f�׽�k>:�=�3�l��>��Y?v�?��9>v�y��04���.���O��#��(C�-b9>&�t?��T?6(�>��=��ཻ2���}<�ٗ�����,�s�<�e���D{>��>N!�=\P��kľ8W?��TlԿ�*���F�
�"?�e>K�?�K�UG<���Y?(�q>���&��ZV��yp��Ҭ?o�?��
?I�о�����	>��>�Ɏ>R��.ഽ�Hb�{)>�"??/��:����v�S��>v��?�@���?�j�ur?貳�{�0�u���`�'��,=/?0k���]�>h/�>�$�=h�{�$x���j��>K1�?��?��?Guq?�F�D�`���,{�>Y{�?�C?X/���¾��=^#?��	��A��@1�C�`?��@�@ΏQ?�ؠ���ۿ�����ϓ���{m�=a3�=���=�ͼ��=)*};@���馉��ZF>:E�>:�P>OM:>'�U>�uC>��L>�i����B͕�^���y&0��������;���i��Ur�f{��瓾�ԥ�]���8��f���z��)������>4�L?y�C?e�O?$,?�lɽ�C�LՌ�|1�>x#�������> �J? %P?�3+?���fu���#`�u���V�o����>$�	>�%�>���>B�>g���LO�>�0`>W�!>���=�	ɽy�^<��1���>oC�>�5�>z��>�b4>}�M>���ƶ�}fq���m�ޫ�=꽝?�䪾��B����PY��ǯ����=W2+?�q�=g���v0ο\���+P?8�M����؃�FZ�=")?��O?�w;>}���E�<��=�����t��Ԧ=�����s��O2��x>��?�Ie>�ԅ>E-:���A�dAV�̩�v�>Ud6?�����54��v���F���ؾU�B>�|�>�.��m�$�!>���qu�)�L�{�=��=?ou?�`ĽkF��˼y��Α��5>�|>���<�ӭ=<�5>W�.۽��V��$�<���=�]q>MP?r'>k|�=�Ф>�G��|O�t��>�~C>��*>^A?u$?s��/���̃�I�+�4%x>�b�>OL>>�H�-��=o�>�yg>�����W�Z�=��`T>nɇ�$^���s�*w=G����y�=
׍=Wj����=���*=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿdf�>p�aY�����5�u��b#=���>69H?�[��oO�]>��u
?�?+e�T���?�ȿ�{v����>��?D��?h�m�$@��@����>6��?�]Y?Yji>6_۾�YZ�c��>��@?;R?2�>�:���'��?��?Q��?4[>n��?Ã?�x�>CH���W2�FT������&�3|T��ٹ=�>�➾A�H�����#���f�q�/�����>�S=摬>Q����̾h-�=Q���dǾ�/�=;m�>��%> ��>�"�>���>���>Rd�>GP�~��ם��l���!_?���?�W�<o���=1w�>���=Ƹ(?[�W?��9�6�7�>��k?��?�J?K�B>�D�fW����Ͽ� ѾU���B=�=�?b�?u�2�p$�� ��Wv��b[�>\��>�'t��l���ܯ��O���nO>��2?���>~��=ã&?1�!?�v�>�>�N������R�?\��>��>�ł?�N!?E鯾�^$�t܋�⮱�s����Z>�{?T)?��>m�������6�
�˭�<k�=R<�?瓀?D�1�@?^n�?�)?�o?��>��m8 �6�4=�j�>O�!?���2�A�Sd&�K�2�?�f?���>-���UֽbQټ����S���?]&\?�2&?���9a�\7þ��<��"��c����;��B�ȹ>R�>Ó��:��=�&>v��=�zm��;6�F�k<	��=p��>v��=�47��Y��A2?n%;�j����">�?���rM�)�>���=]��U��?Ӿ����X��KK��� ���?Ɲ�?P*�?��Żlq�G;?m��?i;*?s�?�ٳ�ӳ	�G�ݾQ,���Ͼ�"��HQ>]�>C��(y>��㯿M���82����~����&��>�>b�
?3{ ?���>��>�>�T�0�_>ھ%X�EZ����L�]�L�}88�O�辋��ʷ�ƛa�Isþ}����j}>w�A��s�>9�?*�>�nk>F\�>.��=���>���>���>-��>	X�>>u�d>q=�=�ѽ�KR?u�����'�B��~���~2B?�pd?*2�>i�)�������?φ�?@s�?i?v>�~h��,+�.m?t;�>����p
?�`:=)��G�<�U����+2�� ����>H׽3 :�M�lf�^j
?t/?���P�̾�?׽����f�=ly�?�1?;$���V�OMs�Q�K�^�(���Z��8���!�چo�\斿��cm���%�rǤ=j�&?%L�?#��b����
��	�h��A��}�>i�?��>���>�Uo>1��i��?�mj"����@�>g�f?8܌>e�E?!;?>6B?_?�>_�M>�9��;!?[4�jw�>�?�l??"�2?�U$?O��>��?��H>|<��l���P뾟�?��?XV�>��>w�>Zᾋ�"��t=�b=㌾�☽��ﻕ�ɽ� �N�����=�i�>�X?�����8�����mk>f�7?��>q��>���)-����<��>�
?G�>A �~r�c��V�>���?����=��)>���=ώ��U�Һ'Z�=i�����=�5���y;�3e<s��=N��=�Kt��*���2�:Ϟ�;)n�<)�>L8?�B?��>%Þ�?=��fa�u������>j����)>+?��9���?˓�?;���~�>��?�3�?��;>��>֮�t�@�$X����9�7\�'�=I��>��+??D[?h�r?A%?M*D?�)]>��E��#����+��ڹ/?(1?"z�>���(���竿��3��4?�?O�p�̛<��2��ܳ�U�0�w҂<v���x}��ಿ�-?���E>���=����?���?p�/<�F���B��~~��(����T?�>��>���>�HU��w�X'����>2�2?RBm?���>;pK?	3z?`[?� h>Mr6��$������x<�D>Ow@?��?�؍?�lu?�H�>7(>��.���� �2;$��[���
��!%6=7�Y>���>q�>aӺ>%��=��ٽ�ͽ�SD����=Xog>�W�>s �>���>M�d>�>A;\�G?���>�\�����t뤾\Ń��=�A�u?���?F�+?�T=m����E�MH���I�>Ko�?���?Z4*?~�S����=�ּ�ᶾ��q��$�>�ڹ>.1�>=Ǔ=��F=c>�>+��>�&�a��q8�\OM�J�?�F?`��=��ſ�ts�"�w�ׇ���Vk<����1b��"���}Z�`$�=l>��Fz�)ꤾ��R�����񫑾I�������~%{�� ?�%�=�4�=�&�=}�<ü�!=�EB=f
"<�=��i����<t�E�qbq�Ǘ��Y�ջYN�;aG>=}�D;ݫ����d?ŰJ?��/?�K?�MG>f+=a�Ƚ�)�>�����?��q>��!=����`J�,D��M���v�-u�W�Z�'ǝ�K��=I�c���>�f>F��=&80>s�=�d���π<�OP�~�<'��=�U
>�=�O>8-i=�+$=B�|?�=�U���C+`��O��c�?���>�����׾�$Z?l?�̅��ſ���E�w?��@�j�?Ӿ?��˻Q��>��վ(�=�=>9k(�ή)>��@>Oi�t�>���>����F��m��'�? �@�CV?����+Gȿ�x>��7>p1>��R�Ѐ1�7S\��Xb�hTZ�݂!?_H;��9̾C�>��=�E߾!�ƾ�A.=��6>��b=y��Y\��֙=W7{���;=��k=�щ>��C>��=g�����=�\J=X��=�P>�@���7�`+�AH4=4�=��b>'(&>$��>��?�_0?�Vd?C;�>�n��Ͼ�A��mH�>C�=�G�>QӅ=�hB>���>I�7?��D?�K?���>h��=��>��>��,�=�m��l�'ͧ�*��<J��?+Ά?AӸ>$NQ<{�A���We>��Ž�w?S1?6l?��>�� ��Kܿ�PA������<y��x`"���Ƚ�~��\唾�
>_F�=y�]>�?.|r>���=�A>;sb>��Q>���>}8>k���T=�DؼAx���$=~�-=-k<�)#���<y�=�S��v��.�r\7=~Ĩ<o�:�l����>���>��=��?q�=�⯾���=�T�'P��y�=���&n���n� 勿M�=�W����̻=�kq<S��o^��L)�>�i>T��=���?�y?�YU=jzX�mP���ŵ����):ǽ.��?�=q����X�y	a���Y��?�H�>��>7q�>َx>�o,�Q�?���l=���iI7���>���R�"�,����q�Zե���6i�i��!F?���z+�=1)}?qwG?�l�?K�>����RӾ*�>�톾���<3��l�YᎽ�`?�J"?S<�>��� E�݇��C@u����>�5_��S��#��130��%=�9ξ��>T�������3�_�������rHI��Ӂ�C��>�)b?�k�?�z`�����cA����N��R�>�\V?w��>h��>5� ??vq���f����A=_kv?��?���?i�=*��=��w�M��>�k?ӗ�?dɑ?,n?8���[�>`�=��K>�O���/<��f=��|=�>��
?���>��>%F���Q��^ԾÙ���o�a�����=� �>��>4X�>s��=��9>LB>4�R>(�>��>c�>�C�>2J�>�N��u��Z�	?�v�=�'�>mm-?&�>��*��7���>_����_�@#d��b���r<*�[>��=���<t�ʽ���>�Ͽg(�?�S�>i7�V�>����8T>�,>�\�>�P>�(?�?���>LF�>w<�>/�>WK[>[>~>�?Ӿ%�>c���o!��2C�b}R�ωѾ~�z>y���	&�~������BI�hk���^�ij�;/��~@=��W�<�G�?4i����k�m�)�N�����?3V�>�6?����*�����>[��>��>�O�����qō�6o��
�?���?(܃>�&�>Ka?�6?�m!� w��A�g���h�fD��t��8A��A��~�����қG��V?�n�?��J?��D=�8>5ڝ?�U۾ȿȾ���>���o�@tI����>���p�L�i$���5�uؙ����<b�S?Kn�?;Z?<��Pb�M<<��B?Hx?Y�y?�8�>���>�@y<��x?��<k��>�#?�??�H?��>�?��Ղ(;�뙽�I���y���I���¨��u=�.��&��=��$>���	_�����=���=t�w����0#�b�c���x�-=�&	>��=�K�>x�^?3�>H��>!6?O�!�p�<��R��t�,?���<����@*���P��������=<j?L��?z�^?��d>��@�� 8��V!>�)�>�Z!>�]a>B��>.���g0��z�=�->m�>��=�Xf��苾3	�����Ec'=�+ >��>{u>�=}��u9>M������Īd>�QN��~��\T�hMF�B1��>z��پ>m�J?��?��=fp�4L���d��B/?��<?�K?��~?��=$���;��I��g9����>|"�;�U��6��o��� 9��H<|��>N"��O����J>*$!�+H���{��;T�'+��8�=uN�S<ț����7�y�i��=r�>Iƻ����:�������^
Q?�f>�㧾�^4�v�ܾ�c�=S֒>�r�>,��GL�_�;�����~�=jB�>V=>��*=#���L��$�����>�>?�4d?ȇ?M�p���w�x]2�;C�����/ҽ �?�ȟ>��?��J>L��O���>��b���"�l��>B��>5� � 3<��^ž�"���1����>"�?p	O>S�?�	M?��>��a?�0?��>Gl^>	�Ƚ류���&?$��?f�=��޽>�S���6���D���>�U*?rA��ؕ>z1?��?��'?t�R?/�?^
>a����@��>Ί>��W��0��`>�`K?Z�>��X?�˃?f�A>~"5��ţ��h����=��!>�E3?��#?� ?��>���>˭����=���>�c?�0�?R�o?Pw�=�?^@2>���>m�=�>���>�?VO?+�s?��J?��>���<0C�����js�1�O�y�;�H<��y=J��-?t��^�@��<ݝ�;}B��D�������D�l4��NE�;	_�>K�s>���t�0>(�ľ3P����@>p����Q���ڊ��:��Է=䄀>��?���>*X#���=��>9H�>���8(?
�?f?��";��b���ھy�K���>�B?S��=g�l�L�����u��h=�m?֌^?d�W�"&���ct?7z?�𵾚?�����^�Pp׾(�|?fz?#�j���>��g?��m?S?��=��]�d����jw��3��w>H��>��@��M��Z��>M~?�?�.�>�ɩ>����W3���;��_�3?t�?p�?;�?]^�>��U�kDٿ�Ҿƙ�0�R?O�?yu��D}?gփ;�)���Eھ�N%����������떤��̾�9���`����Kn�=w/?��f?��?��`?!_��mf�W�h��V��ӆ<��e������L�r�@������^�e���-Ҿ`�����=2�y�IE�H-�?��'?7�3�c�>�����e��վ��Q>c���
?�fю=�ʞ��=o�R=�b��=+��ɬ��J?�ò>���>8�=?�D\�Qe=��1�5�8������->I�>���>��>mz�<�J2����qcɾ�ꋾ�L��"�u>�c?�L?��n?� �sr1�#끿)�!��H>�膨�wPB>r�
>��>��X�w ���&���>���r�.����6V	�� =�2?�j�>;�>��?9�?��	�c��Eey��1��2�<U��>�h?A�>a΄>�aԽY �ݹ>�mQ?��?�>�>M����7�k�d�a�����>*4�>� ?��R>�ܱ�`�M�u��Rc��U�#��l�=�%d?�x��2�{�k>k�??#H�=W%�;+?��K���Y�	��V��2*�=N!?��R=y�=����2��`��t�
�W9+?54?�Ǒ��Q)�@#�>QX'?�y�>4v�>�q�?�ҩ>������-=|�? e?�NP?e�5?d��>)�<��5�XHF��q�=}Z�>3Kl>�9>=�[�=���� `�Z2�n>+=��>����xٮ���<槼,#�;T�<.�I>Qr�|�Y�A?��T$���v���ƥ������~bQ��že�����y���Z��=��g���y�����x����?��?�	�&�Ⱦ����ʁ�qT����y>_\��ʷ������Z�i�7���qȭ��?��s����I��p�f����?�Jd��Uƿ�i��~1��&?8c3?�Uk?���I���0�j�H>��\=� ���-7��(GͿ����e?��>��۾Ӆ��˼>�>���>m�>=����I��0���R�?�2?3��>�}O�f4п5J��.=�'�?o�	@�|A?��(� ��kV=���>z�	?�?>�U1�KI�����cU�>I<�?���?��M=�W���	�Ve?ph<��F���ݻ��=�A�=�W=���:�J>�S�>Ȃ�]TA�xBܽ��4>aۅ>�x"����z�^����<��]>��ս66��5Մ?,{\��f���/��T��U>��T?�*�>Q:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�߅�=s6�ꉤ�{���&V�{��=[��>c�>,������O��I��U��=WN��'˿��"�w���2=�t;;<��ƹ��ӄ�#l(��E���-g�LM۽s�|=��>��W>c�>!�E>�"a> [?�r?�ڣ>q��=:� �y����W����D��듾C�1�`˅����{���=ᾍ�ھ7��Ef�9���о�=�S#�=)S�DА���!�N2c�[�D���-?��>�i˾`�M�0�;*ʾJ���l�u�����̾4!2���n���?�B?����11V��6����#���(�V?�����������=������=���>�m�=�����3�G�S��x0?�P?8b��Q���+>���t=db+?Y�?��b<���> |%?��)�T�c�\>_D3>e��>�8�>�>���hܽ��?t�T?�]�*Y�>��Q8z�cZ^=��>I14�.伏�[>zP�<������Z�����d�<e(W?���>"�)����a�����Q==��x?�?}.�>v{k?��B?�Ѥ<h����S����cw=��W?*i?u�>?����	о����ҿ5?��e?��N>�bh�i����.�CU��$?�n?�^?|}��3w}��������n6?�{p?RfX�5���d�7��u��>�_
?�+�>�'`�q�>hZ?	+�!8����������r�?ˏ@���?�F=�}(<>�j��?q�*?�㪾 p���[�ORc�4���-?n���l����:���)�4??��|?���>u�����?��=},���P�?��?薪�-md<?��0l�߱�����<��=�+�I$����8�H�ƾ��
�ݪ���𿼦��>R@�Y��6�>k8�R(⿒SϿ)��0%о�r���?:�>Yxɽa�����j��u��G���H�A����M�>��>ܲ��p���L�{��q;��#����>���	�>�S��&��ǚ��ӓ5<��>��>5��>�+���罾6ř?�c��@οY���ם�u�X?4h�?�n�?q?�9<��v��{����L.G?ɉs?oZ?�o%�>]���7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�d�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?S�>	�?Q�=�>�C�=�[����$�z">w�=��;��?��M?Ǖ�>%v�=��7�/�);F�9R�S'���C���>��a?��L?��b>)B���4�s� ���ͽ�1���>	?�h*��߽2c5><�=>��>v�D���Ҿ�?Y���ۿO��ސ��w	x?��>�=�>��޾E���=l��?@+�>��A:������r<���?v��?��
?͹�迨���=�3�>��>n����r�<��w���.>ʪA?Q��l��Ő��f��>PF�?u@)��?dHl�%e?	����8��������)�`�9�2>�-?�p�y�U>F]?n:N>��u�/l���`m�+R�>]a�?��?Ĥ�>[�g?��r��'-����=��>��8?�V�>���=�����;>�?)?�ȟ�ޙ�IE|?�u
@�a@�8a?˧�֮�MT��3暾�t��=�>��=k��=z�=�.>gs�=$#ҽ[$����>Ev�>TT�>��Y>�z>5S2>�fU>2K��sp�aN���@����@�fG����g�Ͻ"��[������R�о[ĵ��ݪ�)<ƽX��!#��� ��s���=>�=?;WE?sY?z/?�\�=�ֿ=�����i>��)�C�>��>H	S?�u?��P?B��=�ީ�#}e�^m��P�������?s)�>��>���>�L>�`!=�R�>B4[>,v>�|S=.�-�C�����;��X>�ԅ>a��>�&�>�@4>Rt>ƴ�����j���}�޼����?����yI�MQ��U�������B��=�.?>ݢ��q5п 쭿��G?����+��+T&��>U0?W�V?r�>N��� 0C���>�q��c�+��=�U �a�j�f�)��Q>��?�#>Pi>nB�\A�+g��"Ͼ�ޓ>��#?����`.���~��}<�=/ƾT<>R��>��<f��r���Q���Ir(���=+87?�z?XXͽϭ��<>��+��ǻh>�Uw>p�l=�\;>��u>���[����,���Ƽ�5�=�M�>*�?�$>���=ю�>��h�M����>��E>�'>�r@?�&$?��r����C��/�/�+�u>G��>Q׀>m
>�[H�z �=�X�>ܢe>٬�L����6�s�A�c�R>�:}�m`�Ks��z=�z��\�=�m�=���B�v3=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ>F�>L�������������%�=�A?k,?"�������=��"?1#?�+��b���`п�y����>\!�?��?)�_�҂��X�=���>�u�?��Q?�X�=�紾g4k�S�>6XD?IC?���>��?�s�X���$?���?���?c�A>��?�A{?K��>�2˼�d4�����6����ϼ�c����z>�x�=���<9����� ��>uo�Ml�JC�>�Vk=�Ԩ>|'��+���$�=��������)=(�>
�>�3>3�>\�>(��>1��> }���U�Mה����`?9A�?bd����I�=9��>���<P�?�.V?��\>��z�UW�>+�}?jr�?�!�?��>����(��򧻿���������K>E� ?�N?�
ɽ��%>�A��%�����>�r�>u�=���]�u��.׽�<>B�?2��>���=�/"?�[%?�U�>���>��C�S0��"�B����>���>Q�?���??{��V���M��14���	m�Y��=U�?�^#?\�>�D���ܡ�9Ƚ"
��8 <��P�?T�_?%�>"?�E�?��'?��3?�=�>@������"�ֽ�ey>��!?��O�A�nY&������?�T?e�>5���l�ս�Y׼2���F���?�6\?MA&?*��4a��þD�<�:#��d]����;`�C�!�>�>z����´=�?>�Ӱ=�cm�6�N�l<ח�=O��>�p�= 7������q,?@ ��"觾9Q>��~��J@�.h>�y>
�Ix?�{ս3ⅿ{����읿�[5�8�?�z�?7�?]�9�j��??t�?'�#?��>�ꪾ���n��s����f����&������?�7=���}ߤ�����k��>j,���0�g�>B��>��?߲?�>/�>�[^����J-�����bed��g'�3bA��;��z�溑��ƽ�?�"_��Ju���И>�(���>Vj?�zb>,6g>��>jR�[8�>�x>�@>�x�>Ǣ7>�'>�!
>�j=��J��KR?#���]�'�_������3B?8qd?c.�>:i�{���5����?҆�?�s�?{Cv>�}h�r,+��l?�<�>���+p
?9n:=���QH�<�U��`��
*���c��>�K׽�:��M��if�dj
?�/?m��'�̾8׽`W��]p=Q�?j)?�)�"�Q��o��W��	S�����1h�]Q��"�$�+fp�돿�r��1)��E�(���,=7�*?�?��MgS��zk��#?��cg>�,�>!�>��>*�I>+�	��b1�?�]�5'�Q̓���>�7{?�>ؖ<?��*?u\<?qa\?�߷>��>�Fʾ�i�>�d=�L�>��?F�L?ƪG?��H?��?+�?�7�=��!������/ݾ�'?D&?�?���>�ֵ>Q+���ѾL��y��H~6�+��9u�=ӇT=C�'�N��?a�<��c>�W?W��Ҩ8������k>��7?8��>���>����"��t.�<��>Q�
?BG�>����]zr��`��O�>m��?u��N=��)>��=jǅ��ֺ9<�=}���@�=�|���;��<���=��=�*t������~�:,d�;�ï<�p�>�#?_��>�&�>�&��	��[��ν52�>p+H>ɢ}<���n*r�!�y�^8Z�r�>�w�?���?�"�ϐ�=o�=��+\�ew-�fǽ�}�=��.?d�
?n�T?TԜ?^�H?��?�+>��i��h1��M����Q ?m!,?��>�����ʾ��։3�ܝ?d[?�<a�	���;)�ِ¾��Խͱ>�[/�^/~����CD�򅻸��0��2��?꿝?>A�O�6��x�ֿ���[��w�C?"�>'Y�>��>W�)�y�g�q%��1;>���>uR?D�>��O? 1{?M�[?lV>�78�v��ə�H#���">j@?��?�?�y?��>��>*���3������J
��Te���zX=�yY>�G�>���>��>���=>Ƚ�}���i>����=Aa> ��>TZ�>3��>/w>g��<q�G?-��>]�� ��+줾�Ń��=��u?囐?��+?PV=E��!�E��G���I�>Oo�?���?%4*?�S�1��=��ּⶾF�q��$�>�ڹ>�1�>ʓ=6zF=�b>!�>'��>�(�a��q8�SM�;�?kF?�=��ĿpTr��p� ȕ��<�5��A�_��K��!b��3�= ���(�ٰ���]��Ơ���������B���w�}�=-�>��=�>
��=�1�<��ݼ�o�<86=�g<�y=�{��{j<�@5�D=�$f���8��q+<<�)=��>��c˾�}?��H?e|+?�C?Ƃx>)�>��1���>򢋽��?�8S>��Y��]��1�=�q먾�ϔ��׾�A׾uCc�i��n�>vN�97>�4>@�=�0�<�i�=�!y=��=6�
�}�=�7�=�=�=���=�>�>�6w?I���"����2Q�"m罂�:?O:�>7��=��ƾv@?%�>>�1������d��,?���?U�?V�?3qi��b�>����Ȏ�嗐=�Μ��22>���=��2����>��J>C��QM���u��:3�?f�@	�??[ዿ}�Ͽ�a/>v6> >O�R���1��^���c��>Y��`!?�!;�kZ̾h6�>&z�=/߾6yƾ�5/=�6>�]_=��%~\���=7�x�g�>=�Im=*��>KD>��=-D���ڷ=��L=��=�Q>�`{���<�$+��5=�I�=M�b>F'>Ï�>R�?3d0?�Ud?�5�>un�H(Ͼ�?��$P�>u(�==F�>�ʅ=�gB>ŋ�>	�7?��D?[�K?8��>=��=��>��>�,�2�m��u徉ͧ�ݰ�<���?�̆?�Ҹ>q�S<�sA�B���d>� AŽ*s?�M1?�g?��>���0꿞� ��A&���z�izO��J�<����'��ޤ�5W,�y���9��=Ҁ�>���>���>ަs>��>h5i>H�>_�R>s��#�;��/�<�D�=
^��	ġ���F�c��;�2=�0:�� ����Ѽ$��;cq�;lf������i�=���>��=h�>�)=�aȾ;,>�2�ÐT�=�Y=�֧��tW��a�-u��b>/��@���?>�q_> ������*?�w�>�>��?�c`?�8>9���4`�i���g���_�BX�=��">����S�8i�~�H��پm��>�ߎ>l�>�l>�
,�$?�{�w=��Gc5�x�>fz����� ��8q��?������i��^պA�D?E��B��=^ ~?��I?X�?���>����z�ؾ,0>IP����=��"q�R����?�'?���>��H�D�nH̾���߷>�?I�#�O���O�0����Vͷ����>�����оq$3��g������ݍB��Lr�K��>�O?��?�9b��W��3UO�����(��xq?�|g?7�>�J?�@?2&��z�r��Xw�= �n?ĳ�?S=�?C>،�=M#���$�>�&	?���?��?�qs?b\?��e�>ij�;�� ><똽���=�}>0�=o�=j?�
?�
?PB����	������7^��@�</ơ=���>1H�>�s>]��=\�h=n٢=\>�۞>1��>i�d>m��>f6�>�O��V��;�
?�>p��>q�(?q��>��U>1�B�}�=�o�ټ��s����P��v=7�P=`>��l��>e�ǿ�?�?��b>�K)�:?��ž(e�<Ե����>L����M�>��>*L�>+��>��>�{�=إ >8�4>U�۾t0>���w�(�'�T��S��R��	�p>~�������
�����8�"�f���i��^CZ�$����F���<ȼ�?����/_�y�+��O5?���>�)?�h��
ߓ��L>�?d%�>Ө��hA��y�������?0�?2�$>Ǆ>��i? )?8�-��g��to��>{�"D�����M��|���c������<a���o?�2�?P?&���>B��?6����Pξy��>�M���P�������>�p��о�̽��0��?�s���c>lp?BЕ?t_@?'\��d�K<�-�=�`C?��K?gB�?E�1?R�>
>��PmD?���>U�?�g4?ʎG?/F?#�!?-qE>��<�oo���<��׽�7���ʖ�iW���p�,�%<���=��ۼ6���|=��>ڤ\=Ԉ�W8��#�c�lI��=ê=6>��=��>��T?��?�*�>I|@?Ϥ0�{�[����ZM*?��,��1��Ҿ����J��<��t?�.�?��h?X)9=�n�;=O��ǝ=�?b>�)�=V�(>�P�>()ɽB)M�+D>:T�=��=�2>�*=�]e���r��~TƼ%F>���>�2|>���u�'>�z���+z�B�d>��Q��ʺ�q�S���G�"�1�Ҁv�w[�>L�K?�?�=�_龩4��If��.)?�]<?ZOM?��?�=��۾�9�P�J��?���>Z{�<�������w#����:��^�:��s>T0��<࠾�ր>������䁿�9�Ȧ¾���;�w�Q�=�t�����߂R����=�'>=�������"<����S?�� >�dƾ��W�`����>ݎ�>�<�>}��u���C�٪��ߟ�;7ܽ>�>��v����tI�������>7�B?Up`?�ք?�W��q��27��� �f���FK9��z? T�>�'
?��F>��+=d���V����`�ѹ9���>tg�>5;��sH������WﾞP*��K�>,|?��>�]?�R?�?w�j?��+?�7�>	��>�&���ܸ��=&?䇃?6 �=�Խf�T��9��F�M��>��)?Q�B�ɗ>$�?�?��&?��Q?٫?k�>X� ��@@���>PS�>^�W��`����_>�J?��>,Y?�҃?I�=>y}5�l̢�����Z��=,6>b�2?%0#?��?Ǭ�>l��>%���Y�=�t�>�c?���?��n?L��=gG?��8>�e�>�ի=���>e��>�*?�[N?�Yr?sI?��>/�<j���Ud��li��G�.�;MG2<-Wl=���.ri�x��*z�<��:;4��芼<k꼱�E�!.���X1<�`�>}�s>�����0>�ľ#T��V�@>!��mK���֊�\�:���=��>� ?���>�Z#�C��=R��>�@�>����3(?F�?�?e'%;�b�; ۾��K�S�>�B?]��=A�l������u�-�g=Q�m?��^?єW����\m?<�m?J<����n����(x>��(=���?���>�~��QC>m[[?��i?��"?�]�|����"���h��r5>g*>m>!���T%�1VU>�DC?ɥ�>l��>4d=ܪ��f�����.�>�I?���?��k?Їj>+�V�x¿	��p��Xh?%�>b5���1?�x���۾�+��$�ƴƾ�x���귾����@빾(���o�ʺ�OOs=�?Uzt?# r?Q�b?
����k��~[�?��o�V��
�i�
�m�E�n�I���8��pg�"����,3����=?�^��G�֧�?��%?[
�)
?�����z��fԾ��4>D����wａjl=����Rt<�~x=��K���9��ɼ���#?~�>{P�>�>?��f��~:��30�|�C�Y	��*>��>���>��>T#Ժ��6�祹�p���'�y�;a���u>��b?�K?�pn?L���	1�5��@0!�*�!�rߧ�R?A>>>-�>bV�|��L�%�,T>��r���+ꏾ8�	��u=�;2?2�~>�͜>�*�?��?�;	��>��'hw��1�<g��>jti?{��>v��>�C̽ 1!�"9�>_�d?��>�s
?�u��#�F�od��,�����>-�>&��>7�[����b��&����i�N�0��R�=8R}?�o��rM�	Rc>�4o?}�4�Z���T?���P�q�����Ťg��BK>��??�>gV�=-���xL�>τ�P�)M)?0?J����X*��J~>�!"?�}�>�9�>��?�[�>�8þ���9�?��^?�ZJ?�&A?G��>��=�%��h�ƽ�U'�kW+=~��>�K[>��l=���=���]���>D="-�=�dѼ���{ 
<����sM</$�<614>#�Ͽ��<����dJ0���	�i�?	�����<V��(�<yn���Z��C�սT���5v�<���l\a�Q0z���?z @�;�Y�����e�*�Ͼ=�>�	f����=2J��$�žl���ݾ�����i*�M�E��t�|z���? ���|�ɿ�U���. ���?�9?��F?�	 ����l�[�{/>t�<=	����v �ݵ��=����精 d?j0�>�����Շ�Pb�>'P^>Z}>�d>N�z���� ��=�{?��J?�|�>Ԝ���տ󀺿$�=k��?c�@jbA?�)�y;쾷�]=��>T�	?x�?>&�0����Σ�����>0K�?S�?�"U=��V����\e?�(�;��F�����=��=|e=C��fJ>J��>
]�ޡC�"vؽC4>cG�>��'��j��G_�u��<� ]>��սuT���Ԅ?x\�f���/�^S��]O>s�T?6,�>P�=��,?8H��}Ͽ˳\�O&a?|/�?ݧ�?��(?�Ͽ��֚>j�ܾ��M?�H6?���>�e&��t��p�=��2��'���*V�4��=���>r�>�,���ؓO�-˙����=��;�ſ��!�p����W=	ݢ<e����9��|-���∽xg��-|V��n���y�=2�>ʫv>}e>I�H>vj>�s]?�Pw?��>j=�6�t&�����jǪ<��w�w9Ƚ�m~�O�C�H2~��h�Q��0��a��F����ɾl�:�H�=��U�E_���+��	\���<�%?�� >�M��"�P�;o��|��Dv�����E����W˾��3���r���?/J?/����V��	�Ҩż�Э���P?68��@#�J����`�=q�>����<��>ʄG=�澞�6�W�T��u0?�\?����5^��S(*>�� �6�=^�+?��?�Z<�&�>�L%?��*��0�#d[>i�3>֣>��>�:	>���V۽q�?ĈT?��������ڐ>�c����z�ca=�1>G:5����#�[>�z�<��O�U��J��G[�<3|W?=��>j�!�u����s;����==�Mz?�	?��>r�r?�eE?"�=���5V����^;w�Q?.n?(>�HK��Rᾭn����6?�|q?{i~>�5X�Û���3�����0?_o?X�?�x�;p�w����/��{6?�To?��'��a��vU��1����?���>��?78��;�>x�o?E��=T���~�Ŀ8���?��@�<�?�eL=K���=К�>С�>`��;\���_�~�?�ԾѧM�ɫ>o�w��蚿OG_�A�=�\W?2�?U��>t�L1��:>����r\�?=\�?����I�=���'p��	���ݼ�>�#;��i��������=�O&��&��WǛ�ϙ3����>�@��˽s��>���:�ʿ7����nξ`2���?o��>l�/�.��44a���e�of:�U4�d_r���>�s>YN�� ����{��X;�
���v�>e� �>�>e�S��鵾���6bB<��>�r�>�V�>���������?N���[3οN��į�R�X?�H�?U�?�#?i�E<C�u��z����oG?I�s?�Z?�� �=p\���;���j?�]���U`�F�4�0IE��U>Y#3?�A�>$�-�\�|=�>���>�g>�#/�r�Ŀ�ٶ��������?��?�n�5��>��?xs+?]i��7��>\���*��P-�=A?�2>K���θ!�i1=�Ԓ�`�
?;0?�t��,�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�U�>fr�?��=7 �>���=����gZ���(>�< >M�5�<�?ԱH?�`�>`��=��1���.�D�D���U�"q�dTC�$K�>��c?��F?��e>l«���p��e$����	(�90L��N8��@Z�N����&&>"�:>�`>x{9��˾
�?tҾW{ٿ����Iɾ?@	�>2��>�	�̈Ͻ愴�u2_?ֿw>�<;�峿����bT�A�?3b�?6�?�������F|6>�4�>�C�>�ᗾ�X>��þ�Ն>~S?M���ٞ���!��s�>���?^F@>7�?��U���?�\ʾ�5��Iiw�60��>�<X�Y=��P?ѯ#�(<�>hh�>��>ۙe�����kRn��U�> ��?R>�?؂?�Jc?�Mt��Y%�C��=� ?g�q?L��>K�8>���q�>.8?�����撿s�辪�j?��@�@��n?�L��Ǌ޿����*2��f{���K>s�=z��=��&���]=X�#=�^���,"���+>X@�>�_>��>[_>-�0>��>|j��"��՗�#����:�������镾i��
�,�/� �����I�}��?���A��<߽N0�(3�Zs �ٍ>�O?h'H?.�U?���>&�ʻ>����/C�>>����a>z܂>�b@?+�^?z(?6j�����{�g�\�����d�u��>� n=���>� ?���>\�=�{��>�k>ֱU>��>�O>%�>Q�=�2f>���>$�?ȱ�>�W+>��=>����<Ե�{�v�/j[�߀u��1�?ޅ���h@�?i��N���g���(Ҡ=�z)? \�=�Î�[�οƓ����I?��h�
�/��N�>�Y(?@UT?�R.>r1���1齼��=��D��E��*��=!!(�J����-���F>�%?�h>ʨv> m3�i8���P������>8�6?y��J�9�>v��H�3�۾P>��>�P�l��u��`��j�,�x=�;:?W&?�筽),��a3v�I��S�Q>A�\>1�=��=�HM>��_��ǽ?�F���7=y��=8]>�S?��)>@ �=�t�>o����O�dk�>�B>�C,><3@?�"%?���ᓽ�o����+���v>���>�{�>��>ƞH�v��=���>�Sb>�� �v��<9��i@�N�T>�w��"_�@p��kt=�L��a�=���=�H �]�<���*=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�0�>�U���)���q����y�}�=_��>qPB?)���H���R��P
?�?�I��V��Z�ʿ��u�*��> ��?�3�?��j�Uޘ��:���>A5�?�bR?[�h>?�ܾ̺E�k�>�A?O?�-�>ׅ�"�%��/?j��?M��?DI>�w�?4�s?��>��y���/�$���Ҽ��2Zu=�=;�ǎ>�>C¿��4F�l��Kk����j�q���]c>K�$=�Ը>�߽C¼�$(�=�#��'ר��OV�_�>h�n> �I>��>� ?�>�=�>�=2G���l��p�����[?v�?-��dJ��D
�D�=�t#>��R?��??^���<0���>�^?��?b�}?RP>>�b$�Ћ��7g����ܾ
!p�X0>�0?��?�]����=TŮ�h���(�>��>��?��hz���W� �����>r>?��I>�H<�� ?�}*?��>���>��g�)鮿��7�x��>Q��>٥?��?�?�T�hBܾ�皿�|���4�k�>���?�(!?�>b���A߰��{Ͻ�?��\N�⡞?FR�?M >:H?ø�?�U?��J?!��>²����T�V�齋>{="?���JA�W�&��w�� 	?!?;��>a��/ڽ�t�����h����;?_G\?�%?sk�^Wa�}�¾��<��7��;���F0<Y�C��C>�S>}����A�=NR>�ç=�l�s�6�;Uu<�1�=�G�>C}�=�66�] ���(?|l=\���eJ��aP��
@��>��>�a��?�˾����K���#���!��?9�?o�?5��?-���$g���.?�ܗ?�?��>I.þ����+���8�B��k��)�=�O?��罣���e��ܞ��hw��3:���??��>P�??z?�=�$�>̂��/���!����-v]������F�g�N��M�����P��Dy�'W��<!���=�>^�Խ�՛>bw?L�>u��>���>ARn���>p��>�>s?ƛ�=�h�<�M�=��}�_$�� S?|��s�&��x쾶Ҵ��WC?��e?n}�>ASY�ZD�����y?��?�
�?�g|>�h��8-�^�?�"�>,�{��K?1=��D���<�v��T�(�y����Fz�>���7��L�:�b�b�?{�?�C]��
ʾ�w���o��!�=gu�?
�.?@J)���Q���e�j�Y�3T���y�@���r������i��V����C넿ʶ&�A+�=�)??�X�	���ȍ���h���F����>P�>�Ď>y�>7�]>_�fB�)�U�+�F&����>d�t?�Ҍ>�QI?�P<?�O?]L?���>e�>L����N�>���;��>�$�>��:?v/?�F0?�?�e)?ŅZ>��������h{ؾ_�?u�?ٛ?�?�?�~��0ջ�����Yl�%�r�9�w�Tw=^q�<�ֽSt��m=�U>�?ܢ�C�8�ۊ���1i>n�7?��>���>2ޏ��΁��6�<���>��
?ɏ>����ۤr�W����>���?R�I�=�1)>���=�.��z���ʜ�=�	��5u�=J�����>��"<i��=�m�=�1���4N:r�;˳l;<��<?�>rH-?]�>��C>r#3��'Ҿ�}�Tr�O��>������<u(�_��bG��������>��?ڠ�?�oB���=e;=�@о}4ɽƹ��ƾw��=.�>��?�v?�_}?��?
�_?�|�=�侖���W������[?�$,?�a�>+���)ľ���Un5��a?lr?�]����v�(�?J�����*a>�"*�,
|�H�����F��_l�nc�a�����?��?���V8�ML�ᙿ����B?�J�>
~�>��>/�+�rZj�E��sA>�]�>�Q?���>�O?H&{?i�[?f�T>'�8���|�������!">��??ב�?��?�y?a��>vk>�(*�fK��=��j8�������SU=��X>�ɒ>�2�>���>��==�ƽ����0>�0ڦ=zd>��>/٥>�.�>�
x>K4�<O�G?A��>L\�����"뤾Ń��=��u?���?_�+?kQ=J��W�E��G���H�>�o�?���?�4*?�S����=��ּ�ⶾ�q��%�>�۹>30�>zÓ=�{F=Gc>�>���>	(��`�r8�%PM�[�?F?Ω�=��ſ��q���p�"�����f<�0�d�D���i�Z�[Ф=8���_�#���֤[�#���k�����ߩ����{����>�)�=zg�=E�=��<+Jɼ���<>�J=%E�<�a=%)p��Xn<G9��HԻ԰������\<:�I=\��'þ�?z?SI?��+?[D?6P>�J>b��mΡ>��p��~?�N>M�������{1�����!��ҩ��YӾ��e� L����>IU���$�=�"=>V��=�;a�>�=X&�=1�N;oD=Ț�=_ �=?#�=���=Ŧ>��>ct?/q��s��lAS��Õ�_�0?3څ>cA>V����E?V�E>˴���T��q���?)��??��?�?��x�]��>؉�M�\=�J=���Y��=�؃=>,����>�>#G;��W���&�*|�?�.�?��E?�]��WO˿�<>z�7>G>f�R�1��\���b�?qZ���!?�C;�F<̾;:�>�?�=C߾��ƾ�.=e�6>Qjb=�l��V\�v
�=�N{� �;=�;l=߉>��C>U]�=@L��߬�=Z�I=���=��O>���A8�>g,�@�3=���=%�b># &>���>�?�^0?~Wd?t:�>��m��Ͼ�4���Q�>�F�=oD�>� �=ڏB>q��>��7?��D?c�K?Ix�>኉=c�>���>M�,���m��c�o����b�<M��?�Ć?�۸>/R<pA����nb>��ŽFt?Q1?�h?C��>y[�@A忠���:�b{>j��=��<;��B=l�b�,ހ��#�q�=�f�>�?��>^�>T>��>Z��>u7D>�;.�{о��o���S<=���=hk�=��˼P����x��2� =�F�=ױ����;$��<�i��$L����U<Fe�=�2�>r�=��>r�Q>��ľ3�_=GW��iZ���4��+žt�Y�8]r��{��A?)��*�|k>�\�>2x�#'����?�>��V>�	�?��i?4U�>��>�\���xW��q��M�=���<Yw����l��pa��^P�̇�˾�>��>mH�>�$n>�+�s4?��e|=���%�5�o��>}��q��v>�	q�T�����%i�&H�ʹD?�#��a��=C3~?�DI?Y��?ߍ�>{⚽14׾`�0>Y����;=��:�p�����*�?<|&?,�>+��ĞD��F̾3
��Rܷ>�@I��O��ˮ0�����ͷ�4��>F�����о#3�|g��0���9�B��Mr���>C�O?�?;b�W��_TO�O��(���n?�~g?0�>K?B?u��+{��s���v�=��n?ɳ�?9=�?�>�a�=�۾��F�>;?Q�?_��?�@o?�b)��s�>��<�&>$؆��
>-)>v�=�J�=Y�>���>���><�a����@)��������c=��=qt�>��s>|6�>X�>���='?�=1R�>��>�Q�>
�>���>�H>�
s��!���?L�A>x\�>T(A?��(>B+�=}r=��<�{=6���^Ľ�U���`�Ծ�<ނ8=�UA�|u���
?$cϿ:�?�>J��70?��̸����X��>�ɳ=�=?�'�>� �>���>�K�>[t[>��>��:>�1;S�.>���L-���L���H�1����{f>�L���n(��s��g�f�?�ȏ��Z���_h�����EC��q���w�?�P½-�h��J��
нj�?q��>=r3?Y����D˽� >��?�}>�"�k��ؑ����fى?��?}9s>E�>x��?_3?��]�<����	������d�'�ڌ��+���9������R������}�|?Ђz?0Qi?�N�C>��?��cuϾ\�>��$�w�*��F���q?�վ�������H�ξz����8�=>�z?7ń?��`?[{�����=��K?(�W?J~�?��?%��>k@��[0?)�>^�
?N�^?�]<?7�&?d�,?(h�=�Հ�:2N�L����e۽xXs��罅��k�C=�c�<X�=-v�9=�����|����������~5��%d�<�����\�=⯟=3��>�!_?��>0�y>�6?��b�E����z�,?r �����u�� \������Ƒ�="�s?T%�?B�b?��1>M�7�~=��Y�=��l>��>��o>�ė>�T�K�$��;�=�F>�o>���=M�A~���:
�Њ������)�+>t~�>6��>6,h���>~ ��Ⱦ��>�J��A���=�j�6���&�Q�ڽOY�>!�N?;E?��<('��"��1j���?�c_?JPQ?��?HCټ����`�,]>���cn�> _�����ס��4:���.=;e>�ES�������>�2�wD
�2���I�6�G���_=P��ye������ƾ_vq��x�=m>�A��l��Oʓ�"��r�N?G�=�q�zz&�F�־7]�=�n�>�n�>��=��w;����ԥ�^��=���>��[>��=�<о�K�����
�>2E?�s_?���?�ڂ��s�]+C�)���]���@aѼ=�?e��>��?QA>�Y�=�a��%H��ad��F��>e�>�n�J�G�\J��:)����$����>;?f>�[?��R?��
?�_?�)?2�?��>ܝ��H����A&?,��?�=��Խ+�T�q 9�F�d��>��)?F�B����>m�?�?6�&?�Q?ѵ?�>#� ��C@����>UY�>|�W�ab�� �_>m�J?���>z=Y?�ԃ?8�=>O�5��颾ש��U�=k>_�2?�5#?G�?ѯ�>,��>|���j�=n��>oc?s/�?��o?F��=v�?�72>���>�=%��>���>�?\VO?��s?��J?Î�>���<W:���8���Gs�I�O�5ǂ;��H<��y=����3t��F�]��<�$�;�[���5�������D��䐼U��;z_�>��s>�
����0>��ľ�O����@>F���!P���ڊ���:�_޷=�>��?��>�X#����=宼>I�>.���6(?��?�?��!;�b�-�ھбK�%�>/	B?��=��l�����g�u���g=��m?��^?��W��&��p?)�}?�ξ�7W��I��Y��C�򽜖�?��>����a>w z?�s?~H?������|�	J����d�z�o</�I>�+�>��6���p�Ｆ>���?&G!?>io=g�>"#���މ��IE��a?(T�?�?�o�?���=�x}��ٿ��Ѿ�R����u?�>�B��SL3?mѽ-¾lGݾ}cg���Ӿ�c��e�¾����䶾�'��yW������ż�h?��h?^�[?��v?�� �`o�qKt�sڃ��#5��E������B�n�J�h�;��a��l�R���~���=c�j���K�^i�?g�?�t��F ?�桾�2�Դ꾶1Q>Շ��l%��H=ͽ��<d?`=FX���$�X ���~?�β>{p�>o�B?	�c���=���6�.�=�'��3O>-�>a��>���>d�����1�:��Ϣ��@~���ǽ?�u>�c?�~K?�p?�!�g3��!���#�� %�zF���+@>]w>� �>��W�i8$���'���=�U�p����T"����	����=f/4?o��>"��>
6�?fI?�m
������w�
91�ej]<�»>��g?��>���>нq !��N�>�l?|�?��>�Zݾ��Q���ۨ��F&	?�x ?Hs�>���=b9;�p\H�����꒿gH�+�B>��[?7���Μ���n>�τ?��R=�3�����>������;���&�@�r���	�G��>/��>l��=* ���+�L�v��ǥ��1)?�y?�?���)���~>?b!?��>7��>��?���>�-¾"6�; �?8^_?�J?<�@?k��>"J=S���~˽�")�n�=="i�>Qg\>��\=��=�w�.lZ��� �u�9=��=d���ֱ���9<�̱��41<|�<B>5>75ܿ�[?�D��x&/�(9�������0�ae���|0���<p�4�e�4����8�;ќb�|@���������s�?;�?��	����CK��t�e�����ި�>��¾����G7��,_��o�Ⱦ�=�̲���R�]U=��e���S�{p?�W��u��L'����$�?$�?�k?�����-�J�����=$j=�g%��p��~�����οl¾��i?�[�>E��V��k�>l�>���>�q_>^ ��]7ܾE=o?��-?'%?Qw����տ�м�l|��	�?6�@}A?9�(�R���V=���>�	?��?>GV1�I������T�>h<�?���?-�M=��W���	��e? N<.�F�m�ݻh�=�A�=Q=o����J>T�>��@TA��?ܽh�4>�څ>;s"�Ǫ���^����<��]>��սE7���؄?�&\��,f�;�-�����&[>wV?}S�>_�= N3?s�H�L�п�]�d(]?��?S�?"�*?JӺ����>�c޾4�M?�6?+ԙ>s&�v�o��=�����:صݾY�Z�\�=e��>Q>�a0�Yo�g�Y�5�ݼ���=O����ɿ&�d8"��2D==#�<�WE�Ӟ��X����0���u��㌽��=s�	>tT>��>��J>�Re>*�c?~�?86d>��y=�a�ꡋ�uD�������g�K�"�/Xr�?�⤩�R��'־)��*'���fe��:>��]�=e[�Fj���'�wj\�&O:�L:(?�G>3�پϢH�5\�;^Ⱦ�p����}������^˾�1���h�ȯ�?&�D?}���MP��O�A2�%7��0kU?��影������=(�D���+=���>�=�=�Ѿ�15�]�U��o0?�o?zK��Q��GE*>#~ �=L=/	+?�?:Ye<�/�>��%?H\(�(�w�[>k|3>'z�>C7�>t>�7����ݽq�?�T?�0�����$�>-{���Zz� �]=�2>�4�H ڼ9u\>��<񜌾f�_�3��)��<U(W?��>��)���b����wA==��x?[�?�/�>k{k?��B?Wͤ<�h����S���ew="�W?i*i?N�>Ո���	о�����5?H�e?��N>�eh���� �.�4U�$?p�n?�_?ۋ��fw}�������Co6?��u?iJW��/�����ܲI��R�>ȱ�>^��> �D��g�>�v?��æ��;���+��Z�?��@���?JH�=F+=� ^�@�?��?�����Ӿա��}����<����!?�˥��=����I�\j��^d?��?�4?�V�������
�="���9�?ԅ?����%v�<���ɿj�;j�%5l<t~�=��J���o������8�XȾ��0�����ࣃ>C�@����@S�>bL�m��7:п�ȅ��	ƾ�~��?��>!��A\����g���p��=��CB�M&��hM�>2�>p���B���1�{��q;�l����>��Z�>��S�)$��u���޾5<��>���>V��>+2��O⽾ř?d^���?ο����@����X?�h�?�n�?p?`a9<��v�Ί{����0G?��s?(Z?;z%��D]�m�7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�b�|=�>���>g>�#/�y�Ŀ�ٶ�>���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���J�!�C0=�TҒ�¼
?W~0?{�f.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�Ź>&܄?��=^r�>[`�=�:�������>_�=���j�?�HO?���>��=��2��J,�a�C� 1T�K$
��B�U'{>�c?�N?�'_>=�ؽ�0d����нս�C1���@P1��z���Mֽr�<>�/;>�>p�>��ɾ#?7�ݾ��ٿ�Ϡ��
'��b?D#�>��>j���)@����>�S?���>����¿I����Q齏�?���?�F?� ۾�d?��X>�b?e�=>_1�~T����8�b��=�C?����^��6(�����>%�?�	@��?D8v���
?�d��
W���~�E�󾣅��#�>J\'?O��3X>�q?;��=�o� Ŭ�w�t�j�>�?��?�E�>[i?~	v�D�.����=>&�>��U?jp�>�[#���%�T>�;?�I�47��~Y
���|?@�	@_�@�SR?��9�\ᨿ�=������'O>��t=�D�=��*�0Y�=U�[�wQr��2ؼ/63>�Ū>��p>��v>2K>U�8>7h>����u#!��s�����I	/��+����̹g���;�����������m;�7����5��kL'�"#����O>��D?4?#?gwH?�{?�޽�� >h�����>\<��S��-�
?��e?�S|?Z�-?�Ӥ=����<)��A�r�����%�����>�U�>��?�.w>ěU>.�>!Up>�>0T�=o+�=//�<E��<�u=���=�2l>8��>��>��7>X�>�~��_1��!k��#v��
�����?�����J��:������Pe����=L-.?��>Ñ�; п C���G?񣔾c>���)�>r�/?glS?�>�T���d���>�	�!Df��(�=<�
��gq���,��O>�;? �">v'�>l�I���K�gt�����0�>�%+?邾Auw���H��=�#��#&X>%�>����"��Y��0����F��^=�Z?��>q4����������j�u��?>��/>&�<��<�SZ>�Z�1����M��� ��8=Ma�>S[?;),>yz�=���>�F���P��x�>��A>!M,>�@?$#%?~L������<���-���v>15�>w��>��>�{J�5�=���>Ib>���������9h?��NW>�~���_�uRt���z=���� o�=\$�=&� ���<�`�&=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ$��>ۡ�@���z㌿I�����'>Gi�>��2?����|���e��tr�>A�?s�ᢱ�~�ȿ$��*��>4��?�S�?tQ�г��{J8���?�?Qf?.>/���s�����>NtD?2�`?�:�>t.,�-�4��\%?��?���?';>��?sv?��?^�]�u[�t���u߉�/��=~~�ol�>��(=�Yþ�5�����ē�{Xj����-2X>��>=��>;����û��_�=����ľۿ> �>B:>��>a	�>���>Ͻ�>	��>���Ҵ�\Ku���T���\?@�?{�E&r��4�<%�>&>���>-^F?�$��*!��2�>��`?p��?��_?-��>����}��]V��N�Ӿ���^4>@�?i?�p����5�0��A4��>�>�.�>e��;���R�f�W~K��z�>0L?䇴>$�T�1?|+?���>%-�>��@��ʬ�Z�K�n�?���>�ƹ>΂�?���>����5~�7}��e����_l�נ&>׌?h<'?\��>���������_� =>�e~>�r�?�x?;�/�G{�>�ǉ?�c?SR?}�>ú�gO��mS�s(�>j�!?�����A�[&�D=��?re?� �>M����RֽG
ټ����I��
?�5\?�4&?K���9a�mþ��<��"�C�[�[� <fG@��>\�>�=��I)�=�J>���=qm��D6��+i<_��=���>�x�=6q7�-��6�0?��������=�x���5��m�>q�ѽ�6�T�?�D��p*��e����䙿�嘼�;�?or�?�A�?%Β=��r��M?��~?�5?�-?Z#�� ����9���B��m���W$�^��>8�>j_��& ��뮿L���?t�b�o���4����>�%�>�a?�8?:k>��>r��0)��x�9�`�l�+|$�A%W�!�I����䗾^\�����˾�����>L'����>2?8�>ZZ�>���>�z[����>%D>���>
c�>�U.>4�=�b�=�Z�;�OR?������'����q����6B?wud?A�>�h��������?4��?4s�?�Xv>\{h�Y3+��c?�3�>����m
?):=Y���ˉ<K��s���b��G����>�e׽�:��M��`f� m
?�4?t��ǔ̾܅׽���I}=.X�?]v+?c�(��U���p�S>W���P�4�(�b��n����$�#!o����G��\��o�&��`.=��)?�G�?�-�w��=¬��cj��>��t>U	�>�>�f�>MjP>���&1��\�u)'�������>�z?;�>�H?>8?��L?��K?�ʊ>4m�>⳱����>Q_~<u��>s]�>�=?��1?1 0?5P?��%?�@>�������~/ھ��?}?e?0��>�D�>�<��ѿ��$��Yc��C#s���N���=e�=�ͽ�N��Nhi=��Y>�X?�����8�2����k>;�7? ��>d��>`��-���<��>1�
?FG�> ��}r��b�?V�>~��?���=��)>8��=ߌ��VӺ�Y�=������=t7��Bz;�f<\��=���=r3t�C���%�:���;�n�<A��>?�>?�	�>��;>]�T�4$�Y�k��}�>�k>��N>�y>�wƾ�9�������H�g�>y��?3��?#oq����=�J`>.����
��g@���B�Q⺽^(�>�6�?-�y?F�?��^?�W?o�=*�&�-��&����*ɾB+?{,?q��>�����ʾ���g�3� �?8[?�2a�q��~3)��¾��Խ��>�S/�#(~�����D��d��n��ۏ�����?=��?�A���6�.}�𺘿f��l�C?2�>{T�>��>H�)���g��(���:>ˋ�>�R?*6�>u�O?��z?�x[?�T>�t8����������%���!>��??���?��?>y?��>��>�)���cx��B� ����^R����[=r�Z>���>��>{^�>��=�ɽ�6����>�:��=�c>���>rz�>�z�>]w>K�<��G?w��>����y�<ݤ������?��u?��?�m+?mj=���F�g���@�>Cr�?���?�Q*?R�S�7��=�wӼ궾�Er��/�>���>�ߘ>Y1�=�	J=�i>F�>x��>K���y��n8��N���?%!F?[�=˖Ŀ?^m�������������Q��m�W�������[��+�=������̨��V���ZO���X������;��k?(1�=���=9Q�=�%<�Ѽ:q�<��b=Ǩ�<�/+=P�D�QS<�N�;��0�v��у;�t�<+�=7/����˾��}?�8I?ٕ+?��C?@�y>?>7�3�g��><g��<?f/V>�TP��}���o;����,!���ؾjn׾��c�pʟ��5>-�I�k�>K3>Sm�=j��<f�=��r=��=�KU��!=��=���=�d�=+��=��>X>�6|?U�~��ڝ�)�8�=�@���9?/��>�H�6��ak?���>�B��H3��5��5A�?�*�?��?�*?V?���R�>�V��!Y�=:N>�������D�)>�Z��|��>mV�>�Eb�~F������ۋ�?4��?vO?󄉿�ο8Z>�C1>�>�UU�3�p�m��a�&(P��� ?��8���;R�>���=gBݾ�4þ{==��4>�e`=�!���\�yI�=�f��xi=?�r=c"�>EA@>ޯ�=�`���/�=��Z=���=�I>ꮚ9m�/�ħ��/D=h�=��W>uc>]��>��?�h0?Yd?%)�>�An�5Ͼ�#��-�>���=��>B6�=�
B>Lq�>�7?��D?��K?���>Q��=� �># �>'�,�V�m��Q��ӧ�e��<�?3ӆ?wƸ>PU<�7A�8���p>��OŽWh?�J1?*s?�ƞ>9����v��h"��]�<�Xy=L�"=m�b�i�*�mY�^Vj��o9��>�s�>��>�?�>3��>�u2>�"><��>I/J>�c�����:�꼀d=	��<�1+>�ͅ=<��9�>��
>��;�ZѼ�1���8��6��z<,�J=`��=,��>dQ=v�>һ�=_���)aY>���9[�HiO>hN����G��Yp���5����F>�v>ŋ�:��2�?��U>��P>�1�?��v?���=����a��e��I�������>�pV<��Ӿ_a�L�k�j�H�"�5��>��>��>(2m>�,��;?��w=�F��M5����>�x�����`0�5-q��?��T���.i�	�ȺB�D?�@���4�=�~?�I?L�?4Q�>���3tؾ��/>	���ئ=T��5q�������?q�&?J_�>>���D�mH̾����޷>"@I��O���d�0�ǰ�Iͷ�폱>�����оv$3��g�������B��Lr�A��>�O?��?�9b��W��"UO����U)��rq?�|g?�>�J?�@?�%��z�,r��*w�=��n?���?6=�?�>���=T$���;�>P,	?��?���?y�s?q?��~�>��;4� >򦘽?Z�=.�>���=�&�=�n?��
?��
? h����	����:���^��+�<�ԡ=ۉ�>i�>j�r>���=g="��='8\>�ޞ>��>�d>>�>mN�>�M��N@�8+?x�Ѽ���>w�<?^߫=>��)]>��ٽ�(p����@!���A�����<���=\ީ=��o��-�>J˿pZ�?f�H��TԾ�g?����ed= ��Z��>0.��}m�>�b>c��>j��>3��>j�">��]>���=|�оV�>le���%�(�J�F�M��Ⱦ�ǀ>{-���;�H�����0�A�����#o�x.f�ʠ��q�A���<�e�?f�)�^��L%����	?C�>E61?NT��^w���W> ��>���>s���3����hB�>ƌ?(��?)�~>{m$>}�?�iK?���\�������H�U����.K��<��x���`�������ͽL�k?���?e�W?�G����%>� �?�j��?��&P>T�F����XE>�Z�>�o��a��ϓ��)�׾2��d�>��k?j�f?��<?��3�عc)�7=?��=?f>�?B��>���>p�j��hL?�<>m��>T�1?��L?/;?f�2?;�=���^(p�ɞ�?ͷ��ђ���I��T��F|��=��6=������X<+u�=U�q�F�ͽe��F���Z�<Yf�<w>Ʈ�=羦>t�]?hV�>���>��7?���M{8�侮��/?ّ9=s����'��ܢ���B�>3�j?��?�hZ?uZd>z�A���B��>�I�>�x&>��[>Z�>�DｖvE�@�=�P>!n>�ɥ=[�M��́���	�W���ބ�<�>��>�*|>�)��/�'>A���	5z���d>dR��Ѻ�a�S���G��1��v��F�>��K?��?���=
V�S���Kf�3)?�[<?�NM?�?u�=��۾��9��J� m���>���<���{¢��&��1�:�E��:*�s>�>���v��h��>���ِ�d����E�P~���9��*4�l���j����<E�
>��=
�ԾM�E��P������-�U?Y->����ǁ4����&�=�J?�:�>�z�b�h��MU�Z̾[?�=�?u��==�f�W/��x)�fi	��Ɗ>H@F?��`?�;�?�����v��pC��f�o���E�� q?�(�>�?<�:>�ם=Yy��J���$c���D��>�>R��>L�GdH�(���L���E �?��>ml?2>�
?%�M?B\?.3]?�*?��>	��>�\˽?Ӭ�o+'?N
�?���=4Z��=(^�(�9�w\D��)�>['?uB��Ř>�?F�?Ҁ$?��N?�?���=�d�U�<�/�>���>��Z��ڰ��sb>iM?jS�>:rY?P�?��*>�<�Z~��mm��J��=U�>X�2?��?|�?��>�{�>�����=���=��n?���?+ '?�JL=qgS?ೝ=^��>X.�>��Q>3+?��a?h�v?�ч?l}?4�h>h`=�ru��������������;(��I->珝<�b�=]�>ց�<!N�������|=YCW;I$=��!=	��b�>��s>x��p 1>��ľR��_�@>�ţ��N���؊�Ģ:�C��=z�>��?���>VT#����=���>5�> ���2(?��?�?�N*;Ǟb�<۾s�K���>�B?��=.�l�A�����u�\gh=��m?�^?)�W�����c?�/_?&Lﾝ�9��ƾ �g��F���K?��	?��I��ʱ>Zz?��l?1��>�e��Im�"��a�b�:Gh����=�*�>��bTf����>a�9?��>��i>zu�=�T޾xw|�6����?�H�?XЭ?�Ǌ?�">Jn��U߿d"��֕���`?��>0K����!?Oe�����'����EH�_Ҿ�b���V��)��֫��Q!��υ�yd�0��=[�?]J_?�Yp?��d?X�����i���n�c�}��d�zH���g�M��5:� �:�l(x��X�&D�1�Sߺ�G9��X9��#�?%@?������>3l߾�1ž�^��,�>����#���iP=�9�ͮi<ګ�=���8K�W�ؾ�"?6۵>�+�>��,?Caf���h�:9�o�W���(��z�>��>��o>�w�>��d�+�����n�c�ѾB�A�j)7�;�>xZ?��N?�x?u�)��7�
[��D�C�89;��m����>�@>�b�>)\���9W��w龿�D��_��
��=o��p�^&+�Wn4?��>�� ?���?�=?�5۽c奾4B��o�W�����Y��>��?Y �>�{�>�	��~:���>]�l?@��>��>󇌾0U!���{�~�ʽP��>���>���>p�p>�,�n`\��h��r���9�f��=h�h?|����y`�P�>��Q?$Ϫ:�lS<�W�>�y���!����/�'�Oi>ؒ?��=�4<>@ž|�4�{�W��o�'?��>��]���4��>��'?g�>�Y�>�c�?��>xy����=Q~ ?�)t?��d?�	V?�?�2�=����r����/�K��<d|�>�3>���<w��=����k3��m�̲�=��=�%�<s���δ�@wl��<f=�֠=�>9>��ҿA	N�������� �k��t�|�����Ǒ��̽N����	ž�,Ѿ0� �~���h�;� ���H���g���?~��?x�����V�������y�8�¾lƗ>�����)~�����a%d��E�v&¾�E���'?���n��qu���f���&?ʞ���Vǿ8���L��%�?�r!?V�x?����W$���8���>���<V�N�-�����qϿ����?;]?o��>[=�`����_�>l�>�"W>~Bn>E���rE��X��<|?IZ,?�� ?�q���ɿ{����P�<%��?�@�yA?��(����	�U=���>��	?��?>�D1��H�����S�>~=�?%��?W�L=��W��	�~e?��<��F���޻9�=�X�=�<=1���J>�T�>����TA�C:ܽ�4>ׅ>w`"�����l^�2��<7�]>0�ս@��5Մ?,{\��f���/��T��U>��T?�*�>U:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=s6�����{���&V�}��=[��>d�>,������O��I��U��=z"��Pǿ�b(�� �a��<7P����$��=-�����<����ك�������=���=�]>�x>�.>�>[>�S\?7�h?C?�>��F>�.�����Կ���x�~�f�����w�>���.�N�ʾ��׾1��+�U
'���ɾ�	=�~��=�RR�2C��l)!���b�1F�u(.?�#>/pʾl�M�fm<T�˾�k���؃�s$��;;42��n�0�?/B?AՅ��kV�����u
�����=�W?]�����i2�����=H��~=ۜ�>��=�����2�JlS�.�$?��#?�Ȳ�Q����>'>����� �=A�/?���>s8C�$^�>�t5?
i���\���0>�>t�>(?�>�>�簾�/��l�#?{�J?��ν=B��5��>ɾ��u��9�=��>�hO��T��l�>-o�=�����ݠ<�.��[��<	W?�͍>��)���HS��P�Uj?=��x?9x?�˟>�fk?�C?u��<�����S�����w=��W?�i?�9>�`���Ͼ^z��M�5?0�e?w�N>"�h����h�.�AR�/?��n?S?����TI}��������E6?��v?XC��5�� w�N}�ƥ5>�[?H?*�F�)i�>�a?�WO�>'��gM���R�k��?ӎ@_�?>|�=��OY�=j%?�=�>_���������5[�KU�=��>�h�l�b�Ԕ!�Y+��;?i�?�N?���?����8)>����ڞ�?��?�������G=��R���1�x�m>X^P>[Y��]0y��ξ�oK��J����@I���9�5�>��@�d��	�?�펾����0¿����^��Y�r��?9�>�;=�;\ž�2t�G��I��vN�cYc�Ʀ�>�<>�Z�+��u�|�r3>�Ŝ˼���>J��0�>��=��~��>���e_.<���>�`�>A�W>j'�q�� ��?V)�"Ͽ-���C+ �s_?x�?R�?V!?V�2��}�����μ��D?�h?��X?�~���r�� ���k?|���j��V=�̴A�X�->R�4?Ȇ�>�+1�gq>03W>���>��=��8��#ſbճ��ؾ؄�?�J�?#-�j��>�%�??�)?l���������������6?c>�!����(��;��a���_?��<?+a.�S�$�\�_?(�a�K�p���-�v�ƽ�ۡ> �0��e\��M�����Xe����@y����?N^�?i�?̵�� #�d6%?�>c����8Ǿ��<���>�(�>*N>ZH_���u>����:�i	>���?�~�?Qj?���������U>�}?�#�>��?'q�=�_�>�^�=�|,�n#>��=�?�I�?�M?RD�>!1�=r�8�+/�[YF�9FR��$���C�C�>B�a?сL?tXb>/
��92��!��oͽ�b1����S@��,���߽�;5>�=>�>��D�Ӿ�K.?N���ؿa
��m����(?�\�>Kk�>ga��>�=%-9=��-?���>'�\L���ڠ��G�P�?G�@F7?:�ؾ�,�|0Q>��t>,v�<s觽�<=�N��>�^?Ub���7��km�h^3>[��?a�@:j�?BX��vj?�P ������������mA��	>�7?���X}�>�?٬�=��p�ٙ���x���>��?Wm�?��>�Fe?��i��>�
8_=�i�>��Z?�?�MQ=�����6>cC?������J��|W?W�@�x@_R?}&����ݿW���	��Y��uQt=*�üP^�=Kr����>�����?��35�=s��>�>�]�>Nv^>��=�Đ=cy����*���!���~:�>q��, ��mr���-�;��j}"�u��莿���˻��<��<��@���н�;d e>��<?�OJ?���?�t?�U<�*R=CJr��;�>W�5��=ɜy>�.?�J?��]>񙠾L�g���������hM����>}>X}!?	��>�z>�O>/Z?xQ>�/�>��>�b>^�1=RhZ>}�8>!�>��?_g�>�&<>��>�ȴ�]���h��zw�iVʽ��?�����J��'������4���"n�=G.?��>C ���?п^뭿B5H?�������+�%>�0?`sW?|S>{���9�X�=�>]��X�i�I�>�� ���m���)�1�Q>	b?�a�>�>�����Y����̌�>��?U���a�L���Z��~�c2�>r�>̙�D*��C���=��|u��\�;�_/?{�?�Һ<$)�����oh��+�!>�Yo>\6�=�K >c+?>�����=wӽ�p�=Yc�=�>u7?�R,>L�=�Y�>Z����N�P��>��B>V�,>�??�#%?�
��!��Fۃ���,�_�w>�h�>1�>�>�5J��[�=۲�>��`>�I����PG��@���V>`}�%�_���v��sx=c��t��=%�=oQ��!�<�B�%=�~?���(䈿��,e���lD?T+?` �=�F<��"�E ���H��F�?r�@m�?��	��V�>�?�@�?��P��=}�>׫>�ξ�L��?��Ž4Ǣ�Ȕ	�2)#�iS�?��?��/�Zʋ�=l��6>�^%?��Ӿg>�>e=%���� ���7k��:=�H�>��2?C����9>�X����C>�O?�Y�.٣�S�տ07��AZ?,}�?w9�?$OV��w����k��??���?2QA?�<6��R�#>p��>�4I?�KI?\�O>�6��؁��>R�?;ݪ?tZ>C�?YE�?�>]Hz�m�T���ڿ(��dT��92�<�"?&��>g9���w��.���@g���z��?���`>fD�FV�>%���?雾�4=t�F�5>���������>쓑=@�z>�X�>��+?�	>�ܛ>0��>^i �v%�������L?6��?�����m��<7�=��]���?l4?^��}о��>!\?ȶ�?��Z?�J�>����G��￿�����<SL>���>u��>����GJ>��Ծ6D�y�>8�>�ϟ��ھ�;��w#P�`~�>Y!?Ea�>��=c�%?R�0?�L�>�~�>M�EL��ѫB��_w>��>�*?��?��?��ʾ��'��鈿���� Y�s >'i?X�?e�>�ޓ�Δ�����^�˻u�<��w?ƺh?��O�J��>�^?�?<�:?���>=�D��Z"�M��>��'?q&��	5���"�8�_% ?M?@�>औ�$��c�J*����?J!J?��?���V^f�yEھn��<Y6���U�9�=�%���>x/'>�U����C=M2">t��<��b���@�$iL=�>5Ş>��>	�Q�����,?�	�=H�Ǿ��F��p���e��j�>˹�>�dǾ#�y?8�=c1h�I��܀����ξ�d?V)�?Qț?�@<=�n���>?ɑ?��?O��>�f���>���"ľ������� ���><h�>�&��z��?�������T������8 ?��>��?5��>�
J>�B�>��\���������VQ����;�c�������ȕ9�"��^�ž�|�1{�>�b���>8�?ءI>^Ƅ>Kl�>!�����>t�W>G��>A\�>���>�eE>l�>�<�<;���iJR?*�����'�ε�����/B?9qd?�3�>�i�����i���{?���?�r�?�3v>_�h��-+��l?!;�>Y��Qq
?dw:=e/��ĉ<(R������+�� !�J��>)C׽:�_M��|f�h
?|/?�ލ�E�̾#׽J�����=��?T�6?��(�y�_��r�̪^�o�V�*=*����p�����6g��y���z��74y��"�x��; 0*?�ԍ?��������Ѿݗp���,�?v(>!��>�U�>}�>�VB>��	���,�PHH�d�-������;�>c�?�W�>Kk>?"@?��Y?RN?ؤ�>�Q�>x�����	?�U<���>���>��5?�q#?\.?�?:6&?��,>�V,��f���1վ �?BB�>�?��?:?8�,��ذ�o�>��xT�+xM���g�1�=�t�<``�\��:�f=~(>�4?���<�8�:���;�j>��7?ִ�>��>-'��􎁾j|�<��>��
?�M�>� �Xdr��B��`�>���?�N�:�=*>q��=����*�e�zq�=�TƼ�n�=#M����:���<nU�=�?�=8#0�/#`�c;c�;���<d��>~�?���>
M�>O���� �s��9~�=��X>{�S>h�>g/پ�t��� ���g�"y>qv�?�q�?+Zf=�9�=�d�=�]���?����09�����<�?�7#?OT?���?d�=?�O#?l�>��K��\a��& ��=�?0?�w�>@���a��zxC�Tq ?��?�)?��(���]J��5�<�;=�>�m6����?��Y�@���V�L���~n�<pX�?BV\?�B>u��5@���i�#��"�S?��>:�>�;?��G�E�m�(j	�$�>�d$?��T?�>�R?�Y?/
Y? wC>�U>�����𓟿�����>�SH?���?#�?�B]?A��>8>�]��^߾����Z"��@��ُ�Lѻ=�JM>]�>s�>�ѯ>+��=ml����ɽ~l�'�=��>��>T�>z��>0(c>|ф���G?D��>@��כ�����W����;��u?��?�+?��=�D�0�E�����9��>-r�?R�?**?z�S����= �ּD���5q���>���>l1�>���=z�F=Vl>H�>}m�>�t�Z��6�8�c.M��?�E?��=�ƿ"�q�2q�T͗��e<�풾<e�B��v)[�h��=hژ�#�� é�ȫ[�̕���\���ᵾ����"�{�t��>��=6��=la�=E��<�ɼ��<��I=��<�=�n�#zl<�9�~�ѻ�Ј��c&�	�Y<�G=�p��a&˾X}?;HI?<�+?�C?�z>A�>�/�DÖ>����.�?M�U>��K��]����:����`����ؾ��׾.�c������>�mJ��^>x5>r��=%��<é�=�dm=H
�=3E�#u=���=��=&�=Gv�=(�>E�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�.>�o>�5N���2��#W�� M�2K@���#?�:�-�־ᓆ>��>�uھu�ݾ̭�<�,>x(o=Y
��&W��?�=�ց�Kƍ=��[=���>U$W>Bq�=Wн5�=eR=���=�(E>��<���֞�Ή4=ƿ�=�\>��>�`�>(�?J^0?�od?�_�>osl�	�ξ;��� ��>fz�=	<�>@ƅ=2B>��>��7?ˮD?��K?���>V��=[��>��>�$,�-[m��	侯 ���q�</��?҆?���>�4#<��A��}�i�=�u���Q(?|1?�?���>��>���	`�$�J�]�&�=���L�y�V���m�@�������V��=��59�>��>���>��\>�3>/�Z>�H�>L><�G>�X1>�덽�#�=S>=�[��xo���ͼ���@U��v�1����쑽�:��V���%���`==9�=�| ?y��=홒>-9�<E*ɾ��>H<��sE8�b݅=drn�����`�)���6a@�8�a�D�<>�u�>T��<
b�� ��>���>�)>X�?N�?5C >��t��`ƾ}��N#��:b�<9j>�S���x�`
�^c�4QU�Aݾ�H�>�פ>��>Y�3>�$��&6����=\�:-��>�x��*a=�'������������Kc[�}�%=��B?6��<�=pa�?�;?<��?t�?%Rn��B���>N���?n��-龱�2�.��~�)?A&?%I�>�����C�sH̾����޷>�@I�>�O���C�0���,ͷ�$��>�����оN$3��g�������B�Mr�]��>�O?��?G:b��W��^UO�����'���q?�|g?�>
K?�@?�%���y�r��iv�=�n?³�?S=�?�>�ǿ=Qz��ѹ�>���>{��?�
�?�o?P�8�
��>�)���>�V�:�>W8>n��=v�><�?��?O)?Y梽p�����:���Y�"�<Y�;=f�y>�$|>5Zd>���=0/�<��}=�Έ>8��>>�]�>��>9B�>[؟���&�!?c�� g�>�g:?���>��4>��׽{�A=ܽ_��������@���	���鼹l�=>�?>ɖ�=�&�>� ڿ�|�?��>T��^�>�D.�w���9�=�C�>9���K"=,7V>N��>r�>Q۝>!~;V��>&��=����.>>���S����|�t�Y�V�O���\>����E<�����z���@���O��h ���� n����K������?�pJ��H��4�+5	�c^�>�	�>��A?��9�8��_�@=���>%�>� ɾ}~��Ҵ���%ʾ�`�?5��?E<c>��>C�W??��1�J3��uZ�6�u��'A��e��`�G፿�����
������_?�x?�wA?:�<�8z>?�%��ҏ��*�>7/�$';�tB<=C,�>H)����`��Ӿ��þ�7��IF>�o?�$�??Y?�SV� �@=�>>K=?��,?e(�?��[?/3$?�_=��Y?�� >��>�U ?��:?�,?�?$�>�"�>_��E�!����������]���[;u
;>�Q:�lQ������ͽd����0�M�a���3>��e�=�$�=&�-=��> ��>K�]?�|�>Ɇ>$�7?���\8�-����s/?۔8=r߂����Э�����Yt>��j?���?j�Y?<�b>��A�:�B��>9ɉ>"�&>4!]>�б>�%�{�C�d�=\�>��>�G�=$�E�ڝ���	�Ǳ��7f�<j�>lD�>��|>8h���;*>k~����z���d>��R�����KS��H�Z2���x��x�>��K?��?�F�=���x����1f�t�(?q<?��M?T�?���=�ܾP9�'J�W���>栰<�������`V��n�9�HN�:��t>�J��}����>7n�]���82{�2
0�i�F�O�Ų �� j=�����㾩?{�vU�=��>�ݣ�z#��������U7E?�>p��}^�������qX>Oh�><(�>���bF$���a�s�ھ��=��>�w�=s�������V�@�\�߾�H�>��@?��c?w4�?���wJ�E��(Ϯ�S=�z?�E�>�b�>P�i>��<T��xN�f�O���0�h��>r��>����K@�py����v�-�=G>	�?��->�?�2??
��>���?��@?%�?%�b>�_��/Ⱦ�0?>5�?�Y�=�o��d���q11��9�J�>HZ?/k$���> $?�[�>��?�F?��?k�=u��l�1��&�>���>��`�G���1?H>�[O?]D�>�T?�#�?�y�={#E�𽯾����xf=)�>s�?%�?']	?�>��>�V���?�=� �>hd?���?�aj?K��=�L?�,+>��>�=��>��>B?%N?tv?a^G?�z�>瓓<���&ۥ�jt��Ȼ2�r<֪�:<e�=·���i��|��h��<�;�&��>���6���|ܽ�Ž�; ~�>�Qt>���z31>�ľ��/xA>����^)���1���%;����=�P�>��?R��>?�#�s@�=���>�3�>���(?��?&?o�V;�b�H�ھ�L��>��A?���=��l��}��c�u�>�h=��m?��^?(hW�;:����b?+�]?�g�=���þ�b�0�龗�O?��
?�G���>1�~?��q?���>��e��9n�
���Cb�2�j��Ѷ=^r�>�X�[�d��?�>��7?�N�>��b>�&�=�u۾r�w�r��^?!�?��?\��?�**>1�n��3�>��#���m^?�|�>|����$"?>䫻oYϾ�0���h��y7ᾀ+���g��mm���&��:)��т���̽㖻=?:r?��p?
�`?�� ���c���\������W��Q������E��B���B�d�n�]��1�6��oD=`ٽt�[�;��?�:?����>w鞾�B��z��s��>@M�<�{G��kl����<�:�=���>�[�=~�1��mž�a-?`��>��>��?cr���j���ھ��O�Ĳ/���>��>�v.>�&?�ί���;�ݼP��~�:��=5Av>�sc?̎K?ƴn?`���=1�������!���/��B����B>��>ʨ�>�"W��l��$&��P>�-�r����%j��P�	�V ~=��2?$�>i��>�D�?H?.j	�D^���fx���1���<�X�>0&i?4L�>���>;н<� �%��>�l?���> �>�����O!��{���ʽ�>�έ>'��>l�o>٦,��$\�uh�����#9�#��=�h?����w�`���>�R?J��:��H<[{�>I�u�ڰ!����'�+>�|?�=)�;>P}ž����{��5���E+?�?�o����(���x>�9#?A�>'��>뎃?�ݕ>K�ƾ��l��]?��Z?��G?�=?��>8�=h��tǽf�&�L%:=�9�>"�b>��p=�=v���f]�,!��\7=(b�=BS��\����[�;�9��=��<�=�50>%ۿv�M�ey޾����������g��6e������ڀ���ܡ���U�A
��C��?TJ�vrk��
�������<�?G��?V������ٗ��rz��X���s�>62z�h	���T��v-�	4[��}Ͼ�F��_�QW�e=e��h��?Qb:�p�Ϳ�����-&?�V5?Tw?�c2��ξr�0��T�A��>�d��m�0����=yԿy���ڀs?Q��>��澵�D�x��>�/�>�=�=�@�>�پ˔��U�b>�U;?f?t��>�i��ിݺ���Z�6��?c@wzA?3�(�=�쾝�V=���>ʎ	?ۦ?>�k1��?�j谾)q�>E6�?���?BN=�W��H	��e?--<;�F�J�ڻXH�=��=�=����J>,Q�>z���bA�Q%ܽ��4>|Ѕ>"�"������^��E�<�_]>��ս��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=�� �=AĿ��3�w6)�̀�;�Y=L�$��Q��EU�<�0<1���C+���E��$-;+a5>ߙx>�
�>z#�=��=��P?V�]?���>2�C<���Z����1��T�����k����1�Ո����̾��ݾ���)6����++��[L���=2S��j���c�q�N�	�V�
�%?1
P>����{U�礳��u��(��4�%=?2E�m�ϾO�7�pgz��ҙ?c�H?$���:�]�������K���2_?�������ؾ��c<W\�=��(<�Pe>��=ۄ��4���I�MH?�4?�/����d��V�=e�Ƕ�=��-?r�>�ν��><!?tf/����� (>v^�=���>���>�)>O������?L�m?�P=9���ܲ>f������&/�ж�=��(��C����>T8�<�r���=�J?���K�{iW?br�>��)�$��]���I��4�==~!x?'�?_�>)�j?�mB?]К<	���ߢS���;t=�6W?��h?K�>� ��6,оه���5?őe?�VN>h&e�E���.����.�?�o?��?�����P}�Œ��x��C6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������1�q=�"�>���ev����R,�f�8?ݠ�?���>��������>xԹ�T��?���?�t���J�v#�fl�d%�{�=q��=c��=uA�=Մ�IJ�ٵ���w㾍�W���<�n>�\@�F�>:[[�ٿ��ǿsu���Wþ�s���?w��>������]�O��"���C��>�0q?��I�>)'G>�dI�����t낿��4�N�w�>d�]��\�>~�p>������}u<��>^��>�_c>( ��fܯ����?44��ο���]���\?�?t��?��?�oc�����I��� �A1?�qg?Z:C?�߁���m�����P?Jc��y;l�A�6���2��v�=�=?�5�>~S��o�>�R\>hH�>N�m>:�/���Ŀ޽��q&�һ?���?m��:��>]��?O ?o�վ�@���䖾����x���?)dG>^ ������g������`�> 9?��-=�>�]�_?+�a�N�p���-���ƽ�ۡ>�0� f\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>aH_���u>����:�i	>���?�~�?Qj?���� ����U>
�}?�P�>��?%O�=j�>Sr�=`ð�.'�ę#>&�=��@��v?�M?,(�>�!�=@�8�!/��>F��<R�����C�;��>.�a?G�L?x�b>v"��DU1�I!�r�ͽ^�1�#w鼚h@�l�-�	�޽+.5>1�=>�e>��D�&Ӿ��?�c�֔ؿ�e���'��!4?��>��?#��x�s����U�^?Ι�>�D��.���-�����^��?�K�?!�?��׾��ȼ�:>��>�>�ս�۟�9���(	8>��B?t���;���o���>���?Ӭ@��?��h�t	?���P��5a~����67����= �7?L0�s�z>}��>�=�nv�Ż��S�s����>B�?�{�?��>ۮl?��o���B���1=BM�>k?�s?,Do�󾰱B>J�?!�������K��f?�
@eu@�^?5���J`��_.پ�ܹ��w�>W5Q>��
oH��ג>9��=��h=jD���d�>?��>��>3!�>�@�>5 V>�G>�Sy�
��������W�P��%!��K�c�J�d֨�P�&����K�b9¾�����8���⇾`�Ѿ���hL�=��J?�S?��p?/*�>qK���>>����<<�����=N��>
G.?�g[?�:1?���=����]�������V䗾l2�>O�j>�>���>�2�>���;?�u>�S!>�l>��=}@�����;a�A=�4F>"��>��>x��>旘=�@.>���sh��:�w�:6�%�����?�Ӫ���0�=������(��Fql���?�]>p+��i�ο�6��r�R?��N��-/��W��*�=
�+?,�{?}R�>����C���/>�[%��.��;DG�>0�����Mg1�w]>>~"??fr>�>P�2�^�7��P�?B��Ct{>�x4?�겾ʸ?�7v�[�H�aݾ�@B>�ݻ>]e������J��L�{�D�e��{=h�8?,�?D����<���r��ߔ��nT>i�V>���<��=�X>�o�!�ʽlI�<�M=���=\:^><)?NL7>��=�>�>�h��t�\�e�>��'>�� >��A?2*?���e����}�&�,���|>7�>vz>n4>�Q<�-��=���>H:B>��a��|^����x�H��S>hώ�3d�d߁�9�L=ӹ����=��q=7(�?�>�N�F=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ;E�>�f��m��M��(�u��~%=?�>1H?�����H�Ě=�&�	?T??��¤�;�ȿ�v�j,�>�?AՔ?^�m���=�?����>�+�?�Y?yth> v۾ɵX��"�>{�@?ШQ?���>�����(���?_&�?��?�H>��?}<t?��>o���yc6��Ӳ�����^.=�++<�b�>d�'>�C��͌A�YD��B熿l�g�۾�'�b>}�%=�#�>��뽁�����=M��N�����~&�>��t>�>W>˜�>a��>���>�ʧ>�z$=�5�����������K?���?����1n��O�<+��=�^��&?2I4?�[���Ͼ�Ԩ>�\?���?[?�b�>���>���翿�~��~��<2�K>�5�>:J�><%���GK>��ԾI5D��n�>eϗ>\���
@ھ=+��m@��B�>�e!?<��>�ͮ=�y!?M!$?.�m>�>�AF�?��QSE��T�>���>H�?��?l�?�M���2�aG��裂���Z�+nK>��w?�=?/�>r���ݝ��ƙ���4���Q��?�ff?rd�	�?	!�?�r=?�0??�Jd>�o�d�ھ�_�����>h�"?q�OA�(	&��m�D�?��?���>����|�ܽ>���`���P���E?��Z?$�$?Mf���`�+>�����<R����i�6C<�����&>��>q��9�=�>��=B�k�&_/�:P<��=r4�>�D�=��3��~��1=,?g�G�xۃ���=��r�?xD���>�IL>����^?[l=��{�����x��	U�� �?���?Yk�?a��=�h��$=?�?O	?e"�>�J���}޾8�྾Pw�~x��w�X�>���>��l���J���ڙ���F��T�Ž���<��?��>*>�>��'?n٧>�	?�xi�mh־�]��*��y/�&�*�y ��t���+�z�����������Ͼn=�����>ï7=z�?�5�>\m>w�D>�?�Oͽ�1�>\�[>$G>⌾>H	�>xs�>��Y>��<�p���NR?����C�'���o���U3B?�sd?03�>�i�������`{?Z��?�o�?4v>�}h�&+�Sj?�:�>=��hl
?�y:=���@{�<�R������L�������>�?׽M:��M��Yf�si
?y-?}��҇̾gd׽o���v�=�*�?J�(?�*�R�� o��X�F�R�IQ��!G\�cv��o%���n��(���-���r��b�'��q*=�}*?�0�?�]�-�W���
i�M�<�=a>e��>���>C�>��F>�	�X12��]�2}'�y]���R�>�z?�j�>��/?�"??l�[?�C?��>��>��Ǿ%<�>h�<gK�>�t�>b�?�*N?3G>?��?e�3?�t9>Z@�O����n�?0-?f�)?o�,?Z��>%�R��[�< Ӯ��==&ˀ�:7I�
=�Vv<���#�=O=rk>L�(?��^��2�����B>C1<?���>?��>��m��p��%t-�cſ>v��>ðO>
r��I�n���nX�>q�~?P�μ���<�w1>�C>�M�<�5<hv�=��o=���=�^ѼkJ��2�=��>J�=�A4�h���T�=(L=NA�<ז�>��?���>vj�>�d���� ���:(�=�X>2�S>g�>5پ9w�������g�r�y>�j�?Bf�?��f=���=D��=����9�����轾�;�<Hw?�3#?�=T?���?I�=?!Q#?�>>�&��F���j��������?��+?��>&���D˾:���?$3���?t2?"�a�]��]�(�c�þ�нʎ>��/�E�~�?)���B��bv:Yw�_.���n�? ��?ׄ9��77��+�4m��n|���C?;��>`��>�>U�(�rBg�<e�o�;>R�>�R?7=�>�:?��t?��X?a3p=�)x��!�������"����>W<?yك?)r?jc�?bb�>���>n��A�F�������<���h���u=�`>o(�>�%�>�S�>$��=�6o����!��#�>B9�>1�?#`�>�O?`�?>{���H?DO�>�R��_��4���R���m<��Gu?���?q:+?�_=��s�E�`p��4	�>�8�?�ǫ?��)?r6S���=�ּ�𶾖�q�큸>�>d��>�<�=b�H=I�>�6�>\Y�>���q��^8��+O�`?�F?|�=,7ƿ��q�Afw�f��ys<�͑�όj��䍽��O�qϤ=���@t����X�Z�����M������S:��#b|����>��=*Q�=�F�=�N�<xļw��<-�<=,�n<=�l����<�>�%��K�9;ɻX:<��E=�1��˾�x}?� I?΁+?��C?��y>��>�1����>�m���/?SV>ڨP�n���/;���������zؾ^g׾4�c�pɟ� �>N�H�~>�3>D=�=A��<���= @u=	f�=�|H�[3=>D�=���=z��=���=P >�i>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�`?>��>��Q��0��>\��FX��S�;;!?!�7���Ͼ�#�>�=�4޾��Ⱦ7�(=�K->L#U=OY�7<Y��_�=�z�?=�w=��>u	E>�;�=<(��&'�=W�L=��=�mO>�H<�:���#�H�3=���=	g>��%>�L�>b�?w�7?^�i?2^�>gl��qؾF{ܾ��>��>�3�>�l�=@;�=�|�>RU2?��B?�JK?���>���<S�>�>�u$�F'l�Q��|� ��<�?u?��x?K��>��9=�b2����ETD�����Q��>"?S��>��>c��|ݿ$�4�H3��ޕ��ϲ;�ł�^T����=�Hػ��-�����|�=g?�>G�>�Ź>G]�>���=,q)>��>4{�=�V<=$j=�����9=+2M=�y=�,��]��<m�ݼ/J=��߼Kg���da��l��T����޺6ͼ��=���>:�>�3�>��=���T2>�ӕ�TZL�H�=~���a�A��*d��}�Y�.�E�7�K�C>��V>������*=?O0Z> A>N��?n�t?*�>(����Ծ^T���e��T�D�=�~	>�;�l�:�eB_�HkM�%`Ӿ꫌>C�>�6P>���=	{�j�D��O>\Y�cmH�,��>��T��"�=��ҽ-�v�����?��eaf���s>Sel?��]�=��v? 5?�?1b�>�9h�X|P�:J�>N�H&��H덾����06��[?=R$?�?����ad��C̾����ܷ>�AI���O�����*�0�����˷�h��>������о�$3��g��S�����B��Nr���>��O?��?�8b��W���TO�b��� ���p?L~g?w�>UI?�=?�(��yt�Rt���q�=�n?&��?�<�?L>s��=ڔ@�aL�>�j?6��?��?F\?Y����=?�o`�a�>%#=����F�2>��q>B�P=��?Zn�>��>����������v���f�v��=��A=*̨>���>ԇ�>oC�>S-p>b7>�?>�8�>��>6"?>Tŕ>̛>)�ؾ!2��P?��<�&�>��?>�e>��_>g��Y�w<<>r9���92��CF�K &���>�(�=W��>'1ĿbԚ?�3>=�(�>�3��~����={_�>J>~���>7EQ>�κ=�Z>F�?أ$>!�f>�Y�=5���/P>>
�X���J�UB�����GA>�'��@�@�)	�"����}��;��}���6:d������?��B =�J�?Y��Q\m��*�{~p�yO?��>�F?�^����#"=��>Z)�>*��XI��r̋�U˾�t�?E@�?�Cc>��>��W?�?G�1�3�tZ�$�u��&A��e�f�`�����_�����
������_?��x?8vA?y]�<-:z>o��?W�%��ԏ�-�>/�h&;�Bq<=y-�>(,��h�`��Ӿ}�þ@?��DF>��o?�$�?Y?�PV�`Ww��d>6�??7?��x?t�;?u'?�W���%?�>�n?��
?��#?�1?��?�9>��>>��Ҽ3H���h�W��o����Aƽ!��%�<6�=}�<����ݞ=�r�=����{�Pfc�b`�d�E=/�[=v�o=��=�"�>G�\?��>��>ŕ8?
_���7� :���f/?ۄ!=����&��f ����K�>��i?!�?1�X?�V`>��A���C��7>��>C�(>�q]>�ï>���C���=�)>۬>�ڤ=�W�C��+��{揾���<�[>5`�>a�y>s.���S->!7��A�u��Qc>�_T��
��ǱT�;�F�L1���y�h��>DL?Z�?�ޤ=���ɛ�=qe���'?�<?�	M?�6�?���=��ܾI{8���H������>l�<v�	�k��Փ��#�:��J�;_�q>�+��%�徲�)>2��񾾕r|�n�H�v�޾����(�ф|�~��P���OݾɅ<h�=�Ѿ�3�oF���X��Y�F?Tn�= �(�������MF�=��>4!�>�t�<�wN�#�V��<��錼�,�>�I>�f�=n���I��)��.��>��D?Ka?�0�?tJ���kt��0D��( �89��~ )��
?��>�#?xJ>y�=-����)c�d�B�M#�>F��>�o��$G�I����,���&�Ł�>�?�->IU?{Q?V�
?^?�~&?3�?{��>~ޮ��ϳ�*R,?���?!l�=A;�7�m���6�ڇC�/N�>��1?��Q��9�>��?�?��)?FB?-D?*�=����w�1��[�>;��>�W�'֮��d>abG?��>�3Y?^�?E�=�b<�ތ���*�<��=��/>Z'?��?�?��>�F?�ݽ��Z�o�)��s?(�?�߆?9�>��>��>�J?�>��? x:?vg?�Sq?,?pF�>�2;g�#=�Yɽ��9�͚E=�>=�=��#��*��n��	��7J9�J�<��9�w��=cl=g�p:�xG��x@�t[�?��>��t>������2>F�ľ�}��{m?>���������=�;�h7�=��}>ȷ?h�>�:!��܍=1��>]��>����'?��?�?���;Sb��پFXM��ٮ>*LB?�Q�=�)l�AW���,v��p=h�m?��^?��X��	��Ɲj?�D]?�VӾ�"����ǃ������K?u�?����+��>��j?{b?2J?cT���[��ݜ�Y�Z�aaG���=�܍>N��Ыb����>:�7?��>�&Z>�
>���6���X�$� ?�x?]w�?U�?$�>��j���׿Wξ�N���]?5&�>�oq��k?��м�g�P>���1� ��,��������z� �������[f�9,��V��=Ǯ?DE?�}?��x?s�!�O{��OZ�b̋�&ZS��ʂ��V�Q�[��D��T5�`p����D����> �?W"�8����?��<?:<!�2��>����Ӿ�H۾ӌ>�ú�1�~�s��-;��L���=�I9�0�p��|���.,?���>Q@�>�FN?�P����f�C�D��2���Ⱦ��k>�z�>h�>��>О=#ȧ���	����숾d��'��>zG?˻5?���?�'�	`N���w�IF&���ɽSϠ��0�@T!>�=�v~�emཀT���w=���u��Y���ӷ �����&?�e�>Q��> Ô?�?7aa��K��Gѩ��B<�zY�<k%0>bK�?���>��>���c���K�>��k?,��>�y�>���}t$�Mz�f]��d��>W�>�| ?�J>V+�wg]�-P��KY��Z�3��B>�oh?u���*e��˙>�S?�Uu<4�":t�>��,������.,���>�K�>6܎=�%;>ӓž��	��+~����k\?�H?7�c��)*�^��>�}+?��.?j?�Ѓ?�.>?��ǃg>��L?2"b?ږI?�� ?��?q�>,��Uy��@�R�.z��7{�<�	>d�[=�=��|���ľ�8,�"� >��>R��=�>ҽ~R��8=�>!֩=y4�=z?�PE]��N����T�s��wʩ��m�6�ž����*g�Y#���s���Y�|f���۔�l7m�=���y��i3�?���?8
��+�9��C��9��#��]�>�摾�J��^��NT��c}ھN�{ξC�n�n��@}�iG�8�'?#���,�ǿE����<ܾx! ?�? ?:�y?����"��8�� >q�<F1��8�뾳�����ο���Z�^?u��>	��A����>��>�X>kOq> ��#瞾�A�<V�?�-?��>+�r�D�ɿ������<��?t�@��=?38�&����ֻS��>��?7��>�ͽ<Y��������>�
�?D��?m|�=��K����خi?�t7=��>���D�c�=��{=��;ko��P>�L�>�w��$��)��JA>��>Kd��_;�?6k� �=�<�>����#,�5Մ?+{\��f���/��T��U>��T?�*�>X:�=��,?V7H�`}Ͽ�\��*a?�0�?���?&�(?7ۿ��ؚ>��ܾ��M?_D6?���>�d&��t�Ʌ�=q6�����{���&V�x��=_��>e�>��,������O��I��R��=�B��vοW�*������=�=B����9c����UA=�Ӎ�/�d�a���ڕ=^>�>Uۀ>�4>��=0La?�n?�,�>�T>7}@��B����޾u�<^n��t�=����x��E�޾���h����	���|8�N>��:8=�8��=ER�����l� �|�b�H�F�ߧ.?@�#>f�ʾ�M�M�<�ʾ媾�&������ Z̾��1��#n�ȟ?��A?/݅���V��"�T�j�����W?F����R1��&��=i����$=��>;-�=�'�13�~iS�q�0?	�?@���C���u,>����h�I=�5*?���>�4 ���>��$?�,���׽ղ[>�<>��>�u�>W��=A������(�?��N?;��'����͐>��Ⱦ�덾)Z�=�>��&��!�X�?>���< /��H$<2q��n�F;<$W?幍>��)����C��#���d>=��x?��?��>�rk?d�B?Ǘ�<k;���S���$�w=��W?S'i?Q�>󬁽 оL���F�5?��e?�N>T}h����.��>��#?�n?�R?����d}�s
�����V]6?��v?s^�vs�����n�V�U=�>�[�>���>��9��k�>�>?�#��G������~Y4�Þ?��@���?��;< ���=�;?x\�>�O��>ƾ{������2�q=�"�>����~ev����	R,�]�8?ڠ�?���>&���ĩ��p >��پ�1�?(�?V$׾��~�է��d�#8�?J�>����'P��͎�.�����K��9��:��j������Gal>��@e�l=�?�#����Ϳ*-̿:l�����Pփ��Y6?=@�>������l������G��DG���v�if�>��>�0��ӭ����{��l;�����=�>�M���>ݛS����������9<�ɒ>L��>Յ�>����.ٽ����?�V���3ο�����z���X?5c�?io�?�?��2<�.w���{�O��)G?��s?�Z?1'%��]���7��R?��E�Ev��s�N��\h��M>�o?���>�Q	��R>�&>��&>��C>�@6���Ŀ�c���|ʾ�o�?���? ھ���>�Ĝ?�]7?3�/e������s��>�*?t�>!�Ӿ�p'���F��fa���?-??�ag��-8�9�_?p�a���p� �-�y�ƽ�ۡ>��0��c\��4�����Xe����@y����?9^�?<�?5��� #�6%?��>����g8Ǿ���<*��>�(�>]*N> A_�ղu>%���:�j	>���?�~�?�i?�������:W>1�}?̷>&�?��=^��>���=p��L.;���!>���=v�=��?�LM?���>���=8��R.�<LF��R�4#�ĖC��%�>j�a?�:L?��c>�(����.��� ��ͽ�.�_E��?�H�%����C6>|H=>��>� E�g�Ҿ`?%�p�ͺ���ߞ��/?[�+>B�>�{��[!�A��?��>�a��9���J��{�E�F�?p:@D�>]2��ۏR���%>$|Y>ި�=c���$��;��|�>�j;?��n�~�sqb��*n>gJ�?�B@���?�ep��	?���P��Ca~� ��K7����=��7?�0��z>���>��=�nv�ֻ��K�s����>�B�?�{�?N��>�l?ǁo��B�b�1=�L�>��k?�s?�<o����B>~�?1�������K��f?�
@pu@P�^?���ND��ٷݾ0ľ<��=|�i=s��=r�� ��=:�=�+@�n5,���=�W�>���>�V>��^>��y>]j>�}�����4�������&�O'�FI���ھq6+���) �xJؾaʾF��7w����R��s��9��D��N4>��M?��<?�~?��?IP=�-�A>=S���p>�������	>M?�1?�k6?M�4>
�k���j��Rs�q���_����>أ�=U��>��?G��>�x>̵�>p�:>�v>ؾ�=�a�<j�%>�C;>�Ȇ=�>�>��?Pr�>8C<>��>?ϴ��1��p�h�w�p̽"�?����`�J��1���9�������h�=<b.?�{>���?пc����2H?#���`)��+���>t�0?�cW?�>��S�T�:>�����j�`>�+ �<l���)��%Q>ql?�K>��i>,�.���)���T�n1���e>.5%?����à_�0�u�RG�1|����6> �>G>�;%�o�Q~���_�5�@=<&>?	�>�k��C������f���Q>l>n>г<&��=��K>����m����-,��P/=q2�=��O>�t?bF>,�=�l�>#P���p���>�.>^+>\:?�?����q����^���M�Pߌ>�_�>��(>=��=��S����=�d�>.?a>��}<������ng?��SH>z�ĺ�	n���L�b��=p���#>�j=��򼣛C�m�<�~?���(䈿��e���lD?S+?_ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ��>�Ž�ɡ������1x�Hu�=<!>�7?e�s��;a�w*�>ى?+�%ͪ��yٿ)"���?]��?��?l7�����2�_�>)��?�oo?�wx>�;���;���K=u�?�lh?�� ?D��������7?��?�>�?n_D>N�?��?���>&�X�c#Z�K���S��tN���Z7>r#�>���>W3�|�5�f?��r�k���e�!x����=T2}=�S�>�nU��㾏D>�*��5���jZ����>;>Z�;>fi�>�O�>Yƺ>+��>*�>���l���0��L?���?[���sm�-׻<�Қ=��^�+�?�34?�dx�nоM�>�\?��?��Z?�ϔ>�� ?��u���놴��(�<�aK>.�>|��>���%!L>�*վ��E����>�{�>� ��dھQ䂾(�M�<{�>Un!?c��>�E�=�.?(�"?GL�>�;�>��X����ҁN��I�>��>X?&̈́?���>��ž�~ ��������^��>�o?�!?:ۯ>�F��ZӚ���̽"���+YU��\�?�x?3k�GO?��?�t>?z9?��>4y��X�N�)n�>c� ?L�E�;�3�����,�?V�?g�>���iQǽQ�(����A��}?�0X?9�#?����^��l¾�`�<2x����::��?<�,��>�>Q}��8�w=ٽ#>��=\�l��+C�\�U���=݌�>/�=̦G�Z����+?��$�Ǒ��3��=�ss���D���|>$�L>z"���^?/B:���|�>����t��ݝY�{��?�-�?㓖?�����h��<?�Ĉ?Ë?��>4���̝ݾA޾�Ov�d�}�bk���>�ݾ>�Ɖ�D��M0��A	��Q�����˽��N��S�>p�>�Z�>BY�>�a>od�>�Z���4�/K'���3��(���;�1����꧍���\�Ѽ>ݶ��RQ�*�v>p �:�(�>�$?�Ͷ>58>���>��<<J>L�>�>f�>�ʼ>
��>��=�Y*=�].��1R?Zҿ�=�'����g����"B?��d?s�>�@b�Uq���^�K�?���?Mf�?&Tv>/Nh���*�\o?�=�>'��
?�{5=�*��l�<���������A���>�YԽٺ9�b�L�&/g��	?*X? <��̾6ڽKBľ4Ϗ�2�r?O&?�}?�(oT��wm���[�MN�{��s�}������&B��k�w-��D�m��^��u�8�Fi��kL&?+.y?�q��p���v�K-N�� f�g�>��>�>Kw�>&�_>%�ž�JF��xd��&�T���~�?���?�l�>K?��7?��J?-7O?�>:��>����\,?���=l�>���>�H8?�(?�p2?�t?�+?��P>
���w��+�оЫ?��?��?	�?B?vo��E����Z�I�\�e��#���(�=ʬA=
��k{T�M��=�vU>f�?W����7�t���d n>;�7?�z�>�j�>ȏ�X�����< ��>$:
?�m�>�e��#�q�Ƌ�Ӿ�>�H�?&��uO=�J)>�E�=�l���8:�J�=�Ҽ`��=?�'��,���b<���=ڑ=����,|�;7&�;�b<>C�<�t�>F�?ד�>�C�>f@��� �B���f�=�Y>S>9>�Eپ�}���$��<�g��]y>�w�?�z�?ܺf=��=Q��=�|���U�����5��� ��<	�?=J#?)XT?X��?��=?yj#?�>+�iM���^��x��ͮ?k",?᎑>Y����ʾ�憎R�3���?�V?`7a�ļ��9)���¾r*սD�>#X/�Q&~�����D��;������x��x��?���?�@���6��p辁���Ac��[�C?��>�[�>��>i�)�'�g�!�BE;>}�>�R?tj�>Q�M?�|?4:[?��E>��<��������ekG���5>�C=?�с?Q�?�m?�]�>�>|1?��H��I��&���=��a����=�(l>O��>Z�>H��>�C�=Z�ν�e�dX���=2�^>K��>$��>R	�>Gh>���<��F?Y�>�L��?��H⚾��y�K���4�y?���?>]'?(�2=��b'<�.6��>J�?W�?�=)?�QF����=Y���Ļ��у����>e÷>p&�>�_=��<u> �>V�>Zj����cD;�`�eB?a&E?2��=0�ÿ�l�Ǉy��鋾���󕾨\]���ý�eo�C��<�k����2���þ (W�Ȩ��b&����ľ�5��㨋����>QB=�$&>�W�=���<�������R|>=�} ==�=Q����\2=��H�O���������<� ԻX�s=
뮻�˾.�}?�2I?��+?��C?��y>�Q>B;3����>���-?f<V>ݔP������t;�쨨�0����ؾdf׾S�c������I>�KI���>VB3>�@�=��<��=n�s=���=0XH�s=��=�7�=���=�=�>�~>�6w?S�������4Q�"Z罫�:?�8�>~{�=|�ƾp@?��>>�2������tb��-?���?�T�?:�?Pti��d�>I���㎽�q�=�����=2>���=t�2�=��>��J>���K��ဳ��4�?��@��??�ዿ͢Ͽa/>hh->R�>��N��D-�!N���P���I��a!?X8���ھ�l>�2�=)(ܾ{�Ǿk7=�&.>�PT=�f��V�q>�=LW��N7=�-=�u�>e�J>!�=��Ľ'y�=��=�~�=Ae_>�w�;6�;��}��=��=:�j>�4>%��>�w?�m0?(Td?zS�>�k�x-;a���v@�>d6�=�+�>�]�=�B>��>m8?�`D?7iK?�!�>^�=�4�>a�>�+���m�߯�&g����<Q��?
��?H�>la<��>���l=�3_Ľ?�0?��?]��>L����翓�0�,�0��	�5��<�F<�3���ƽ��0=-�A�cY����=*ؤ>���>`��>�Rx>��8>>C٬>��>C+=��=u|�<�]a=�!^�c� <���p��=m�'=��8��	<�X>��a%���#y/��+��oV�J_R=��>y>}��>3�1���;,|�=K��8�'�S���Τ��Ǭ?�-@b�5���.�?�������H>((�>Gw2�~͏��3�>?�>��>+�?��?�З>�7Ѽ�ھ�ذ���վ��=�J�=8�>�af=�^��bZ�e�[�Y�ݾ�>;ʗ>��c>� >�<�aI�N<�๾�k���>��]�k�%��i%��*y�k��B����4N�:��=TXC?t䆿rb?=�Ȍ?�.N?0�?�D�>������x�>�̾�l4�tھK㚾f��2<?�!?%��>���J>F��H̾2���޷>�@I���O�d�#�0����ͷ����>����F�о)$3��g������ߍB��Lr����>[�O?|�?d;b��W��(UO����c)��Xq?�|g?��>K?�@?�&���y�,r���t�=�n?���?A=�?>�;�=D�=L��>��>�B�?��?��j?\\�=1�?A2꽯I�/��=N�7>��>��G>�^Q=�Y�>UC?{��>��Ӽ���O̾F���*���="\�=�P�>��:>���>BB>�-�=�o<>�!�>�b�=�J>I�>���>DS�>k+����+?i0�=g��>��3?;�>ċT>"<���켽���0�;<�'̽V+��V��h=#�:=`Ce>�H>-��>�,׿�#�?t�4>�Y���>@���J@=�S�=��>_ؽ�h~>3}>��>�9N>��>��=e�>TX�=S��S�=�����)�,�H��K���2>wB�����0Vݾ]nt� 斾Ht�����h�]瑿��6�b(�=^�?�8v���w�U^�y�r�_�?��K>ŝF?z���ۥ�<��=>�w�>�E�>�_����'ڢ��y��u�?�8@�Ac>P�>�W?��?��1�3��qZ��u��&A�e�`�`�����ϝ��͓
�I���,�_?S�x?�pA?�
�<z6z>w��?��%�)ˏ��"�>w/�";�'�;=��>K ��6�`�ݪӾ��þJ��<F>͒o?�$�?zQ?QV�O���}�&>�)?�X?&�u?:>?�s>?��ǽq�?;�>�V?�?�y(?�r8?a�?��8>.0>5<������uH���h��B����<���==�s�<� �=HY�='���E˽d���
�<ȃ��[=��b=AX�=��>%�> �`?��>���>h�;?���x�+������;?Q��<|����Ǆ��&��2�Uh,>:qg?�F�?UP?�G>�0=�:D1���,>+l>��>1f>I,�>  ���^)��Ͽ=O|>D8>J��=�μ��x�#�I�����=�3>>�>���>�?���n5>XQ��k��E�Z>��S��ḾYV[��YG��'0��1�����>?�I?�g?QMp=%��|&���1d��R'?�|:?�LK?�?IJ�=+�վ�V:�LM��� ����>��<�
�U٢��,��b�6��Y�<|�g>\���hh���[Z>���,�;�pi-�R�b����VE^�����Ӿ-(���ݾT9�ym��p3�=�ž�7�Q>��yc��yj1?$q;>�w��,C�Oqľ�f6=�]�>h��>�f�<%V����h�Z���2R=U9�>f �>�6v�I���Ʌ?���ؾQM>��3?��\?�8�?�/��楌��Cy��\2���ž�ý�*?w�>�i�>�Պ>(NI=ἰ������e��cT���>*x�>*7(�_�,��r�R\�s��L_�>!��>3Im=�a?�tS?�&?��.?hAK?o?��>� ��%��S�#?G��?<�=JB���V�v�8�8�E���>iP&?��<��͙>�l?��?�O&?��O?V�?R�>6R��@��4�>���>��Q�8î��l>�N?š�>�9[?|��?��I>bx7�����(�W�=�t%>l34?�A#?r�?譹>`X�>z&6;�n=n�<~b?�l?D%J?9Rj>.KD?���>&]�> �5��w�>��:?��9?!�[?p:?�K`?���>�f��B�鼋!ܽ�TA�Cu4��3��}V=�{�=h|S=J�&=V�>��>O=2V�=Ɩ>)b'���=3)3���<��\�>6�s>s�x11>�ľ\��ޤ@>K`���P���ˊ�!p:���=Lv�>t�?L��>�F#�6��=���>/%�>���\.(?��??
?ħ4;w�b�#�ھ�hK��+�>@B?r'�=��l�����@�u���g=C�m?��^?�~W�
��Z�b?��]?�g�g=���þ�b�l�龃�O?C�
?��G���>�~?��q?���>N�e��9n�"���Cb��j�hж=ir�>EX�I�d��>�>4�7?O�>��b>�%�=�u۾�w��q��.?L�?'�?���?F**>��n�4�%>��t�����h? ��>��̾1�?�K����о�喾g�J���ƾO�� 瑾j�����վY�M�����Վ�^E�=��?�b?��Z?�[�?U���]�'0I�����y���	��i ��'d��'��6��/w��j���Ⱦ�g@�[�7e/�\�?�H?��B�4��>�Q��|H��y�^��[�>
�����=qH��X�=��=`�*>�'%�㬾���?1՚>!m>�D?��;���h��U8�8�^���#�)��=���>��>�>@8=�`��eP��(ݾ�7����~�xt�>	_? r=?^�w?�����8��􄿕�����۵�^a�=^;�=�<�=m���ڽS�G<�<Qw����k�p�/�g�9=��?��>�>kǔ?<X?1��\��"9¾57�y��k��>b�h?�a�>�6t>�� ��>�j��>��l?���>��>󋌾�[!���{���ʽ��>Lۭ>���>�o>R�,��%\��g������9�qX�=5�h?}��S�`��܅>�
R?��:lH<�t�>�6v��!�����'���>Ss?�f�=��;>��žc"���{��.��!|(?���>-� �4��F%�>�)?�s�>�ݿ>1��?+M�>��B)+:ם?G�Z?n�]?�W?�t�>��>�Px<K���RG����}�R�>���=��N=�x9=<��g�[�
�%���c=7n����m�M��9@�;�8}<���=H!>�~�N�]����������E�=��6+��M���֡�8�����:�3ﹾ.���Aaڽ�i�ʁ)��ͳ������V�?@��?K����鮽�"��B����	��%<>%����s,��n����(�ҾA��%�ܾ_n>�зg�>�����s���'?�����ǿٱ��^Aܾ� ?�= ?x�y?��q�"�*�8�6� >ˡ�<&����뾡����ο������^?���>��_����>$��>B�X>iXq>����ힾ��<�?��-?$��>:~r��ɿ���`�<}��?��@}A?��(�<��c�V=���>?�	?��?>_i1�G����>M�>
8�?E��?�mM=��W���	��se?�m<b�F�f%ܻ|�=�)�=�b=d��T�J>�E�>*p��?A��;ܽ��4>[ԅ>��"������^��^�<o�]>w�սG��5Մ?+{\��f���/��T��U>��T? +�>V:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?8ۿ��ؚ>��ܾ��M?_D6?���>�d&��t�߅�=o6�Ӊ��{���&V���=[��>b�>��,�ߋ���O��I��S��=8���oԿ�R1��R!��{�tm=D.��l���+�k8H�������(���.���q�??�=/l>���>Ҷ]>Ѹ2>�e?H�p?�څ>��>唖�|��yӱ��[ �͕��-v��xږ�GA_�P�ѾZ�����#�%�GO)���6���پU6>���=aZS�� ���X �Hqb�A�F�5�+?�%>��о��L�O�{<�Ͼ֓���l��ƛ��<T̾6�3���n�r��?e�B?UR��5�T����c�!�G����OT?�����[ ����=�YἙ]�<��>x"�=0��.5��[T��a0?H?U��<���uf+>V����^=n�+?Y�?9�s<�Ѫ>"%?�Z)�����]\>��4>�ۣ>���>�}	>�㮾m۽�S?/GT?r��✾�=�>�,��Z�z��M_=�_>f6�]&�H�Z>�I�<�����Z��㎽���<P(W?⛍>��)���a���f\==��x?_�?�-�>p{k?��B?qԤ<�h����S���7dw=��W?#*i?й>����оN�����5?ܣe?��N>ch�S��O�.�}U��$?	�n?�^?Ry���v}����X���n6?��v?�k^��u��1���W��3�>�Z�>��>~�9��d�>+�>?#�~E�����Va4�͸�?�@��?I�=<�O����=+>?Hd�>�O�YTƾ�8��hz���Yq=D)�>�n��1av����A,�V~8?՝�?5��>g������o��=�/žP�?�A�?(� �)1�/���������m�<uV>5mD����;�ȾNT�{�TA�Ao��+���/l>V�@�u���k'?����߿.��	���c��n�ɾ��	?U�U>r t��p̽p�+�nGh�3E��A�X���&�>Z0>b���6���k"{�s;�_ר�iP�>��,��>LW�����b��O`<�C�>���>x��>����L�����?}��%�Ϳ��������X?��?�K�?��?މ.<��y�*}��q!��	G??is?P�Y?��$�;�]��7���S?"�����C��
}��I
>��(?j~"?m^��=I��>�i�>�@=�R&�?ȿ�η��6���?ѝ�?����x?�U�?�5?p��%����>��V	�M�{�'�G?���>����i�&�,�W̫�P�>��B?�`�R�5���_?L�a�}�p���-���ƽ�ܡ>v�0��f\�uH�����3Ze� ��<Ay���?m]�?5�?���� #��4%?�>Z����7Ǿ��<3��>)�>2&N>�N_���u>��s�:�.p	>���?�~�?Ph?ܔ�����tZ>��}?'�>�?�p�=5n�>^c�=J����\.��S#>��=h�>�[�?+�M?�>�>�@�=>�8�8/�w[F�BFR�(�Q�C�"�>c�a?�L?cb>��_\2�	!�lͽ�f1��&꼊d@�$�,���߽�5>��=>x>��D�pӾ�?�] �к�y�����׾��*?��(>g&#?�B.�t=���,� �D?���>�{��}��3����D�?�@;�>$���[i=�#2>���=�ɀ>p�;~<J°�e��=�t?QV�Ň��nB�g�<>�2�?��@��? ����	?��Cv��H�~��	�m6�RP�=�38?�򾜹y>�d�>���=,8v�զ����s�U��>�j�?�b�?�<�>�Nl?�&o��vB�o�7=���>��j?b�?+�1��F�X�C>`	?�����������e?��
@�{@�0^?O��(i��a��KQ�~���ЖO;3��=X�(�z9�Yg:�-�=�Ξ��}>�d>�.>��>���>}F�>��c>�~��Z!��j��vr����Y�J���}����8q�e���ɾ���;�پ<A1�/����F����;�D��]��M�=�:O?��O?��r?z�>O"�S�=�-�TP���D��+>��>H8?x!J?.!?�
�=���֭b�L怿͊���~����>Ȣ>���>T� ?�s�>��=���>G�{>/|>�:�==\����{�!�T=�v�>ρ�>�p�>�z�>A�@>��>򳿌���1�f���x�Ԓʽ֢?ܦ��z�K��@���?���R����=��.?-� >+���п���zG?����F���.��4�=��1?yjZ?%�>������I���> ����h��@>^����l�i(�	�Q>E[?:�|>b�>;�.��(,�>�I�����<�>�[6?:)����Y������S�u5��U0>�l�>��#�'2���~��Te�K� =C�:?���>��׽\9��"�������:>�Rw>|��<A�g=�ma>Mp���ȽC/L�w�r=�W>`bS>g�?;�,>&�=�7�>%h��#�L���>^A>+{->d�??;�#?���Y���ނ��)��8y>v��>�$|>�-�=�>G���=���>˶]>0wڼ��k�����<�ي[>�f~���b�p���V='��k��=�Е=�, �B>�#�"= �~?���䈿��Sd���lD?g+? �=��F<��"�H ���H��4�?j�@	m�?��	�ԢV�)�?�@�?�
����=�|�>�֫>vξ�L�Ʊ?��Ž�Ƣ���	�q(#�jS�?��?��/�Zʋ�l�a6>_%?��ӾL��>��𢧿gB���~�n�;rMo><V?s�y����v����>9�?���.����׿re��v��>�"�?J��?�@W�z�`�nΫ>��?��h?��>�� ��@B�Y'`>V�X?�xF?��>�q'�;*��ʃ?h��?���?��<>r[�?�s?v�?y��/Q>�{�������I��;v���`�>��=�;�R3�Ra��m���#q�Zz�2�>B�)=��>m_�6���(>�=����Ⱦ�ׂ�Eý>6@>1�?>��>dg�>�>A��>0�=��-�»�������K?i��?����2n��[�<���=�^��&?�I4?wW[���Ͼ�ը>ʺ\?V?�[?�d�>4��>��迿~�����<��K>�3�>GH�>$���EK>��Ծ�4D��o�>�ϗ>����r?ھ�,��܅���A�>�e!?���>�Ү=� ?��#?y�j>&*�>j`E��9����E����>���>�H?T�~?7�?�չ��Z3�k���桿z�[��9N>��x?�U?�ʕ>&��������@E�}@I�����p��?utg?�X��?�1�?ڈ??g�A?�+f>����ؾ����>�>M#"?�I���@�1%�����~?S�?��>E:��Qս�� ��2�������?�A\?w�%?~����`�*�¾��<F+�(�V��l�;��b�\6>��>����A+�=��>;!�=�nl��3�2�n<��=��>���=R5��"���?I��=+Wľ����)>���f���>[��>���wQL?W��=�i�
������"�ؾ}D?��?�k�?�
�J!l��H?AM�?K�?U.?^�ؾDǾ����^(������J� �r�e>���>�2��Vо/8���)���4���<Ͻ��q��=?W��>��>���>��y>i!?�U>��Y��#��H��Y���%�9�S���X+�-���䀾�e�`Ꝿ��ƾH��>���2�>�z>?*�>ł=�{�>�E�=4��>���>���>�?:s>��>
@>��>��NR?������'����ԛ��X5B?�rd?�3�>֤h�񃅿����y?g��?Gr�?�Mv>�uh�G.+��l?�7�>7���p
?WF:=p���<�P�����d䆽f�����>(#׽2:�	M�$gf�(q
?6??x��Ƅ̾%<׽���P�=Æm?�4?� ��=]�u�s� :g���M���佺ox�]া:v0���n��\���ew��l��y�9�c��>�'?><�?��Ǿ����,���N�3�?��å>�=�>"��>���>���=cF���)���U��#�n�Z��C�>�F}?�`�>�7F?W�A?VL?p�??�7�>���>~��Lt�>X*G=�ә>d�>�C)?�F)?}�-?��?�B+?�J=>!c��8��mݾ�?��?=�?�Y?ȭ?��H�M��<2ƛ<�Q�("v���N���=�k=��V�=��`w`=!|O>gZ?_����8�����/k>��7?e��>���>�󏾆���E�<5��>�
?T�>g����gr�]��[�>s��?`�ʖ=��)>���=DZ����Ѻ]$�=����=3����;�_ <Ǝ�=��=�gs�m_��k�:�3�;:Я<�t�>+�?!��>�C�>(A��F� �<���g�=DY>BS>�>Fپ�}���$����g��\y>�w�?�z�?Q�f=��=5��=�|��AU��s��������<ܣ?/J#?XT?E��?L�=?)j#?s�>	+�^M���^������?,,?���>���_Qʾ&ר��m3���?lc?i2a��_�[�)�=#þO�׽�&>�(/��~������<D���y������ڌ�?"��?	�B��u6�+�����o��y�C?���>� �><;�>̓)�u�g���2x;>���>��Q?�H�>�B? Vf?<=l?_��=5�[�C���̖�@pڽu��= DI?8�|?Ӂ?�Of?��>(>�OZ������v�;��ڽ~t��Ei=�K}>)��>-�>��>c3�=V�x3��X�H��<��=�(�>��>Y�>�N�>���=��G?���>�J��g���٤�N���m�<���u?O��?��+?�m=[���E�u���Z�>&m�?o��?�1*?,�S�V��=��ּ�޶���q�d�>�ع>l*�>���=L.F=�;>��>��>�)�Y��l8�A4M�5�?YF?.��=��ſ�q�	�p�J�����`<�,���ae��	���.[���=����a~�*���Q�[������n��絾�Ɯ��2|�}��>?T�=���=I9�=5O�<XǼ	�<4L=��<J�=�zq��Aj<l 9�ݐ׻����!�yp]<�5J=�F��ʾ;R|?��J?+?�^B?х>�>���@��>v�n�Y?�Y>��s�>����7�2���጑�fLپ}ؾ�mb�����ʈ>�T��e>[L8>E�=;�S<&J�=:�x=Z�=n��;j�=���=�=�-�==��=�J>�t
>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�m8>W>�[R��0�j+\��d���[�� ?~5;���˾Z�>��=��߾�~ƾZi.=\46>��[=�,�n�\�8�=�-z�"�9=6n=W��>WE>�ݷ=dĭ�؃�=<�F=���=0kN>�Jʻ]D��e3�10=z��=fc>��&>+B�>��?�1?g-i?�t�>uY�J~޾�+����}>�8�=�o�>���=��>=�>�0?��<?�@?N><�<6��>��>�u�rRe�6q����b����<h��?bR�?cF�>�a��Csh��6��%F�$����,?z3-?q� ?�]�>q�����ۙ1��zA�Y[��,�V���3e���>ؽ!���A��'Ž->�=}[�>[��>CL�>31�>�7\>R)I>l?�>t�=0�=�[>y�<�:�=bT<�9�=����@�>��A��� =��H�� g��{�;��$�+��<�9¼��E��^�=���>�>3��>��Q=u'ɾ�04>�L��]�O��ϗ=����9�:��~`��/��o6�Y�]���I>!�O>C[��̑�">?��{>%�6>SJ�?�u?�>�*"�������x����7.����=��p=���l(2��,n�lL�|�ľGk�>̖�>�n>��=�L��LR��g>�ٚ��o;�rĉ>;/2���=�꽛���C���a��R�Z�閼��E?�p���G >2�?��*?�ê?~�?6$E=���_�>��ξõ>�w1���ǽ-Fc�K�/?�=?�9?>tIξh���H̾q��m޷>�>I���O���v�0�q��Vͷ�)��>������о�$3��g��������B�Nr� �>C�O?l�?�9b�SW��UO�M��!'��q?}g?[�>K?5@?�)��/y�sr��Au�=�n?���?!=�?�>�v�>�#]�l$�>ak?8�?�0�?��x?��޽��?��>�=>��+�;��=���>{�?>�>���>V1�>���>��Ž2y��񤯾ώ���Lｷ�D=|
�;r��>�a�>��>˟�>��6>��>o�>	��>��?�̏=&[�>�>w���9�׾�4?/Rp�m�h>�w5?���>��B>5��<w75�p�ؽ�q�=�+��@P��N�1�H�*���Y�>���=:p�>�.ݿV%�?ZÍ>��
��$�> �7���Ƚ�V�>�]?96�;Jמ>�>8#?��c>���>�B'>�&�>��"=�/ ���>�k
��  �g�F��b�B��g�)>�綾���:�Zq��m$H� ������Iq�j7}��U�ۼ�%�?:������_���P�ք??&�>��}?i�����'>`2*>z��>��>��ھI|���$���Ҿɛ�?X�@��i>�A�>5�U?��?'+&���;�"]�Oht�`�?�Yrb��_�lߌ��e��s���ώƾ\?Pt?��=?��;�'|>N�?�$����O�>/�,��m:�7�x=ڃ�>0���+v��׾��Ⱦ<�#��AQ>K^k?@{�?��?��L���k>1$8>�t�>���>Q�p?g�8?��?�~���3R?�>�>�A>t`?��U?"''?s|1?��?�; =M�R>��`=׹����$򋼫�B�M$�:�`�<�Խ�������?h��|��.����������]�'��+�=\�=�N�=@K">ٛ�>3}]?Ү�>��>ϛ7?��M58�0���A/?��==�|������������'�>��j?�?�	Z?�c>}�A�#tC�r>���>&b&>��\>�6�>ɱ��D�/�=$>]�>3��=�TK��Ɂ�Y|	�����9��<��>u�>)|>������,>%袾��}���`>N�T��(��lS�&�F�1���x��7�>>CK?xY?���=���m����e���(?��;?�L?��?���=�ܾ��8��2J�Ҋ��p�>���<+=	�8�)��G�:���:�cu>�E�.\�>��y��� ?�kQI�{������=�վ��������㩾ɟ��>��:=�O��u�+�Kh�������s3?�g=�图%�j�l�Ѿ�7	>��>�H�>^n����ŧN�Qw��?�h<��>W�A>��3��۾A�;�}s�ף>��A?��T?���?�Q���w�{�Q��}�m���0�#�q�(?���>V��>�U(>��f<_��'
���\�X�>�Z2�>�{�>OE1�dG���-�4c�o=�>#>?�u>?�>��X?> ?sVG?l�?N�?r'4>n��9f��d�,?+4�?S�K=�ߑ�S�'���:���P�k��>�)?��@�7��>!�?f�?�x!?=�C?�D?̭�=����4=�`1�>��>�v^��宿��r>�E?.�>�vL?H�?
++>	�?����.���w��=.">C�1?P�?�?w;�>�2?�޾���=��~>�Eb?%k�?�4�?g��>�\�>��*>��?���>�#$?NX?�6E?\Հ?:�M?f�X?�3`>�}�;�_����0�[���%�ݒ�5!�=��=f��.���*�<k�>�,u�	=O�=�>�F=?Qнq��}c�>=�s>3����0>v�ľN��w�@>�֢��J��
劾��:��׷=�>��?���>�N#�᳒=���>`=�>���37(?y�?�?-�$;~�b���ھZ�K�y�>�B?���=i�l�`{����u�Ƙh=y�m?�^?��W���F0i?O�\?����$+�$�Nl�	�b�9?�?N�:��>��{?�k]?Ee�>yEy��]��ٚ���a�^�����=h;�>�D�P@e����>�2?>��>�E>��>H�۾0o��qh��y9?K��?vf�?�z�?C�>$Tk���ڿ"�򾐊����g?Q��>�{��[�?��<����?���b־�;#b��]򍾌���R[B��G����mX=��?hSY?Fnd?�I�?~����u��a�a�p��Cu�z&��
�'dJ�_�D�5���b��A�Pa뾩�;j�����O�r	3�9�?�B2?*8��}�>�s�e����߾�>�j�.��<i��:ca�=�?�<�}ڽpX�;R&+?���>o �>�Q?��>�jlZ�>����C��c�=;$�>�Z�>� �>}�`:P�������q���HP�uܺ��X�>��Q?�$?�^u?|}�j�B��̀�zL$�8�L=��u77=�F�>p�H�������%W��}?��Im�Z�	��������E>�@�>�-�=�F�>�?�G1?�v��S�n�d�>���?�;E=ܑ�>|?��><{�>��>�����>��l?��>�8�>C���~h!�.�{��˽-�>��>֨�>pQp>��,�(\�ya�����9��<�=Z�h?�|����`��̅>PR?y��:2�I<p}�>�av�a�!����l�'��>6i?D��=��;>�>ž��>�{��,��XK"?޸�>��K��%����>ñ=?ZU6?���>��j?�G>����e�>p�q?��k?�o?���?Ds?��=��]��w��y�h��-<�i>���<{�*<o#��A��܃�q���S�<6&z�2�B>�p-��%M��=�r�<-e�=ja.>|��]�Z"
�o/�ٶؾ��Ո�ey���5��$u�qI����d�}�fx���Ͻh&P�K��-B׾E����?O��?��]��ۼ�H������"C�8��=Ȇ��Y��f5��6	��C��}�'�cľv�1��q��͂�	?m�Y�&?�H����ǿ�����h޾�7 ?<�?}�x?��P�!��8�d>7��<��FN�ٚ���ο����c`?�	�>B_�Mv��pg�>��>xX>Q|r>�S��A!�����<��?4�.?��>�l��sɿ�ͻ�3Z�<0$�?q@jmA?V�(�����NL=eF�>�	?��C>�-��*�^������>H��?�3�?�HW=�uV������e?E<��F�߿�6��=��=^�
=O�f�H>���> c��B�Sݽ�B5>�[�>=[�!���]�{H�<Z�]>��ؽ���5Մ?*{\��f���/��T��U>��T?+�>Y:�=��,?Y7H�`}Ͽ�\��*a?�0�?���?$�(?:ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=[6�^���x���&V�x��=_��>b�>��,�ߋ���O��I��W��=i��jҿ�/<���*�xz�=C��=��k�M�ݽ*���c��kAm�e����>#��=@�G>2I�>�5\>�6>ÞX?.�w?���>
�i>��;�	���luľvcR��x���R�"��eƒ�e���,j��iW��I�X1��I@�����1�<�Oď=a5R��\��FX ���b�.�F��^.?q$%>$
˾�M�Ё5<W�ʾW���Ǌ�v����̾ �1��.n�|��?��A?�څ�D�V���{�ַ�ވW?b����+w��Tw�=􎴼�=�0�>$�=F��3��jS�a:1?ӏ?ә����<)>Op��!
=̈+?=?��?6�>J�$?��+�z�׽r\>��5>�C�>F�>H� >
k���ѽ�i?q6S?�3�����p�>����v�$�j=nE
>a�8�:���([>��
=OŊ��+�����n�<�*W?瞍>��)����^V��lE���<=*�x?W�?^+�>�}k?/�B?���<�c����S����?w=��W?�$i?��>�x���о@�����5?��e?
�N>�kh���s�.��[��$?#�n?�\?Xy��o}����1��Oj6?\k?;�V�؟�[^�>W���Ջ>)��>�?�UL����>M?b!�����l�����=���?�@���?���=kn��l�=�?�\�>I�l�R?�=;���g��;Mi�>����Ri���hY��P�+?���?GN�>�����/��=����?/�?��־֝�a�/�I�n�!����=xj�=[R����Ѿv}8�qF�U(��?������<�>�@לS����>�:�X	ݿ�пm����ા�♾�k?tY�>h�,��Y���6b�"5����F�K8��Ј�)��>�?>=�������ܵ{��`;������ �>�Z�	M�>��S�m��� ���� =<��>��>�z�>�����ڛ�?����ο�����z���X?�w�?ty�?w?�A<8^v���{��$��mG?��s?�Z?��$�q�\�j6��@c?�꫾(f��v>��%U���:>8+?��>��8�ۛ=k(l>6��>5�=��,��ÿ`z���_��;h�?���?�p�~��>���?)5?#�eU���&��R3���=�A?	�">p ��_k'��O�������?ȷ7?*�-��C$�U�_?N�a���p���-���ƽr�>�0�W\�[�������Xe�X��H/y����?D^�?\�?2����"��3%?��>�����9Ǿ��<�x�>�&�>�N>:_�ҳu>��j�:��^	>���?|�?"g?���������]>��}?�L�>
�?7%�=as�>��=u���;�O�">N��=��?�>�?��M?��>��=��8���.�2[F��JR��)���C����>��a?FJL?8�a>�Y����0��� ��!ͽ�J1��V�@��,��߽^=5>��=>>6�D��Ӿ� ? �'ڿ�˜����o ?p �>Nf?����TV�\� >;?�\>��;�ߵ�𞙿v5��2�?���?���>�_־�J>=�H>\n>���=�Z�I�=�M���0>��Y?���pK��R�Y�։>6��?%�@��?� }���? ��"���
����i7����=2�8?Ҥ��d�z>]�>=��=�hv���Vjt�(/�>�?nr�?�u�>Ϊj?ԡn��@��k"=ן>[h?R�	?��������F>��??��d��"�e?��
@�-@��[?i���߿�.��J���*%۾��:>[��=��>'���i�=<=W�Z�����y >��>��>���>^Y�>N�d>(�X>#ہ�g< �,"��m���� #����1\�5�u���
�:	�����kԾ��S��4���|���Ƚ�µ�ܽU�>�|S?<�U?JZ]?8��>F�<��*>s��>h$>����\<&>��?i]8?β;?j��=�F��Jh��/q�?à�Ō/���>@��=~��>a�?'�>���g>4��>�ɞ>�yx=7�
>�M�<��=�JB>�5�>�<�>*e�>5O<>�>Rδ��/��G�h��w�x2̽*��?�|��L�J�J2��w6��)����t�=�_.?C~>����>пK����/H?u���&�f�+�%�>��0?sgW?�>���9�T��8>�����j��`>� ��|l�+�)�#"Q>�k?��z> b�>�`2�r�2�T�K�� ��:�j>i�3?�r�[��v�XJC���޾KqX>�R�>�&���a��>����A�q��Z�=�<?<t?7{���ʤ��B����?�S>.GX>��4= o�=�)g>�MQ�zTR�X�=���G=r��=d�a>�?^�+>��=y�>J]���P�Ȩ>��@>c+>�??��$?���]���0��܍,�69v>���>��>`3>4J��)�=B��>!�_>�
���x����ƭ?���W>�Sw��A`��a��A�{=����ϋ�=�q�=�����x=�2�=�~?|��䈿��]c���lD?h+?�=�F<i�"�P ��}H��X�?f�@m�?@�	���V�2�?�@�?�
��8��=�|�>
׫>�ξ��L���?)�Ž3Ǣ��	�P)#�<S�?��?G�/�mʋ�l�L6>_%?ܰӾ0x�>�����T�����s����=�"�>�]0?�|��_ g�*O�����>���>�g��T���z̿���(�>�g�?ne�?��G�6f��%U����>?�TR?i��>u�ھ������>�?^?�F^?�q�>�7*�7$����?I��?�;�?�N>JL�?�wj?��?��e�
IM�0N��;ۖ��l�=����f>"�>G࿾4u5��������h�j�eY	�)�3>���<��>�������f?>��<����!,;��A�>�|u=��Q>d?��>{˻>7Y�> �>a޽���FK��.K?�B�?�� ��R��b=%ͬ=$�f�?��=?rŽEoо�0�>��Y?LW|?��d?��>����K���U��\�ɾ�)�=�&�>Ǝ�>a�?�S�<�ˋ>�������[�>���>�4�4�v���}��>ѓ�>��?y1�>��>�	&?�x#?��j>[��>v�9�%]�L��j�>Z��>��?�)�?��?�Q���r-��ᑿ�⛿,%U��8>��l?Eh?Iߖ>g����s���C=≽X��ƒs?v1p?���� ?���?s�8?��6?�=>Lٽ�{��½�&�>�V"?���A���%��T�Ȃ?W�?��>=M�ٽv��'�����3?�#[?�X&?1~��%a�rľ��<G��ΣK��$�;�{m�I.>��>[�����=�D>��='Kn�ϑ6��y<7�=�Ñ>�T�=�D8������?�C'<�7��nqc��玿K�`���M>���>�k��2X?A�ƽmvj��A���n�����?�Q?n��?��?��=Сg���E?g��?�S?�u�>g�����L���ϼ�ky��,�ˈC����>#�Z���޾�y��𶿯�v�Jz���9q����>���>���>OD�>�ze>BW�>%f�J���V����E�e�+.���f�ww)�����=�?�>�{���Ex���>p�(���>׹;?�Q�>~z�>h��>M>���>�x�=�d�>�?4�>�æ>�E>:��=#:��NR?5���*�'������	$B?^gd?�G�>�h�������Zx?^}�?�o�?\mv>�ah��$+�'O?��>D0��7w
?ļ;=Q/�T�<8"��@$��T����6̎>t�ֽ�:���L��\f��
?f1?2��ik̾.�ֽ��������VO?7c<?;=�AX�2�f�8�o�9�Z���"�3T��l?��bv9���l��􁿬xw�⤀�I&4�V���l�.?�z�?����y2���!��\L��P]���=wX?#�w>�b>�
>�C�4X,���H�`G��_ʾ�K?�e{?�%�>5�Y?��??�[A?ʠY?��>�c�>��+?��I=��>���>��>?θ+?;�<?��?��?��(>�J�4&��9Ѿ�=?��?�]'?*O?^�?DC������f�=�U=Y�@�R޽�X�==v�<v��� F4��=�t>HY?$����8����Kk>Ԁ7?�~�>���>����-��D��<��>�
?�G�>�  ��|r��b�|U�>塂?^����=��)>~��=���*Ӻ�[�=V�����=�E��&�;�\<���=N��=#t����l�:2i�;�b�<�t�>��?ꑊ>|A�>�B���� �B��qk�=\Y>�S>�>gEپ�}���$����g��Zy>�w�?�z�?i�f=V�=ӛ�=�|��V�����w���'��<ߢ?HJ#?{WT?^��?��=?�i#?I�>+��L���^����b�?�,?A��>���[�ʾ�񨿋�3�͛?/Z?�9a����\<)�v�¾|ս[�>]/��.~����	D���������m����?п�?�@���6��k�N���M��֐C?B�>pQ�>��>�)��g�#��;>���>
R?�%�>�(Q?�[z?�#_?��O>��;�N~��m2���`�;Y	>[�=?�?�Ɗ?-�q?���>�0>�36���ܾl��K1&�����;��Hj=�fi>�D�>��>���>���=6��������[=��6�=5�d>��>ܴ�>[��>#Rf>���<��G?���>5'��M���q���#��tu:���u?x��?�k+?i=�q�sE�����f�>�o�?P�?�A*?S�S�-$�=��޼W붾�tq���>}Ϲ>��>i�=V+C=Q�>�p�>��>��_i���8��@O���?�5F?tm�=H#ſ�sp�����9�̀�����j�m�j��n�u���=�!���H�躾�ق����X���>Ǿϔ��
Ԍ�(�?�d�=��>��=��<Z�߼bb��P{s=�\
=�N=fR��C/Y��a��F	������3�ݲ�=坔<A¾+�o?@*R?�-?�2?i(�>(d >4���\�>E�;��_?��
>�K������t��A��G��?�����P�1����>���.>�Bb>�r>��d=]��=�"!=_*U=]����=
W>2�=�F�=�0>GH>�E�=�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>#:>�'> �R�k21���Z��c���[��!?��:��̾�F�>�*�=;}޾�OžW.=��8>l�`=����w\���=>�x�Մ;=x�f=�Ԉ>�[C>���=Xc��x��=F'B=y�=N>腟��4���(��3=LP�=��`>�4%>3�>e?�=1?�f?I�>|kr�ɂѾ���}W�>{��=��>�+�=�4>�h�>�4?�3A?��I?w̬>�;[=״�>*n�>#D1�&�j�6�ؾV���nA��?A=�?���>K��<CJ7��u�x>��[��Ft?�3+?G�?>�>X�c��hd&�8�.�OF���1�8R�*=Kbr�=�U�B��q�����=1��>���>��>�y>�:>��N>j�>��>���<���=ͫ��� �<�w��L�=	����8�<w�ż�Xo�M$�m�+�D2���}�;���;��X<���;�E�=���>��>˩>�7L<[�̾��*>A����H�I!�=�����+G���g�����~6�F�[�E8> p>9���Y����?� �>�m>�=�?�w?ɾ6>t�/��*���9��z�}�c��;�=�J�=�'*��6�H�j��J�n�þFڙ>R�>���>���=�R9��.K�]��=��Ծ�#"�+��>^���3� ��|������a��3�`�ı�="OQ?����y��=�?��T?���?�>?vb�<�_޾1r�>�J��|~�E$���4���\ ?Q%?7��><�ؾ��*�/f̾m�����>�I���O�ɻ����0��p$��ͷ�#P�>/��*�оH*3�Qk�����ՏB�n�r��к>j�O?��?,	b��M��=^O�k��l���l?��g?f*�>"M? ?Z<��1V��H��"�=@�n?=��?7�?'�>�*�=��<�B�>�o�>U�?c��?l�?�伽�j?&l�=���=�WY�>�s>Yuj>�Rl>�k>��	?��?S��>R2�ͭ��[���Ӿ��r���(=@��=���>� L>�?>���<V��:��>ՒU>X�}> ��>U�T>^)�>8Oi>���H|羦�)?J�����>�0?�x�>�f>�$>
E�>A����ˮ����oqýh����G��Ř<��\>��
>/8�>3ʿ���?%��>��d�>���_#s���>���>��,��>�\!>�P�>\�>�Ho>�Ni>x�I=`߷<����b�P=߾��	�q�J��0�6dܾC�N=�J���6�6��}���렾��k����i��M���96��u=��?2 ����a��%Z�}��=�!?V?�>�jS?v�Z�ި�=��=|C�>9!�>�\��'����E������ώ?�q@�9c>��>��W?��?��1�{3��tZ�s�u��'A�Je��`�����C���,�
�4��x�_?A�x?otA?��<j;z>̢�?��%��Ϗ�c+�>G/��&;�D6<=*�>�)��N�`�@�Ӿ��þ�4��FF>�o?�#�?6Y?�SV��xM�> �@?L' ?�y�?͛B?7�E?0e��B7?��>�_?$�?��4?��4?�A ?B�r>->���p�
=�����핾v��2�����<��=��>�5=@В�;3�=\!�p���r�4�?Ø=#T;=a&�=��=��=�C�=Ҧ>$�]?�7�>-��>��7?����o8�j���O7/?�n9=�܂����u���o��(	>U�j?��?9NZ?4d>g�A��CC�%>3Q�>;7&>*\>�`�>1S�l�E�fI�=xA>2>���=-�M��恾E�	��u��o��<�>P��>�@|>Ӎ��'>�k���z���d>��Q�{���r�S���G���1�%Av��a�>��K?0�?���=#[�Dd���?f�5%)?�W<?�FM?��?�+�=�۾`�9���J��(�h&�>z�<��Ӽ��o ���:��Z�:��s>i"��{⌾�>��C�](������\��uj��s>wf���=#+�*��Z4���>��>�玾E��*�����9�@?C�d=��<�������Ӿ�=ʝ>��>į��=�o<�5�+��=��=���>q�)=��!���n����X�>�YM?ǽL?ջ�?�L!�3S��"�1�k4�Ё���.^�V�%?l�>!�?�t�=MYU>�ʂ��d�+�Y�N.w�}T�>_"�>v���3�ؗ���� ��%%���>��?2�>���>��c?��>O�F?%�?E6�>{^�>�w[��/�0?I�?7��<j��<��콿�R�^Te��?jO?(%�~��>��?�%�>�C?.�`?�y1?�o>�/�Z�D��ژ>Љ$>��X��������>�g?֎T=��]?K��?r��>��?����򖞻,�>|I>h�a?��\?�}?ɬ�>x,�>�+C�ϲ�>��?��d?"~�?�[�?A��<t,?�cY=�R?:q����>'E?��?��\?��|?kmA?#b>�-)=�̽ߖ���x߽pD��c��Q��Ed̽_��������=�z�=�Ú�F����T����	=�<]r=��g�e��>�	q>�W���/2>vǾ�5���bC>���gP��W��p�>�4��=��|>8V?%��>S�"�n �="��>y��>F���'?oh?��?)X��M9c���ؾ�I�J�>_�B?)��=��m��_v�vu=%.m?�]?��[�$���N�b?��]??h��=��þ|�b����g�O?=�
?6�G���>��~?f�q?T��>�e�*:n�*��Db���j�%Ѷ=\r�>LX�R�d��?�>n�7?�N�>0�b>%%�=iu۾�w��q��h?��?�?���?+*>��n�Z4࿇G��]����V?���>&b�� )?)������q��-b���ԾT����Jپ�hW�`B���]�����Μ�B8Y>�!�>l)�?)u?��x?wﶾ��t��Ez�ֶ����M�iVE�;�-�T�M��xy�S���m�Sx����첾�u=:�P�A�n��?�'?@0�5��>�������~;�C>�t��e���r�=�����@@=o�Z=aih��e.��O��) ?�$�>�E�>��<?��[�-5>���1�~�7������3>�ݢ>K��>�B�>;�:+U-���G�ɾ�Ȅ��qӽէN>��_?6uX?�ۀ?%�G�5��Ps���!�����+�L$>_>ѵ�>V˹�Ugս ��_+�A�������u�ڏ���Ct��I?�l�>���=���?��?#���g���=şA�j�'>���>��?�iE?�L)=�jg�._f�ĺ�>.�l?u��>A�> ����U!�'�{��;˽)
�>��>��>A�o>��,��-\��m��؂���9��i�=W�h?�����`�{օ>kR?̄:��E<�>u�v���!������'���>G{?Ც=��;>Ytž%��{�u@��w�.?T�$?X�z���!�;��>%�%?�_>�q�>~�?��>�̰������<?y�[?��[?�Q?T�?���=�	���.
�-u��|�=�շ> Ԛ>��>�6�>D�^������'I�,J�n8>Z�'=$0Ž8�=O�ۻZ����S��r>T���c�3��@N	�`��|	��vz�n[$>H]���h�|���f�cr���#��7�.=�-���f��(v�N4���?�+�?_\��MR:������Z��USӾ���>�����g�_w��ľ=:G�$���I:��� ���&�r�M��_���<?����Ŀ�����]��9��>ˏ?�8/?�/�b˖���F���=�����f���E��@߿������T?F��>S8��4���>���>s�>I ��Ӝy�5ނ��0�<��,?�?u�?����vѿ����NX,>���?�k	@�|A??�(�����V=���>.�	?�?>�Q1�}I�����-T�>s<�?���?�~M=.�W��	��e?9�<T�F�w�ݻ�=�=�=�O=���ՒJ>�T�>����RA�x?ܽ۴4>�م>ȉ"����7�^�H��<z�]>v�սw;��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=lG��6ȿ;*&�^���=�����F_�%ҫ�*/����b�"X��{�Y����<Ku=/5�=W�O>���>%�T>��`>BZ?�ol?%.�>�s>u������	̾�dl<z7����2�Qd���[��H���L�4�۾+5	��#����u�˾�e>��k=�GT�;�����"���c���B�Ǳ1?6_>�fξM��4$=wEٕ̾���j�>���l�ɾ�E/�}�k�ן?flB?1���XR�^��'~I��E��U?	�3���ϭ�z��=���1=|��>�K�=[v޾��1��	R��y0?�?�.���d����->q���M=�u+? w?�n<�ͩ>1�$?0�%���޽��]>��6>��>,�>s�>�����ڽtc?�uT?.� �����ڒ>'���s�|�1�[=�>�D4�u��٣Z>�6�<�6�Q����<�W?L��>��)��%[��,��i�==9�x?q�?I<�>�k?��B?`�<wJ���S��$��~w=U�W?7#i?�>������Ͼ������5?8�e?��N>2,h����f�.��L��*?��n?3_?�2r}�s�����sv6?��v?s^�ds������V�b=�>�[�>���>��9�)l�> �>?]#��G������Y4�Þ?t�@���?��;<!�+��=�;?�\�>��O�?ƾ8z��������q=�"�>�hev����UR,�2�8?ؠ�?y��>`������g[�=:��?���?�V��\��< � ��if�+��Eҽ0=��]�&������.:�I�ؾh?�Ga��y�z=�Hq>�t@J�>�c��>�L+�#�ܿ5sϿ���]˾�־�g�>�>3��İV{�7s���>���L�.e{��9�>?�>9����ᑾ~�{�2;������>�b�k��>��S�ֵ������8<�ْ>���>��>T=��\�L��?�I��b7οڟ��=���X?#b�?�g�?Gd?a><l�v���{��j�KG?�s?LZ?��%��z]�'#8�" }?�����H��X1�i�V�X�s>a�?�@r>��<����>7�=i�0>&�=�B^��󷿂����>��Ra�?��?�߾��?W��?�u)?b�N�R��H�:��H���<?l4?��[>��¾�'��B��o���$?-C<?�E��!�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�
N�����Xe����@y����?N^�?i�?ӵ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>hH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�#�>��?�q�=
e�>�i�=��-�)k#>�!�=z?���?��M?L�>�U�=��8�//��ZF�HR��&��C�'�>��a?�L?nKb>4��K%2��!��uͽ�a1��E��R@���,�]�߽(5>W�=>�>v�D�aӾ��&?#�'�Fֿ-����Z'���/?�}w>U�?v���bB���缴!Q?��>���ǲ��؎��H2����?���?q�?E�ϾЮ+=M�!>�ҍ>בֿ>v뽉IF���j�'�B>Ң@?c@��I����i��F{>��?�@���?�*]��	?���P��Va~����7�d��=��7?�0� �z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�O�B���1=7M�>Μk?�s?�Qo���j�B>��?"������L��f?�
@u@a�^?*�m鿢���zо�<ھ�>?a�=��&>�������=�>ҕ�=�p��>�=H�q>�R�>�4�>W>�V>@_>�ɀ��2 �x�������*��B�����r#=5��$���=��hd�ѾH ǽ�� �fg	��/��dc-�$��=���=�EW?f�C?�b�?5*
?�7����=[1ھv��<��xkF>8R�=��*?�3?B�:?�8> ����(k�^�����i�D��&�>'�4>jB�>��>�ł>v�%�O1>��6>/>L�Y>,ۜ�wƼ��=v>�ٗ>���>��>��j>��b=K���d$��mB���kξ�:�=Mf�?k�Ǿ���T2��=˸�@��1 ;�.2?�$>WE	ٿ�{��zH?�+��G�ܾ��پ,�>a�S?��C?�k��OI�}v=�n�=��=����ru�%�������l���c>: ?+�f>�u>�3�\8���P�����y|>756?q鶾_=9���u�E�H��fݾMTM>ľ�>��C��g�����]�U[i��{=�p:?!�?�Z���갾��u�:��>R>dT\>C
==��=�TM>��c�m�ƽ� H���-=-b�=ș^>}q?>�*>�Y�=I��>����pP�땩>�@>�t*>�V@?��$?#4�qB��&����/���u>���>i��>��>cK��=a��>�c>��=^������@�v�V>ѻ����_�8�s�yw=���'�=��=����>�c'#=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ���>@���\�����z�u�W%=ە�>`�G??���d�J���=�L
?_�?"w�V����ȿ�v�zB�>���?aД?��m������?����>|�?��X?H�j>6�ھ[BZ�n��>�@?�?R?��>	G��'��&?�?���?zp�=2ڏ?.��?-8�>g`2��Y޾�7��(;��onɽ���0�
�(T=�g@�~0\�QQ���S����+�m�=����>���=�h>����.r��b�c1�M_E���:�o��>���>�>la�>d+?ছ>͊�>W?��d<�<)������K?���?��g$n�"��<��=p�^� ?`T4?��Z�^�ϾC�>��\?[��?�[?���>���E:���ݿ�J�����<r�K>i=�>}3�>���R�K>��ԾfD�'\�>}З>�:��/ھ�+���᣻�[�>�f!?�r�>C®=ٙ ?��#?��j>�(�>DaE��9��V�E����>Ϣ�>�H?�~?��?�Թ��Z3�����桿��[�f;N>��x?V?sʕ>a���생�kE�YBI�%���\��?�tg?}S�1?92�?�??]�A?�)f>ʇ�(ؾz�����>1�!?z���A�kL&����}?5P?���>�4����ս�8ּ���~����?)\?~A&?���,a�� þ=<�<��"��%V��
�;�uD�{�>ގ>؋�����=>�ְ=bNm��F6���f<Rk�=��>�=}-7�Mx���E-?F����0��{j�=F1w�C�0�>�.>��ž�a?�g;���|��𫿶����i��?�5�?tڕ?:���0mh�>?���? �?���>��C�Ծ�����z��|��_���>�Կ>.��!�4���੿N���Cҽ{9����>��>���>���>�i�>Ӌ�>���F20��x���Ǿ�g�li��y'��5�jj#�F?��.ޥ��f��վ��E���>f>g�Z�>UD#?��=>Eĥ>���>QN�<�*�>��Y>���>�O�>�h~>B�=	4$>`��=p�=��9R?����'�j��3���f7B??dd?�P�>xi�{����]�?΀�?�k�?kv>�vh�+�'r?uO�>���0V
?�>;=�����<�j������$���p����>N�׽�:�Y(M�uaf�Lo
?>0?x@����̾TC׽e��k�=��?Qx%?����E���v���Y��/T�&������榾x.��hv�}���Pӄ������"�!:�=��!?Cg�?�1޾z��<����	g�B�5�>�w�>��{>�ɭ>�. >]}�ˠF�#f��A%�+Y���>��l?W��>*�R?�1?9@E?K�q?X��>t��>xڰ���(?/�T=��T>|�>ɔd?=�>?26G?�(W?�f?�>x�Ľڂ������{�>?R?�Y�>���>;�7?k����Jn��\��vJ>8�¾^����Q>]G���$J�^�a=�W> P>�_?F$���8������j>U7?ep�>���>gZ��ο��j�<r��>��
?m�>� �7�r��r�	��>x��?%��˫=+�*>���=VL��a�[-�=����=�耼E:���!<���=�͔=�'t��'�796-;�ܤ;���<Iu�>��?���>�C�>�A��%� ���!a�=Y>�S>9>vFپ�}���$����g��\y>�w�?�z�?��f=7�=*��=}���T������������<w�?�I#?�WT? ��?X�=?5j#?L�>0+�;M���^�����b�?�!,?c��>�����ʾ�񨿯�3�ĝ?[?�<a�����;)��¾~�Խ�>�[/�j/~�����D�����:~����?⿝?�A�A�6��x������[��1�C?�!�>�X�>��>)�)�z�g�B%��1;>���>:R?Q��>b�O?�z?2-\?�oU>��8��୿�v��)�1���>�B@?�&�?}͎?͋x?�?�>ŭ>�*�����k��|�<j�n����V=�'[>��>�a�>�ͩ>���=�$ȽgG��b<>���=/�b>��>剥>"��>L#x>)Q�<�iJ?���>�h����d����k}�����v?Av�?je1?�T=�8��2-���Ծ��>''�?���?��(?P-u���=����Z"���풾�ھ>M��>i�>(�=Y�q=�w>��>��>�L���	��X/�3�Ľ�?�KQ?�Q >�b����a��
޾�ui�
�w��������_>�Ɖ�+�)*���)�>&�l�<�Ԇ��#[����<�]�I�����?��>���OH">�Ag�p����=1O����=1%>>�A�.��=��e��'\=��:�5��;1��<�o½�f˾P�}?%(I?��+?��C?M�x>��>�Y3���>񳄽1]?;6U>'lO��_���:�
c��0��(�ؾ36ؾ@�c�܍���>Y4I�R�>��2>���=�T�<��=�r=��=oi6��s=���=(�='ث=(��=TZ>/�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��>A��=N�V��(����-ă�ţL�h)?��7�ܢھKe>OH>L��X���*4=��1>��r=3i��W��$�=��?���'<㛍=�Q�>3@*>m�=�������=E�=g�=�V>�P\��J�B���e=;�=��T>se>#��>Mg?0?6De?��>k�r�W"ϾO���5��>�=I��>뙌=,C>7'�>P*8?�:D?��J?��>�1x=���>�=�>}�,��mm�$��O����<,U�?I!�?c�>�<G<�m<�����M=�}�ýof?�j1?�?w��>��m念\(�\-�]b���z���=^q"��s]�tk������:��f3�=ͦ>��>�H�>��Z>M8>��h>
p�>� #>قO����=u��h���6
��W> �*�0�%�Κ���}=�%�3��������/�[˵�6�h�vw>���>[p�=f��>o|�������i�>���r�Z���L>���J�Z�K�9���N�$~�3#�=�ep>#<T����?�m�=~��=D��?-�?��>�M�<w��蒿��̼L9D�� O>�[�>����[3�)9=�O.6�`��-��>odq>u�>qs>؟?��9�A�=����+<�5|�>�񈾵�н�)���}�>q���⚿N�b��=O|G?h|��i�(>�g?��C?�s�?C}�>�󘻍D;`>�К��-;=���x�?� ��;�y?_�?>��>�����#G�?G̾R���ݷ>�AI���O�_��0�E���ͷ����>������о$3��g������H�B��Nr���>v�O?[�?::b�WW���TO�����%��?q?�|g?Z�>�J?�@?}&���x�Rr���t�=��n?г�?g=�?O>ػe=W�C��p�>���> ��?��?)z?�]��/�>��(=9�h>��7">��A>Ն(=z��=~?�e?��?�^���3�A��#����D���T=��.;��>뜉>Ťj>�>���=�Ϣ=�,s>PO�>f�l>�iT>є�>�>����j�S�?�%��l>N�V?6u�>��'>�1b�5�>�� >]Ԗ��I=nS�;��\��5�g(�����>�UR>���>�jͿvE�?�>`���{�>�*��;>��>|�=h���Ut?	����;>J�>�V�>˜�=6x>)w�>�%ӾHO>
���}!��)C�,sR�wtѾ3dz>����ͣ%���A����GI��k���Y�_j��5���:=�'��<�?�?�1���k���)������?8(�>��5?���8����>��>���>vB�����G΍��w�&�?1��?1$c>�'�>)�W?��?�l1��3��}Z��u�$*A�Ye�x�`�sލ�O����
�|���_?��x?voA?�H�<�+z>^��?:�%�ԏ�[�>�/��);�;;=�-�>a1��8�`���Ӿ1�þ=��E�E>�o?w#�?�G?~VV��I�v�!>l�:?��1?h�s?�E6?B??8�Y�'?(h(>��?-c?��4?Ip4?9s?�L>R>s�<�?�<;#��E�����gM۽n�G�&� =?�U={�'��fR�k$=�F=S
��[{8���"�G��c#B<��G=��=���=Ֆ�>��^?=%�>]%O>)�9?pO�BC�$�����??�l�==�h��䐾�gp�A�Ѿ
�/>m?!#�?$$[?�jJ>	D�h.�	)>�?�>�J>@�>9�>a����L���O=4G�=��>^��=��.��i��}��Ε��r�<��;>���>S0|>,����'>Y|���0z�̤d>��Q��̺�\�S�Y�G���1��v�UY�>�K?��?Ɯ�=-_��-��?If�[0)?�]<?�NM?��?�=��۾��9���J�+?�q�>�[�<��������#����:�O�:$�s>�1������9�j>r�O�橾������b�3ƾ]>�>�Z)�`&y�>�H�d�ݾ���"N>�
>K�ξ9s"����Ź��ZO?=�>KQ��HE�I3�uJ�=љ�>RE�>S�+��?���P�S��XCS>�_�>{��=��<=����[�_��VC~>�M?��g?0��?�%\��s�����l��oA��5Su� O?.� ?��3?��>��h>�
U��CϾ�zJ��r��0�>���>��[ (����� 0��QE����>G�>@CY>-�>r�W?��>��=?��_?��	?���>������"?�l�?ƃs>>�=ց�(B�yXk��a ?��=?2y�Q��>��O?,m?�?�iv?�3<?���>��8Z��Y�>�U>�C�$���9�>G�Y?{�r=�\m?[��?��>	�N��-�1���o6�D�?=�c?��8?4d?g�
?���>����>�"�>kbB?_f�?a��?��	��;&?�5����$?��I>��?7/(?�?�Z?��v?��?���>P|=�%#�$b��$sw�����ƽ�ǧ=w_>��I=-粽Yl�;�l==R�<.7n;Vp��^���&F�%��=�E =�[�>,�s>�񕾽�0>�ľ& ��п@>����	A���늾�:��=^�>��?Ԩ�>�x#���=��>-i�>E��m,(?��?v'?a*;��b�n
۾	�K���>��A?���=@�l�2���_�u��{g=�m?*w^?��W��'��H�b? �]??h��=���þU�b����a�O?8�
?�G���>��~?e�q?Q��>%�e�-:n�&���Cb���j��ж=Lr�>NX�X�d��?�>z�7?�N�>_�b>t%�=nu۾�w��q��q?��?�?���?+*>v�n�Q4�
\¾����N�Z?י�>����L>?	?�������s�%kݾ]�־[u��c̾8�ʾI��x�y�@ia����;bj>{�>�<�?zn?gn?�ͧ�W�i�U�W��F����m�@��5J�&�c���i��uF�����\���T�K�V-��~���A����?�'?�0��+�>�Ƙ��K���̾;:B>�p��@��T��=�Ō�B A=�}X=g+h�ٛ-����� ?|��>��>�=?�[��/>���1���7����D�3>aޢ>���>ӛ�>��|:�0-��L�b�ɾ-ل�=rӽ��o>Z�t?Fc?�Q|?�j���k?�퀀��JN��h�=�D��>���=��}>!`$�U0@�9��74���x��41�]p��B�3���C?���>J��>���?�?_п�������=[�W��5�=y{�>/}t?,�;?fM�>o\�ړ����>�l?��>َ�>Fэ���!���{��˽!��>���><��>�Ln>�a.��\�8h��$x����8��;�={�h?�儾��_���>�1R?���9T	@<uע>���N�!��$�@�'�6�>~+?��=��:>�žĺ��|�6����)?�?����T*���~>i,"?���>��><�?F�>�g¾T����?��^?�8J?�]A?"�>��=/���7ɽ��%��l/=�>S�Z>��o=��=ʮ�B\�4�Zr>=S��=�м�ո�6��;̼��gJ<1�<��3>�ʿ)�M��B�Fd��Rƾϴ�؋�|4S=`袾���<1ھ�Tw�
ԾE���F�'<��B�l���`ԕ�Kf��L#�?j*�?O��j<�o��;�w�����
0�>�C���I���5��˓��|۾�U�0���+��CQ���v��v�r5N?N�h�x^ǿ54��U
���x?c@�>��?��^�پ�Y�`��>���ݛ��о?ڟ���l���z\?�J�>N	���cG��o�>�O?��c>#�=x���䃊�:��>%�?�,%?1'�>��^�^�Ŀ�ÿZ��=�N�?��@�yA?�(����v�U=���>`�	?��?>8L1��E�y���tX�>H:�?���?��M=��W���	��}e?-�<��F���ݻ���=�A�=[=�����J>GO�>�h�!VA�/zܽo�4>�ׅ>2b"����h^����<r�]>��ս�2��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=������ƿ@Z!�g���u�<�����<��W ������=����S�]��x4�}��=m�>JK>1]>�F>�IW>vu`?+q?� �>	�w>1�p2��
þD�<U����1��+��u�ཉ�ݾM��𱻾B��b����۾c�'��uu=�h��6���� �>h�?��%9?�Zt=���^4Y�~��;���'��ȧ��m�!��L�<��t��$�?��U?Cʖ�=C�@0��䆽^��J?z(��z(�0�Ǿ{b;=;ҽX�6=*R�>xg;��־�zD�<Jc�Ct0?�^?Mm���S���j*>�� �|�=F�+?9�?{�^<�&�>�N%?��*��/��z[>��3>��>+��>tE	>U��jM۽T�?_~T?��?�3�>����ֽz�9a=r0>"5� ��$�[>ő<k
��vAW�	��l�<�LU?O%�>9a)�����֎����m=��v?�N?T��>�l?��@?��<q�;�T����0�i=\\Y?l�h?B�>�5��%ҾԬ�Ef6?��h?C�Q>ERV����|/���6�?y�p?�?9L�ɑz��ꐿ��6?��v?s^�xs�����R�V�d=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�$Þ?��@���?��;< �X��=�;?m\�>�O��>ƾ�z������6�q=�"�>���ev����R,�f�8?ݠ�?���>������� >y�1���?y2�?
d{��hx=k!�Yeg�IC��s�}�����&�^�3����O��������_΢��׼�x>�@�n�����>�*&�[��ԓſX�������aj����>�N�<����mе�����2z��<T�?RQ�ež�7�>�>�ꔽ=D����{�+';�������>�}	����>=�R�,���p����-<���>���>�p�>꤬�w��v�?�����2ο�ƞ�Q���RY?�m�?���?��?:�?<- t���z���л�G?�Zs?��Y?�'��w[�"5�LV}?�*��.Z���X��2�8�����>T ?Z�T��K�>��|գ>����g���3����ޯ�rC�r��?���?�ﾼT?C��?�X?+]g�����G���/�v��>1>�W$>s���(���X�C��:?*U?l�q����]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?Ե�� #�g6%?�>d����8Ǿ��<���>�(�>*N>lH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?$�>��?�s�=kc�>�e�=U�p�,��h#>m!�=�>��?èM?M�>�Y�=��8��/��ZF�nGR��$���C���>��a?\�L?�Hb>!���2�f!��ͽ�`1��/��V@�Վ,�b�߽�+5>�=>�>g�D��Ӿ�: ?u���oؿls��? ��2?{��>�J?k_�!f����^?�e�>�����j<��
)�Z��?x�?<�?"�Ծ�:���=>�^�>��}>}ս� ��f9��:/1>~rA?4��s��y�n��>Y��?�k@���?D$f��	?���P��Wa~����7�y��=��7?�0��z>���>��=�nv�ݻ��X�s����>�B�?�{�?��>�l?��o�J�B���1=1M�>͜k?�s?�No���N�B>��?!������L��f?
�
@~u@]�^?({�ؿ�W��T�������=���=�^_>h뽱6�=�x����4�*�y�=�s�>v�]>�x�>D�4>�MQ>�&>����"��_���Ȝ��6��c��������>�������7��_�K|�������,m ���v�G�(��_����=u{Y?��W?l?��?���9h9>����=Ic�#>�İ>q�1?�C?k�?�0�=kl��(_�����l������K{�>��R>�p�>��>��>�_�=���;��> ��>\ >�)>��O=Õ�=nz�>��>6� ?�C�>j��>�{I>�;��r���������c�J�o��?-���0&�����:�������=�^?�S�=,�������ص���=?߿��N�⾁��;��>�F?�'?�.+>��Ǿ���=��D>�Fs��f[�@�h(��x��C�o�5�>��U?2�g>^Fu>n4��8�ʕQ�6[��=;|>�6?������9�Nv���H���޾��M>�{�>*�P��b�<��ԣ�bh�px}=��:?��?�����n��fht�g��o
P>߃]>t=���=��O>�+b���ƽ��F�%�*=���=%�]>�O?��+>c��=���>wU��
�O�~��>ًB>�=,>r@?�+%?QN��[��9p��*�-���v>�D�>�/�>��>VYJ�2n�=�b�>a�a>��I������?��vW>�<��_�GZu�`�x=]<��d�=�2�=J �R=���%=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ��>�1l��뒿�E��E�h����=ݭ�><?��ﾷѩ���⽻��>Ʌ?�Y�*t��jjƿPn�c��>�`�?�R�?aye�����)AQ�(9	?:N�?�?Z?���>�ើ��X���>��=?B�f?*�>��	�9��]I?� �?�l�?0�l>�\�?i2�?#��>X�Ƚ��J��%���;����T�P�ľ��=�0�|�����[��3������# |�}�$�徘=?1]<G�>�/,=D�S��� �"h�������	v?00�>�dC>�b�>Os	??�?�Q�>�b�=~{׽,����g����K?���?*���2n�"O�<W��=#�^��&?�I4?_k[�w�Ͼ�ը>�\?j?�[?d�><��O>��F迿6~��5��<��K>)4�>�H�>�$���FK>��Ծ�4D�ep�>�ϗ>�����?ھ�,���R��HB�>�e!?���>�Ү=9?g,?�Z>i��>�_D��ĉ�%V,�Jd�>&��>�`?X?x?�C?t۴���1�+Ӕ��A��8S��Kv>`}q?��?C��>Tk��%�&8�=�/�=Kp<��?�n?�I���*?hh�?�,Y?No`?�8e>������b�ǻK�>��!?��L�A��H&�:��~?UT?���>X����ս�ռp��@r���?�(\?IB&?��j)a��þ' �<�_"���R�y�;2�D���>�>�������=�>���=ZIm�*P6�?�f<WL�=�v�>q �=}*7����oS,?��.��?��?�=��s�BE��;}>1K>Q��B@^?f?��|�#1���ۜ���V�ux�?�8�?.x�?�#��c�h��)=?)�?�q?p�>�E����ܾ��� gv��?z�D�4f>��>�@��(�wk������)����aʽ������>�5�>�I?�K ?�P>�%�>�혾b�&�u��� �\t^�����8��/�����Ҡ��G ��� �Um¾��|�gV�>S	��c��>�O?Csh>�~>���>���L`�>pR>��>�g�>*�X>�S5>�>�}.<I�νE@R?�����'�n��9���A@B?Qud?�7�>��h�(�������y?_��?nj�?�v>�~h��+�z?�J�>K��BK
?C%;=�6���<6����������Mn�>��׽�:�t
M�(�f�4t
?�,?�i����̾d׽8}��y�=%C�?�)?�&�V\O�.q��xY��mT����F�s��c��+ )���r�����(F���<����(�Y�= )?w�?�Y ��쾜/����m��=?��\F>8
�>n��>��>�0>����0���c��+'����R�>��t?�Տ>4dQ?V?�<K?�?;�>��{>FG�/�F?��>~�>r�?C0I?.N?��<? ZT?�Q^?�>��؋��]���} ?�43?���>B�?��V?`1���d����Q=����[EA��b>��X={�b������=��>`Q?K���8�_#���k>L�7?C��>��>�#���Ԁ����<i�>��
?.�>^ �}�r��`�Խ�>��?ŋ��^=3�)>�{�=̼���&��\�=������=	��rK=�E(<�6�=P�= !h�W{�,v8;��;#�<u�>:�?���>�C�>�@��F� �g���e�=rY>"S>1>Fپ�}���$��{�g�~]y>�w�?�z�?h�f=�=T��=�|��`U�����4������<ģ?7J#?XT?W��?l�=?Uj#?/�>+�eM���^������?>",?��>����ʾh�ۋ3�;�?�[?=a����<)�Ɠ¾fսe�>V\/�B/~����|D�Uτ����)s��S��?���?�KA���6��u����hX����C?^�>US�>��>��)��g�R%��8;>Ԁ�>ZR?^׺>�cP?�h{?�]?TCW>�7�EX��e��Ds�j�>��A?���?�Ɏ?��w?���>v�>�_(��8������g���dȂ���[=��R>��>ד�>ڭ>+w�=q���.w����8���=�Hg>t�>�O�>���>��{>rAb<��G?h��>k��h_����4Ȃ�mπ�G�v?Xf�?�b,?S�&=����jE�G���i"�>GO�?���?��(?�V����=M[ռ�ͷ��v�6W�>�Z�>�-�>kv�=e�W=#>��>�>�	���xv9���V��?�2E?X��=J�ſ��s�~s�k:����<�!��=c��l���^����=�)��h�&��¤T� ќ�|ϑ� ܵ��ۚ�B#t��l ?�%�=��=C��==�cۼ@��<�yl=��A<)�=�k��4pe<�ԁ����Af�.b�;Y�<R�8=jj����˾ŏ}?�;I?�+?v�C?5�y>�<>6�3�r��>v���A?�V>ɗP�)����;�����9 ��Y�ؾ]x׾��c��ɟ�$H>�`I�_�>�73>�J�=�U�<��=8s=�ǎ=1�Q�d=%�=Q�=h�=k��=�>�T>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�7>`#>��R��1���\�M�b�~zZ�\�!?(I;��J̾�7�>��=^,߾l�ƾ��.=��6>>gb=�i��V\��=��z�=�;=��k=r׉>��C>�u�=�/����=�I=���=]�O>�����7��*,���3=,��=j�b>�&>�f�>��?�'6?��j?�>q2��/۾�δ����>��=��>��(>6;`>m��>�nD?@�F?��M?�̖>�ü���>[)�>�j$�]co���̾󶘾��Ľ���?�c�?�y�>�y˼_)�R�+� �?�$��K�?zN9?RN�>�v�>yZ�iLܿhU���M�����jԽ<Ø�e�Խxq���*>U�뽅m)�A$�=�>۴�>3j>�1>���=3��>���>���=��k=&�">�
�%�ٽ�Ea��!U>�?���#�>�W=�Q �X��=}�wg;z�g�͉���'���</ >� ?�>��>�70����W8/>�q˾�zL��R�=�����>�_�w������A�������W>$7g>%��
D��Q?W�=�Z>D��?��?w�>���Bj��������d<ϧ�8�>���>�n\��$9��S�D�B�|�Ͼ�r�>Sƞ>���>'`3>�M��FW���%;�)�O4�Q��>m���C��������8��bÛ�x�U�&9�=�C?�͇��p >�p?�oO?Ur�?܎�>4�v<�>	�T�1>_+��z=g	��x��=�*?I?P ?����H��G̾��1޷>|AI���O���G�0�8���ͷ����>���~�оI$3��g������:�B��Mr����>b�O?o�?�9b��W��UO�����)���q?�|g?��>�J?�@?'���y�^r��Zu�=��n?³�?b=�?�>���={����>_��>�+�?+��?.Y}?�:N��W�>���9�V�>kԽ2GF>�9t>0��=��>
!?]?�(?3���������ğ徜�h�q�o=)�&=Z��>�a�>/�>���=�[[= � >~pq>���>?�n>Vs�>�ѐ>�Bk>X�q��l߾��?q�����>;Mk?8��>�z>V򚽫�y��;���6%�5�<I�
�"�J�'��q�=���>K�E>gc�>8ۿ�x�?k	? ޾s?d4�h��=�j9>��:�
��I�>)M��i,��?|j�>��=��>��y>��Ҿ�>'��zt!��<C��vR�s�Ѿ�{>�䜾��%����#���\�I�����O�
j�#>���W=��,�<S?�?�0����k���)�Y����?�&�>��5?wь�e���Q>���>ȿ�>ؐ������͍����L�?���?�;c>@�>[�W?%�?��1�b3�$vZ�%�u��(A��e�`�`��፿;���m�
���	�_?i�x?�xA?�P�<�9z>}��?��%�ӏ�g)�>i/�5';��-<=K*�>�)���`�7�Ӿ�þ�8�PCF>��o?�$�?�X?(VV�Ե=+��9CE�>h�/?�P@?/C??�tw?z�-�e�;?���=��#?���>�bI?VQ?�?J��>�4A>�eE�餹�Cy�-�4�G��eN���C���{=Z�����Q;X｡�.<D��,�Qƌ���_�Cޕ��.ҽ"�=&��=��= ��>dI_?��?Z}�>�GO?�%��Z��.*��SQ?XJ>��+�w_%�����p۾Хp>^�?���?�<?��,>��S��B1��,�=�7>N��>�>�>�f�>����$i �i�>��=�̫=��}>[ּ����F�N�¾�q�=��>���>_,|>!��X�'>|���*z�٢d>d�Q�j˺���S���G��1���v�yW�>{�K?y�?ܜ�=�\龶"���Hf��0)?^<?}OM?��?�=I�۾r�9�"�J�@�#�>�9�<�������#��T�:�5Y�:�s>�3�� ���>�U��Hw�Z������^Z`����=p��Ḛ=6Q�T�6�����)�Ԁ�=,��M�q?���R���8?%�=Dv�ٱ �E��܁�+ʐ>{N>$*��᧽�^u�uHȾ��=I�,>YNU>�&�r)��{y�E��;,�>[??d"k?�ŭ?'�3������E��x׽6~� q�}�'?Fy�=�
?!�5>�D7>$�%��@���n�O���>�/�>7����=��g�r�־��n�4Pm>Q#7?��>��
?`��?�E�>��V??x?A	?~L�>C�!�6��%+?�I|?�(>V��=�"}=G�^�m����5?��8?�>�#�>��D?��>F6?7�?\}0?g�{><�
���V�;��>*?�>}�,ƿg��>��G? I�=��N?�>�?{��>��?��՗��Ղ�_&�=nC">hx?�C�?C!?x��>���>�ޔ�A�L>F۲>4�0?1��?o�?$�<�	�?��y>܉,?~��W�>��'?�j?a�@?4�K?�:(?ڈ>�M�=���O;�rg���=�b=zJ<!����潶E�=�T=<P<(4н�I!<,ؓ�]��O���Nz���t=���>�"}>
�Ͼ��%>ܢ侥i����<>D,
=Y���0z����j��0>�>���>h�n>�)����=�Ĭ>u�>�5���?�5�>�$?����lz�:����J��r�>#�@?k�<$�k����&Z�H=�e?�XQ?��K�V��:�b?��]?h��=��þ�b����P�O?*�
?��G���>��~?Q�q?#��>Q�e�,:n�!��Db�z�j��ж=6r�>\X�;�d��?�>a�7?�N�>y�b>T&�=�u۾��w��q��{?��?�?���?+*>a�n�W4�!x��Ѐ���O?��>W���{�)?�)�����b�����̾�վ��0S��C۾�6ؾ(S��S G����=ImS>^"�>�a�?}b?�x[?]����~d�3?m�������j�u-0���S���o���Z��]����@��1{��ξ�(����~���A���?��'?a�/���>���?���̾5�B>d#�����\G�=�����a@=JZ=�g��-�ޭ�F ? ��>o��>��<?c�[�/%>�Մ1��7�N���u3>���>P��>^<�>M��:`o-�c꽊�ɾ�{��ϛӽ[P�>}�f?�`?.��?��J�sJ!��s�� �DMĽ�P��V�=<���6�=@���UY3�M!���G�J�����7���H�^���o۽�6�?���>۽q��t�?��]?=�ܞ�{l)<��P�-��>�V�>� E?��4?��*>jA�=�`��6_�>�Nl?���><��>�捾�\!���{�^�н��>���>��>;m>M,2��]�h���">��	9�:��=�ji?�J��F�]�,��>
2R?��;��x<�ȣ>�Zw��|!��=񾔺'�Z	>�?0�=)28>�eľJ�e:|�
4��)?�?:7��C�)�,�>��!?З�>矣>�4�?q��>2c��6<�:?� _?ڥJ?�A?���>��%=񰳽�aȽ�J'��/(=�>n&[>�Tp=ѐ�=2��V\�n� �@=]��=`�Ѽ庾�Q��;%@��P�;<pD�<5>�A̿H������: ��o�ܼu�-(<=­u����E���xW��}��n���k�ۼɹl�.�B���]�D�_�?���?聩��v��yc����n����a�>��f�L�Ľ^;��_�)=����W��!���@�	�*�~�S�yHH�*�??ڶ��(Wɿ�ϩ�ɩ���?nj�> AV?C�3�[Sj��i����=����z���������ֿ�U���bd?�[�>*�ӡ���ۗ>\��>l8!>���=���� ���A&�-g�>�?]H�>�G���,�����`p��S;�?��@PfA?��(�Ws�8�T=�v�>�	?��?>)I0�(�tﰾ�K�>V:�?`�?��K=�W�����fe?��<��F��ջ���=���=a�=����I>��>����A�!�ܽ�3>lw�>�N#�����)_�]�<.]>�!ս����5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=���D{ȿ+������a�Mj��r�?��A��ν�HH6��������`;��Z>��>��+>Ʒ^>̄P>4�B>�k?�I�?oE�>q2)>�P ������*���={&/�U�"�󹄾�6��ؾu\�)�ɟ�l�����h�ľ=�4�ޞ�=�-Z��^����#��%^��:���1?Ձ>�(Ⱦ��G�|��=��޾t���w���JνQ%���`(�2@_�tC�?�H?����XI�����0��Gˎ��tE?�5�#8��\�V>jN:����<�+�>*ٯ=��ؾr�(��N���0?�?�8��Y�����4>���3L�<�,?��?Nğ<�ɩ>�`&?k�'��vݽ�^a>�{9>	٧>���>�v>���A߽
o?nuV?(����I����>�6���qv�)%7=Տ>��/� �μ��X>�1�< ӌ��f¼2���t�<R�V?�J�>vt)�<:��8��E"�ƕ?=��x?Mc?�Ԡ>�:k?;�B?���<�6��O�S��,�i5y=@�W?�vi?j�>L����оCl��5?�Ie?�/O>\]g��Z�@�.�(��>�?�un?�q?�'��΄}�	���uE���5?��v?s^�ws�����P�V�e=�>�[�>���>��9��k�>�>?�#��G������zY4�$Þ?��@���?��;<��W��=�;?m\�>��O��>ƾ�z������(�q=�"�>	���ev����
R,�d�8?ܠ�?���>������}��=�W��?~�{?���>��<��|v�<
�^��(�����:�㽝[��|P�6��	��F�����<�e>i�@TL=�A�>�����ۿ�Uÿ7쓿"��"���.�>�&P>&H�����\w���|�4{X�)�Q�$�r�##�>�<>�N��_(����{��0;��_���.�>����b�>G�S��赾l?���n.<42�><�> �>ᮽB����?r%��j)ο����z�o�X?r�?�q�?�}?��<<�9u���{��R��[G?��s?D�Y?&$�T2]�e8:�Xx?�ߘ���W�70X���D���=��>���>A�;�]�=^��IBg>���0b������Mt��\�/��h�?���?�T��	?�2�?�+?��2�x#���c}���0���>`��>�g�>������I��7�j�[�+F?�F?����I�]�_?+�a�N�p���-���ƽ�ۡ> �0� f\�N�����Xe����@y����?N^�?i�?Ե�� #�g6%?�>d����8Ǿ��<���>�(�>*N>iH_���u>����:�
i	>���?�~�?Qj?���� ����U>
�}?�"�>��?Gi�=�\�>_�=��۬,�Zo#>�"�=�>�ۡ?ҦM?�M�>�W�=��8� /��ZF�4FR��!���C��>Q�a?��L?bJb>���*(2��!��jͽ�n1��5鼩U@�T�,�ߞ߽�.5>H�=>�>z�D��Ӿ�0?�5��aؿ?����'���3?�N�>��?lY��Jr��I��V^?�)�>����0���[��Pt�d��?�6�?c�?
;׾9"��	>8>�>��>tNֽ�����S��83>�nB?��$��/p��p�>I��?�z@�	�?*h��	?���P��Ta~����7�j��=��7?�0��z>���>��=�nv�ܻ��W�s����>�B�?�{�?��>!�l?��o�M�B���1=.M�>ǜk?�s?iQo���e�B>��? ������	L��f?
�
@}u@^�^?+��޿0R��`̾�&پL 
<2��<HnR>եν�%=X��=RTx:F:���>z�>йj>Xo>>�P>��U>_>�ą��!��9��Gx��:�N��&���ɅH��N��U��_#��d��fM����� �����M#�E~;��2@�q�=}�U?�R?�Ep?� ?�0{�Rx>�A���� =�+$�|w�=k��>P]2?k�L? �*?�$�=<Ý���d��o��y-��9҇�hm�>}I>,r�>$�>��>)�:.YI>�F?>K��> |>��(=����A=(aO>[C�>��>�c�>ܛH>�<)>� ��Zy���v�W��������۞?����UYF��f��X��<ž�Vm=�(?��=���^\Կ�a����D?�����=��5U��$>S7?C�B?w>�⻾ҧ>��g>�7��F���>k���痾Uw-�0�>i'!?`g>>�u>��3���7�,kQ�/����|>�	6?�L��&b9�PMv�*H��!޾�hL>|N�>�|S�Mj����;3�h��{=�g:?9?+���WS����v����\gP>�\> }=���=��M>�Oa��{Ƚ�~J�H1(=?#�=~_>�n?>�P�=�J�>������A�7��>��Q>�$,>��=?��$?쟼mK��vƅ��.��j>���>O%�>�>T!A��4�=��>F9f>s��é���k��?��]T>�5}���j�QT����p=�#�����=��=�O��2�0��=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾrS�>�1�5Ȗ�=��>�r���h=���>1H?,���:.ͼ�1���?��?SP���Dǿ��s�f��>||�?&��?�:j�2��D����>T��?L�[?qf|>��ʾB�\���>;?1T?���>v��;��y?ެ�?f:�?H�9>Q�?�R�?�|>@�;�����͐�۵������ᬾ�.>T����V���W�Ꙣ�ە��T���B��j�>^�F=�f>H�l�_s�J�)�I�a=�6���p�=%C�>���>��}>���>l�>Ҋ�>XU	?�L9>+ 5��� !����K?���?-���2n��N�<Z��=)�^��&?�I4?k[�}�Ͼ�ը>�\?k?�[?d�>=��P>��G迿7~��G��<��K>*4�>�H�>�$���FK>��Ծ�4D�cp�>�ϗ>�����?ھ�,��[S��GB�>�e!?���>�Ү=- ?��#?'j>,��>�%E�8����E���>�D�>%�?{c~?��?�G���c3�v,��%���AD[�#�M>*�y?o ?6��>hv�������h-��:������҂?[�g?D��O8?���?[_@?�B?غg>XY�d�־#/���M�>~�!?D���A��L&�B��?�S? ��>�&��-�սP�ռ����u��(?J'\?�?&?���"'a���¾>�<�#�MW�"��;��D���>��>`������=[>�԰=dRm�hJ6�JGf<�i�=�}�>��=B*7��y��>,?�GG��ڃ�ט=�r�sxD�İ>2L>��*�^?Bt=�~�{�����z���!U���?i��?	l�?z���>�h�C%=?H�?�?�!�>�>��[n޾	�ྮVw��nx�v���>���>mk� �X�������|H��D�Ž�"����>�׽>��>u��>��u>�>��}��f!���Ǿ뾸�Z��R�1O2�U8��E��袾 ����q=��;��~�K�x>���c��>,�?�i�>"Q�> �>�1^����>�4>툈>Q5�>8��>j#�=�W>�.�<����GR?�����'��辙���#1B?Znd?�7�>i�����p���?y��?�o�?+v>)~h��(+�p?WB�>����n
?5%:=x'��$�<k[��$��M����=��>ir׽f!:�!M�_{f��c
?+?g��V�̾Nf׽������=��?�2$?6*!��I���n��b�l�W��5 �n���F��SL*�Fpv�YY��Q􇿘ۂ���!���=A"?���?��Ҿ���p���h�&�1�	� >��>�q�>x^�>�>3�����[��/-�E���]��>{x?B��>� L?!.?��x?շ�?C�b>��D>F����?�?��Y���t>���>\e?�B"?��G?L/s?��l?�>�>������0澜�Q?�O�>}��>�?�
>?>aҾ�Q��k
=�R�=�v��Yά=�5>�n���g5=�}��{��<Qd	>~?�ݽA�2�5E��F>��=?1��>���>W����bZ���=-�>b?^��>Y.��t�!>����>n9�?g�#��&ϼ?< >�E�=j�l�f��<�t�=!5C����=�j�P���+�<(�I=��z=X:�=���J�=s �<n&�mu�>�?-��>�B�>�A��\� �����`�=�Y>S>�>&Fپ-~���$����g��[y>3w�?�z�?�f=.�=���=�{���S��&��	���V��<f�?�I#?�WT?���?Q�=?�j#?ͷ>=+��L��N^��|����?`,?%�>u�X�ɾ�`����4��?�)?�Na�[�p�*�����Sh۽}>�.���}��گ��VE�����5�r䙽w~�?�Ҝ?P�6��Y5�"�W��V��~ C?���>� �>���>�(���g�8^���7>���>��R?L�>��O?�5{?>�[?eT>F�8�����ՙ�Z�1���!>$@?���?���?_ y?E��>,>��)��ྪO����{f����,V=e�Y>�{�>4!�>���>Ҕ�=<�ǽxz��4?�`\�=�Sb>�p�>�s�>	��>�Cw>�k�<miI?�}?�}�����:5�����4�����?A�?�X?��=�����5���¾���>��?F|�?:�%?�|�����=�Z-=��ľ��	f�>���>H��>	��S�=�X�=k�>p��>�����GH�c~�v�? �[?�!)>���� �W�:٨��g���x�����;�O����<�y_���=�������<�ɾLJ��:����7��k����GQ���?x>����gp�=��l0����=��i<會�u�J=D7
��5=0����k;�����<�'�{[=��#��˾��}?�;I?ʕ+?��C?x�y>�;>�3�P��>*����@??V>�P�̈��v�;�;���| ��&�ؾx׾�c� ʟ��H>�`I�"�>�83>XG�=MM�<=�=�s=�=��Q��=�#�=�O�=.g�="��=�>
U>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>w2>��>]V�=�1�-�h�"Pf�YV���!?�89���˾7�|>� >�9�bg��I�={+>�qW=*���W���=9�D�nz�<���=7a|>V+>�,�=x'��{*�=ub=�@�=&�H>	�,�pN9���q�`�N=6^�=�_>�M>c�>��?�e0?Ed?�@�>�n�0�ξXq��_�>�=�߱>H��=:D>�4�>g68?)�D?��K?�5�>�Ň=a��>!��>/�,�s�m�����ç���<Ԁ�?ҳ�?
6�>i�M<0�@����a	>�֫ý�3?/91?s?~��>�������Q@���B��e�L~Ľc�=_�ռG�G��5���ߘ���i= J>j_�>��>B��>��b>��=�k_>���>Qǝ=H���b��=2w�.�9=�k���)>� �<�K�=����l�Ē�j=�=LO�<N��<U��O��;�h =P_�=��>K�>lq�>� B=�'���'>�ȕ�aK��Y�=� ��!�<�W_��*��k�7�&S@�0�)>��d>E6;����D?�US>��">���?��z?��c>}#���dξd���.�TMG�KB.>|fM>N?8��0:�0U��nP��Ⱦ[��>�פ>�N�>[�>��0�����ۤ:l㾈�.�ɤ�>\*������zv�7�����������Y��z>f�v?�����<>ks\?�&?yB�?:�?��>��/��=W�(��zS>�ھ�`>bȊ>i��>o��>Q�>5���X��D̾��bշ>CI�X�O����0�zB��η�Ϗ�>g�����оo$3�nf��������B�Nr���>
�O?a�?�7b�(W��QO����-D���q?�zg?V�>J?H>?�2��y��v���q�=��n?)��?<�?��
>�ȴ=��L�>E�?3h�?���?6�o?�˅�u �>G�輈Y>Z`���	W>�
`>8 �=�!D>��?�6?>, ?-�ǽ:���

��I
�����r�<Q��=�V>��>K�H>7�%>��>���=*��>���>��)>D�=G�>z�y>�萾%���?����t�>SbP?5��>�Xv>|>S���ӽ$�=�������s%U�l
.��v��� =�*>9P>���>�?ѿ���?(U�>T�����>_�u�~=�X#>q��=;vd��d
?P��<��S=>��>0��>e/]>0��>��Q=�Vb�!27>�k)��s$�	�_�S\����5vg>�-��c��
F�1>��:
����¾|�����s� ���d|��B��{Ӈ?Srz��/\��Z�P�>*jr?��N=�?O����9>-��>z/�>nȾ>�� �sQ�������I܊?r��?�;c>c�>|�W?�?&�1�H3�
vZ�h�u�k(A�9e�\�`��፿���D�
����F�_?g�x?jxA?�X�<�9z>E��?��%�wҏ��)�>�/��&;��=<=�+�>S*����`���ӾԹþ46��HF>�o?�$�?9Y?tUV��=@>]���?lR?a�M?�o_?�$}?�C��~�?�q�>�,^?�>�c?�Uc?�!?]�>���>�1>Ę������:�6IȽ5��� �x�_�:=�w�=�/�;�=�H<��-=��=_��!<	���u�^�=�Dk=.��<�}�>�Gh?�q�>��X>�\?�Ad��VT�M���a?�i>�NS�:���?�^�T��	�>u y?+ŷ?��[?�>x4G�ҷ>�	@�=��>؊�>_1�>Y?�D��!I)�cz�R�H=0�k>�F>:d�9�W��["��q��;N��>���>�.|>����'>�|���/z���d>��Q�\̺���S�]�G�Z�1�҄v��X�>q�K?��?��=�]��)���Hf��0)?�]<?�NM?��?�	�=)�۾N�9��J�r@���>C>�<�����$����:� ��:��s>�2�����>�>Κ@����TϚ������z:��P>),;�l��=ɫQ������ﾌ+�Y��=7���-�^1��������C?yAϼ
9�<W㩾4Ծ<C >���>�8e>L����3W�ԝ"�;���G>&�q>e��=B�
=���z�K�9����>�F=?+`w?@��?%:M�Hyi��<�L6�������d>I�'?*�>].?_X~>ީa>W�������&�*�o� ��>	��>m"0���J�/ �Cn�y�o�?��>��>T�>� ?�?���>�j.?-@#?�!?��\>��c;��n�-?��{?��S���U<��<D�]��z���2?�?V�4>��>=�6?h�?-'?6�o?�<M?L�H>��پ$Q@��b�>	1�>����䯸�E��>�(?Q�P>!��?�f�?=V��#;�X8������F��>��~?��f?�?!��>EѨ>��^��>;2�>��I?���?8_s?���=�!?�B��?[Ǥ�w�>��O?'�3?�wI?��~?Iw.?Q}�>�+����m��&ͻ���r@�	O�:EJ)�vg�=Ӟ����=���=u\;=������������=�O�e� :ü���8X�>��s>����0>K�ľ�?����@>'䢼�L���Ŋ��`:����=�v�>;�?s��>�y#�籒=ϱ�>�S�>~���$(?��?�??%;��b�۾xK��&�>,B?���='�l�����u�h=��m?
�^?��W��'��O�b?��]?@h��=��þ{�b����g�O?=�
?2�G���>��~?f�q?U��>�e�+:n�*��Db���j�&Ѷ=\r�>LX�S�d��?�>o�7?�N�>/�b>&%�=iu۾�w��q��h?��?�?���?+*>��n�Z4࿹~ƾ'��:P?g��>yz�� ?�󁽪}���9��>�a��p�$��歾�̾���^r��Y��I��'t^>@h?�B�?��?N�]?Rپ�l�AX\� ��(y[���<�� 4�k�}��C�@L<�,�{x��<<�쏼��a3�͵|��@@�'��?K�)?�t/����>�w�����&�ξtlD>08���*���=%ㆽ��I=��Z=�h���-��N��s�?�Ը>�	�>e�;?$[�n9=�5I2�[E6����f�2>Ӣ>v�>V��>���:W�-���ʾ�Ё�OBӽjW�>�o?L}?��?�"��)/���}��-#��:���©����=�R�Z��=׵�vK��W�$�@�4�����&���}��"� >����?}~>��X>箥?}��>��	i<q;,>�C�(>s��>@�?�d6?�9�>/[P������>�l?�S�>B�>���P!��{���̽���>G��>���>��o>�-�H\�xz�����#9��Q�=��h?⪄�EC`�>�>MR?��%:�vH<hf�>�z���!�-�򾖀'���>�i?f��=�;>�dž� �\�{��`��!)?�c?�J���*�s|�>�"?���>���>�B�?P:�>l�¾���9+@?��^?�QJ?�A?�s�>�S%=������ɽ±'�y�1=0�>�~X>̊s=�J�=!��X�]�~���G=��=xtۼ�����<��ƼJZ<& �<��3>�Ѿ�ʔF����+��"I�@���:�$' ��E��b桽j�ྪ�J��,��ܷ��F<�A@�/�%������d*����?M��?�|��C=�ȗ��m���v��V��>�¾k�U> �!�*���
��n��(�ʾ0&��e/���T�׺W���A??����ǿ���� ��.�?��>\2?E7�%�q�	�K�1�㽬<]�8+t�yn����(�ῥů�B-?7��>k���W|T��>�Њ>�@p>��$>�Ⱦ픾R�޼ղ?��?�ǭ>����%ǿ�
��h��<���?^@�hA?��(�/��S(T=N�>Ε	?%�>>P/�|��ㅰ����>�S�?/��?P�I=csW�C�	�=ne?[�<�mF��ػ'�=��=Fj=N����J>�N�>s��6FB��wݽ��2>�>��"�(5�O�]���<�j]>�Xֽe0��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=�� ���ſ�`"��{"��7<1R��ʐW�� ��&��yŴ�W���y�T��vʽ�=���=F�[>5w�>J�N>	�`>4�]?yg?C��>�@>[Ͻl�Qľگ�<R�������s��U�A��"o���ǾW^��g�F���ξ�X�:�dю=�U���t�"�Կd��HC�� /?�>�þ�O���<pξ����x��dd��s�ɾ��1��dl��à?�]D?�܅��>T�݁�Z�L������OV?с� ��s�����=�M�{}�<y�>!��=��⾡�2���S�_1?Lc#?��Ⱦ��~��V�>������4?�z?�(��;-�>M�-?Ҙ�kzܽ�d�>��l>���>�#�>.�>������-w!?ՓJ?/&��:�w�>��ʾ���8,=���=�q1��%��H`�>��.=�]����~=��S�9=3V?��>��(�������M����<��{?��?�c�>xg?�F?b.=P��f5N�U=���=�GX?� h?�4>pВ�2mɾ����|�2?�ed?��S>��w�����.�|��x?q(n?g�?�kϼ��|��琿����T5?��v?s^�vs�����E�V�j=�>�[�>���>��9��k�>�>?�#��G������xY4�"Þ?��@���?[�;<��@��=�;?p\�>��O��>ƾ�z�������q=�"�>���zev����R,�e�8?ܠ�?���>�������|>:�I�+֧?�ar?l�|��o�<W���]���µ�&�R�ctA������� K�U����&�x졾^N�<4�[>�@��=��>�E2�d�ۿ�p���덿��þ��=��>i��<E�㽂瀾�˅�Zu��:<Q��W���־P�>-�>�����5��U�y��<���C��>h�wW�>�L�?<��!�����b<,�>bD�>s��>1뭽��\`�?����8Ͽ�M��4���V?&�?IC�?�!?��.<#x�T�{��=��E?>t?Ӊ]?M����8^�.�+�Z+u?ⳇ�{�i��G>�^ra�C�>�
?9�=��6��LG=Ֆ
��e�>6K���b��Aǿ�ʨ�V��^��?��?�d�j�?LÐ?�A?��Q�������g��u5�UEX>��>�>�>S4���=��W-�j����R?��m?��g��/��]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>gH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?f$�>��?�l�=Fb�>�`�=��,��k#>� �=��>���?��M?GK�>�U�==�8�f/� [F��GR�{$���C��>��a?L?�Jb>V��&2��!�xwͽ�d1�@Q��W@���,��߽
(5>��=>>��D�\Ӿ_�?�o���ؿOj���x'�+34?޵�>��?���J�t�����4_?o�>�:��,��&���^�d��?�F�?h�?�׾��˼�>�׭>vC�>��ԽD����w����7>m�B?L��C���o���>/��?j�@^֮?��h��	?���P��Va~����7�X��=��7?�0�3�z>���>��=�nv�ݻ��V�s����>�B�?�{�?��>"�l?��o�K�B���1=9M�>ǜk?�s?�Po���n�B>��?������	L��f?	�
@}u@]�^?&�3߿Du���A̾�^۾PM=5.=�U>u^	��1�=C��=�r=۩R=�
�=̓�>�/5>Gc>*�_>h�
>�H8>���r��hS��`政�!E�`5"�x�^�z�g�h|��Pu��댾�㠾��������׳���Q�%���?>4S?�O^?eh�?�!�>=���2F>����SC���g���=�r�=��4?3C?V�-?NB�=$a��]�8���/������Ҽ>�T>쯿>j�>���>Z��=SbP<7�+>�B`>�>P�e>�F=0;V<%�>>څ>!�?`>B�>c�]=�䦿P����y��󻷾�mֻ�:�?d\
�����̪��x{����s�¼�C?���=�B�����'���HO@?:(���W��z�7�>��g?�?��=�����*>��=�僾#El�p� >W�_��!��L�<�>�9?�Mg>�u>�H4�Rk7�~Q��ϲ��}>G
6?�I��[�6�� v���G� ޾�J>�_�>nH�< ������~���g���=`�:?Q.?�)������`u�ν��K�P>�X>�=
ݨ=�LM>,�m�"�Ž;oG��(&=�y�=һY>?j�>�0�=���>�S��1}/�s�>��l>6->܋D?-!?��<	����P��Tz+��Y>6�>�s�>6�$>u6��3z=���>�	x>��üC|�������V��K?>�B��(G��q�,�-�l=���!r>��=���D�7�P28=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�g�>ol�HY�����R�u���#=լ�>`5H?�Y��)�O���=�rr
?�?_�G�����ȿ�zv���>��?S�?��m�?���@�Љ�>���?}fY?�i>\_۾�ZZ����>�@?�R?�'�>05��'��?�޶?���?�g>�^�?���?�P>�*o���*�=���:���c�(=SϜ�݂��Eо��Ǿ����V��񘝿\��/���ᅽ��;G��>��=���0���B5\�� ƾ�dL�^�>%�>�>�J�>���>�	?i��>h��=�<=�����龃�K?���?-���2n�CO�<[��=.�^��&?�I4?�k[�}�Ͼ�ը>�\?j?�[?d�>:��O>��E迿8~��7��<��K>*4�>�H�>�$���FK>��Ծ�4D�ap�>�ϗ>�����?ھ�,���R��DB�>�e!?���>�Ү=˙ ?��#?��j>-)�>�`E��9��U�E����>��>hI?@�~?��?-Թ�=Z3�����桿x�[��;N>U�x?�U?�ɕ>r����tKE�HI�J���p��?�tg?2O�?=2�?]�??'�A?++f>��dؾ���� �>m�!?��ϺA��M&����~?�P?<��>�6��S�ս�Aּ���Z����?�(\?HA&?����+a�E�¾A:�<��"�_�U��
�;]�D��>�>l���'��=>Q԰=�Om�G6�a�f<�j�=��>��=�-7��u��6=,?x�G��ۃ���=��r�xD��>iHL>��g�^?�l=���{�����x��P
U�� �?Ġ�?3k�?	��*�h��$=?�?]	?"�>�J���}޾���0Qw�o~x�tw�F�>���>�l���$��������F����Ž$}���?�l�>�L�>�I�>Փ>��>y��u�&�0�۾��¾OXh��/	�M##��v<���"��#��h�Ƚ��%=��ؾ	S���>���I��>ǚ	?��A>,��>"8�>s|a���>_eC>/�>���>���>��>_�>y@|='-ν�HR?����-�'�G�辙����5B?krd?p0�>Fi�͇��|���z?%��?�r�?))v>�h��)+�.p?KC�>r���i
?�\:=��Z�<X�����M������%��>�H׽�:��M��nf��l
?.?����̾4@׽v�����=oY�?y(?�0(���P���o���W���R��D��n��j���U%��q�dX���ք�g���=�(�ы/=3K)?���?� ����Z����k�b">�s\>fZ�>�@�>Z0�>d�<>���9�/��F_��'(��Ӄ�{��>�zw?�\�>�P?zH?r�F?�Do?��>"��>wz�[:)?0���/a>�b?�d]?{�:?��F?$�B?�f?��>s�=���~���	9?�|�>��>A?�p??�ɽ�Q�̲s��HV=�[��,��H��>�I�<
��e^�QY�<d�U>Z�?%=�ތ7�O����bl>-�7?#��>�z�>�_��Q�v�S��<*�>��	?e�>{���<r��
����>j΂?u���<�.>���=ցi�2��%��=F����=�=����%7t�84_<
��=�5�=��.�9`�:�?�]�;�_�< u�>6�?���>�C�>�@��/� �c�� f�=�Y>=S>|>�Eپ�}���$��v�g��]y>�w�?�z�?ջf=��=��=}���U�����H������<�??J#?)XT?`��?{�=?_j#?ϵ>+�jM���^�������?�(,?j}�>�����ʾ�憎�3��?P:?�=a�x���;)���¾��ս1>�n/��/~���� D�O�p���������?ǻ�?�B��6�)U辺����E��zyC?��>�a�>���>h�)���g�����;>΄�>nR?V��>��O?s�{?��]?��S>Ժ8��:������[�a��%>L�??�|�?��?��x?0F�>LE>M�)���S����=�7]���쁾�?\=@LY>�>M��>��>M]�=�1ǽ���Y=���=��c>�_�>�D�>a�>P8|>n��<D>K?ۊ??�־*���@н�b¾�=��W��?��?&'!?_��=M�о=��Q�,9?��?f��?3#?Z�E�*^�=�U�<%���2�W�#d�>�A�>��>%
�<�o>�8����>��>�K���v*�Q�4�)���L�?\�L?��>��ſ5�q��5q������c<>s����d��Ȑ�P�Z���=D���b�����vi\�i��ຓ�Z[�����L�y�J
�>�N�=���=��=w��<Cռl�<K�E=r�<�=�&z��Vv<B�9��Z�P��}���*�L<?G=�򻴈˾ƍ}?E;I?V�+?��C? �y>:C>��3�嚖>ؑ���@?�V>�P������;�2���-����ؾCw׾��c��ɟ�uE>}cI���>�:3>qH�=5Q�<'�= s=��=.�Q��= "�=�K�=�a�=���=Q�>`T>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��7>�>�R��1���\�+�b�@|Z�ˠ!?�E;��9̾�2�>N�=+߾8�ƾ0�.=^z6>�xb=�`�N\����=w{��#<=�Bl=T։>M�C>�]�=�T���ζ=�gI=ȅ�=��O>'%����7��,��3=q��=īb>�
&>}��>dR?�F/?
m?0�>S����@����o>��U>�;�>�+>�F>���>}�<?X!D?N�@?�Ѯ>9��<K��>���>��A���y� ��^]����
�R!�?�s�?@��>ՔE<*w-��#�ֶ7�����.?B�9?��>\�>����Jۿ���3DG�g
(�\X=� �=۩��k�=a �=��=u<ۺ7�W>8Z�>G2f>>��=�b�>���>���>�J�>V�>�2z=��t=��ڼ3�|��Ր��P�<�<{��Ї�ݰ9���<A�1��|ühu=Η=J1;��4O�K�Ż4�=���>�>
��>��u=q���@�2>�\���_M���=?����oA�6�e�A(����1��v<�̹=>�T>��Y�X���^�?p�_>�~4>�!�?��w?bZ,>������־���NT���Z��S�=�)>̠7��:���]���J�AvӾS��>*��>��>b<�=!�T�����Z>�(@��A��B�>}�=�H�������'��򕿉�K�P����d?�ݒ����>P�p?U��>au�?lg3?�L>���v=�����1�>d/'�: �>l�>��
?&��>V��>�W����<��̾RD��_��>�I�F�O�ַ���0��^ �j���>�����о�*3��j��@ ����B�:�r���>��O?+�?��a�>D���:O����~��Uy?�jg?�.�>�.?�5?�;��v���r��J�=��n?y��?=�?o>@d�=}<����>��>P;�?�ٓ?F�u?�+�m��>��+<sbv>����=,�B>n�<�Ix=��?v?��?��ǽ#��@ྊ���OH�`��:�,<�l�>���>ro>�K�="f�=��r=,M>���>?B�>�`>d�>%w>������?�>���<�>cPD?N�q>C2�>�6��`�6>�>%ս�/���hi� %��Y��?�>�e)>���>+3ݿ�?��s>����hث>��$�E>ͳ`>L>�Ծ:�9?�/�=��̽I�?�y�>�>��)>�Z>��Ǿ	�>:r��(%�&B�
&O���о��x>��3���������S�]f���k��Rh��D��&@�|�vҎ?br�/n��u*�H���LH?Z��> �.?�7R��&>H��>���>����ཕ�̀����1ύ?B&�?�;c>��>O�W?�?��1�+3�	vZ�'�u�k(A�Be�_�`��፿����
�����_?��x?yA?DS�<
:z>]��?��%�Pӏ��)�>�/�';�1><=o+�>,*��+�`���Ӿw�þ�7�_HF>i�o?/%�?UY?�TV�����v�Q<30?IU�>�E?�Kq?��l?�v\�m�)?�����~$?g@�>��#?qFZ?�?���>�K�>�^>��Q��F���i�>�۲ʽ�`Ǽ)��=v��=؅2��Ճ���I=��槽�౼�&=e����ג�<uz�<J���Bm�>�h?��>̔>�Kl?���W�q��d*=:�q?�0̽;�:����Z/<=!��T�>!�?;>�?_f?�I>�d��L?���>��n>���=��>"��>�o��a�O�R��|�� �=���>��>��ɾb�4��q{�O7�=��d>���>�1|>�����'>�|���2z�2�d>��Q�κ���S���G�6�1���v��Y�>��K?0�?i��=_�9��SHf�}/)?�]<?�MM?��?��=��۾K�9���J�d?�X�>*o�<	��e���{#����:��ݛ:��s>�2��{⌾�>��C�](������\��uj��s>wf���=#+�*��Z4���>��>�玾E��*�����9�@?C�d=��<�������Ӿ�=ʝ>��>į��=�o<�5�+��=��=���>q�)=��!���n����X�>�YM?ǽL?ջ�?�L!�3S��"�1�k4�Ё���.^�V�%?l�>!�?�t�=MYU>�ʂ��d�+�Y�N.w�}T�>_"�>v���3�ؗ���� ��%%���>��?2�>���>��c?��>O�F?%�?E6�>{^�>�w[��/�0?I�?7��<j��<��콿�R�^Te��?jO?(%�~��>��?�%�>�C?.�`?�y1?�o>�/�Z�D��ژ>Љ$>��X��������>�g?֎T=��]?K��?r��>��?����򖞻,�>|I>h�a?��\?�}?ɬ�>x,�>�+C�ϲ�>��?��d?"~�?�[�?A��<t,?�cY=�R?:q����>'E?��?��\?��|?kmA?#b>�-)=�̽ߖ���x߽pD��c��Q��Ed̽_��������=�z�=�Ú�F����T����	=�<]r=��g�e��>�	q>�W���/2>vǾ�5���bC>���gP��W��p�>�4��=��|>8V?%��>S�"�n �="��>y��>F���'?oh?��?)X��M9c���ؾ�I�J�>_�B?)��=��m��_v�vu=%.m?�]?��[�$���N�b?��]??h��=��þ|�b����g�O?=�
?6�G���>��~?f�q?T��>�e�*:n�*��Db���j�%Ѷ=\r�>LX�R�d��?�>n�7?�N�>0�b>%%�=iu۾�w��q��h?��?�?���?+*>��n�Z4࿇G��]����V?���>&b�� )?)������q��-b���ԾT����Jپ�hW�`B���]�����Μ�B8Y>�!�>l)�?)u?��x?wﶾ��t��Ez�ֶ����M�iVE�;�-�T�M��xy�S���m�Sx����첾�u=:�P�A�n��?�'?@0�5��>�������~;�C>�t��e���r�=�����@@=o�Z=aih��e.��O��) ?�$�>�E�>��<?��[�-5>���1�~�7������3>�ݢ>K��>�B�>;�:+U-���G�ɾ�Ȅ��qӽէN>��_?6uX?�ۀ?%�G�5��Ps���!�����+�L$>_>ѵ�>V˹�Ugս ��_+�A�������u�ڏ���Ct��I?�l�>���=���?��?#���g���=şA�j�'>���>��?�iE?�L)=�jg�._f�ĺ�>.�l?u��>A�> ����U!�'�{��;˽)
�>��>��>A�o>��,��-\��m��؂���9��i�=W�h?�����`�{օ>kR?̄:��E<�>u�v���!������'���>G{?Ც=��;>Ytž%��{�u@��w�.?T�$?X�z���!�;��>%�%?�_>�q�>~�?��>�̰������<?y�[?��[?�Q?T�?���=�	���.
�-u��|�=�շ> Ԛ>��>�6�>D�^������'I�,J�n8>Z�'=$0Ž8�=O�ۻZ����S��r>T���c�3��@N	�`��|	��vz�n[$>H]���h�|���f�cr���#��7�.=�-���f��(v�N4���?�+�?_\��MR:������Z��USӾ���>�����g�_w��ľ=:G�$���I:��� ���&�r�M��_���<?����Ŀ�����]��9��>ˏ?�8/?�/�b˖���F���=�����f���E��@߿������T?F��>S8��4���>���>s�>I ��Ӝy�5ނ��0�<��,?�?u�?����vѿ����NX,>���?�k	@�|A??�(�����V=���>.�	?�?>�Q1�}I�����-T�>s<�?���?�~M=.�W��	��e?9�<T�F�w�ݻ�=�=�=�O=���ՒJ>�T�>����RA�x?ܽ۴4>�م>ȉ"����7�^�H��<z�]>v�սw;��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=lG��6ȿ;*&�^���=�����F_�%ҫ�*/����b�"X��{�Y����<Ku=/5�=W�O>���>%�T>��`>BZ?�ol?%.�>�s>u������	̾�dl<z7����2�Qd���[��H���L�4�۾+5	��#����u�˾�e>��k=�GT�;�����"���c���B�Ǳ1?6_>�fξM��4$=wEٕ̾���j�>���l�ɾ�E/�}�k�ן?flB?1���XR�^��'~I��E��U?	�3���ϭ�z��=���1=|��>�K�=[v޾��1��	R��y0?�?�.���d����->q���M=�u+? w?�n<�ͩ>1�$?0�%���޽��]>��6>��>,�>s�>�����ڽtc?�uT?.� �����ڒ>'���s�|�1�[=�>�D4�u��٣Z>�6�<�6�Q����<�W?L��>��)��%[��,��i�==9�x?q�?I<�>�k?��B?`�<wJ���S��$��~w=U�W?7#i?�>������Ͼ������5?8�e?��N>2,h����f�.��L��*?��n?3_?�2r}�s�����sv6?��v?s^�ds������V�b=�>�[�>���>��9�)l�> �>?]#��G������Y4�Þ?t�@���?��;<!�+��=�;?�\�>��O�?ƾ8z��������q=�"�>�hev����UR,�2�8?ؠ�?y��>`������g[�=:��?���?�V��\��< � ��if�+��Eҽ0=��]�&������.:�I�ؾh?�Ga��y�z=�Hq>�t@J�>�c��>�L+�#�ܿ5sϿ���]˾�־�g�>�>3��İV{�7s���>���L�.e{��9�>?�>9����ᑾ~�{�2;������>�b�k��>��S�ֵ������8<�ْ>���>��>T=��\�L��?�I��b7οڟ��=���X?#b�?�g�?Gd?a><l�v���{��j�KG?�s?LZ?��%��z]�'#8�" }?�����H��X1�i�V�X�s>a�?�@r>��<����>7�=i�0>&�=�B^��󷿂����>��Ra�?��?�߾��?W��?�u)?b�N�R��H�:��H���<?l4?��[>��¾�'��B��o���$?-C<?�E��!�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�
N�����Xe����@y����?N^�?i�?ӵ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>hH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�#�>��?�q�=
e�>�i�=��-�)k#>�!�=z?���?��M?L�>�U�=��8�//��ZF�HR��&��C�'�>��a?�L?nKb>4��K%2��!��uͽ�a1��E��R@���,�]�߽(5>W�=>�>v�D�aӾ��&?#�'�Fֿ-����Z'���/?�}w>U�?v���bB���缴!Q?��>���ǲ��؎��H2����?���?q�?E�ϾЮ+=M�!>�ҍ>בֿ>v뽉IF���j�'�B>Ң@?c@��I����i��F{>��?�@���?�*]��	?���P��Va~����7�d��=��7?�0� �z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�O�B���1=7M�>Μk?�s?�Qo���j�B>��?"������L��f?�
@u@a�^?*�m鿢���zо�<ھ�>?a�=��&>�������=�>ҕ�=�p��>�=H�q>�R�>�4�>W>�V>@_>�ɀ��2 �x�������*��B�����r#=5��$���=��hd�ѾH ǽ�� �fg	��/��dc-�$��=���=�EW?f�C?�b�?5*
?�7����=[1ھv��<��xkF>8R�=��*?�3?B�:?�8> ����(k�^�����i�D��&�>'�4>jB�>��>�ł>v�%�O1>��6>/>L�Y>,ۜ�wƼ��=v>�ٗ>���>��>��j>��b=K���d$��mB���kξ�:�=Mf�?k�Ǿ���T2��=˸�@��1 ;�.2?�$>WE	ٿ�{��zH?�+��G�ܾ��پ,�>a�S?��C?�k��OI�}v=�n�=��=����ru�%�������l���c>: ?+�f>�u>�3�\8���P�����y|>756?q鶾_=9���u�E�H��fݾMTM>ľ�>��C��g�����]�U[i��{=�p:?!�?�Z���갾��u�:��>R>dT\>C
==��=�TM>��c�m�ƽ� H���-=-b�=ș^>}q?>�*>�Y�=I��>����pP�땩>�@>�t*>�V@?��$?#4�qB��&����/���u>���>i��>��>cK��=a��>�c>��=^������@�v�V>ѻ����_�8�s�yw=���'�=��=����>�c'#=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ���>@���\�����z�u�W%=ە�>`�G??���d�J���=�L
?_�?"w�V����ȿ�v�zB�>���?aД?��m������?����>|�?��X?H�j>6�ھ[BZ�n��>�@?�?R?��>	G��'��&?�?���?zp�=2ڏ?.��?-8�>g`2��Y޾�7��(;��onɽ���0�
�(T=�g@�~0\�QQ���S����+�m�=����>���=�h>����.r��b�c1�M_E���:�o��>���>�>la�>d+?ছ>͊�>W?��d<�<)������K?���?��g$n�"��<��=p�^� ?`T4?��Z�^�ϾC�>��\?[��?�[?���>���E:���ݿ�J�����<r�K>i=�>}3�>���R�K>��ԾfD�'\�>}З>�:��/ھ�+���᣻�[�>�f!?�r�>C®=ٙ ?��#?��j>�(�>DaE��9��V�E����>Ϣ�>�H?�~?��?�Թ��Z3�����桿��[�f;N>��x?V?sʕ>a���생�kE�YBI�%���\��?�tg?}S�1?92�?�??]�A?�)f>ʇ�(ؾz�����>1�!?z���A�kL&����}?5P?���>�4����ս�8ּ���~����?)\?~A&?���,a�� þ=<�<��"��%V��
�;�uD�{�>ގ>؋�����=>�ְ=bNm��F6���f<Rk�=��>�=}-7�Mx���E-?F����0��{j�=F1w�C�0�>�.>��ž�a?�g;���|��𫿶����i��?�5�?tڕ?:���0mh�>?���? �?���>��C�Ծ�����z��|��_���>�Կ>.��!�4���੿N���Cҽ{9����>��>���>���>�i�>Ӌ�>���F20��x���Ǿ�g�li��y'��5�jj#�F?��.ޥ��f��վ��E���>f>g�Z�>UD#?��=>Eĥ>���>QN�<�*�>��Y>���>�O�>�h~>B�=	4$>`��=p�=��9R?����'�j��3���f7B??dd?�P�>xi�{����]�?΀�?�k�?kv>�vh�+�'r?uO�>���0V
?�>;=�����<�j������$���p����>N�׽�:�Y(M�uaf�Lo
?>0?x@����̾TC׽e��k�=��?Qx%?����E���v���Y��/T�&������榾x.��hv�}���Pӄ������"�!:�=��!?Cg�?�1޾z��<����	g�B�5�>�w�>��{>�ɭ>�. >]}�ˠF�#f��A%�+Y���>��l?W��>*�R?�1?9@E?K�q?X��>t��>xڰ���(?/�T=��T>|�>ɔd?=�>?26G?�(W?�f?�>x�Ľڂ������{�>?R?�Y�>���>;�7?k����Jn��\��vJ>8�¾^����Q>]G���$J�^�a=�W> P>�_?F$���8������j>U7?ep�>���>gZ��ο��j�<r��>��
?m�>� �7�r��r�	��>x��?%��˫=+�*>���=VL��a�[-�=����=�耼E:���!<���=�͔=�'t��'�796-;�ܤ;���<Iu�>��?���>�C�>�A��%� ���!a�=Y>�S>9>vFپ�}���$����g��\y>�w�?�z�?��f=7�=*��=}���T������������<w�?�I#?�WT? ��?X�=?5j#?L�>0+�;M���^�����b�?�!,?c��>�����ʾ�񨿯�3�ĝ?[?�<a�����;)��¾~�Խ�>�[/�j/~�����D�����:~����?⿝?�A�A�6��x������[��1�C?�!�>�X�>��>)�)�z�g�B%��1;>���>:R?Q��>b�O?�z?2-\?�oU>��8��୿�v��)�1���>�B@?�&�?}͎?͋x?�?�>ŭ>�*�����k��|�<j�n����V=�'[>��>�a�>�ͩ>���=�$ȽgG��b<>���=/�b>��>剥>"��>L#x>)Q�<�iJ?���>�h����d����k}�����v?Av�?je1?�T=�8��2-���Ծ��>''�?���?��(?P-u���=����Z"���풾�ھ>M��>i�>(�=Y�q=�w>��>��>�L���	��X/�3�Ľ�?�KQ?�Q >�b����a��
޾�ui�
�w��������_>�Ɖ�+�)*���)�>&�l�<�Ԇ��#[����<�]�I�����?��>���OH">�Ag�p����=1O����=1%>>�A�.��=��e��'\=��:�5��;1��<�o½�f˾P�}?%(I?��+?��C?M�x>��>�Y3���>񳄽1]?;6U>'lO��_���:�
c��0��(�ؾ36ؾ@�c�܍���>Y4I�R�>��2>���=�T�<��=�r=��=oi6��s=���=(�='ث=(��=TZ>/�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��>A��=N�V��(����-ă�ţL�h)?��7�ܢھKe>OH>L��X���*4=��1>��r=3i��W��$�=��?���'<㛍=�Q�>3@*>m�=�������=E�=g�=�V>�P\��J�B���e=;�=��T>se>#��>Mg?0?6De?��>k�r�W"ϾO���5��>�=I��>뙌=,C>7'�>P*8?�:D?��J?��>�1x=���>�=�>}�,��mm�$��O����<,U�?I!�?c�>�<G<�m<�����M=�}�ýof?�j1?�?w��>��m念\(�\-�]b���z���=^q"��s]�tk������:��f3�=ͦ>��>�H�>��Z>M8>��h>
p�>� #>قO����=u��h���6
��W> �*�0�%�Κ���}=�%�3��������/�[˵�6�h�vw>���>[p�=f��>o|�������i�>���r�Z���L>���J�Z�K�9���N�$~�3#�=�ep>#<T����?�m�=~��=D��?-�?��>�M�<w��蒿��̼L9D�� O>�[�>����[3�)9=�O.6�`��-��>odq>u�>qs>؟?��9�A�=����+<�5|�>�񈾵�н�)���}�>q���⚿N�b��=O|G?h|��i�(>�g?��C?�s�?C}�>�󘻍D;`>�К��-;=���x�?� ��;�y?_�?>��>�����#G�?G̾R���ݷ>�AI���O�_��0�E���ͷ����>������о$3��g������H�B��Nr���>v�O?[�?::b�WW���TO�����%��?q?�|g?Z�>�J?�@?}&���x�Rr���t�=��n?г�?g=�?O>ػe=W�C��p�>���> ��?��?)z?�]��/�>��(=9�h>��7">��A>Ն(=z��=~?�e?��?�^���3�A��#����D���T=��.;��>뜉>Ťj>�>���=�Ϣ=�,s>PO�>f�l>�iT>є�>�>����j�S�?�%��l>N�V?6u�>��'>�1b�5�>�� >]Ԗ��I=nS�;��\��5�g(�����>�UR>���>�jͿvE�?�>`���{�>�*��;>��>|�=h���Ut?	����;>J�>�V�>˜�=6x>)w�>�%ӾHO>
���}!��)C�,sR�wtѾ3dz>����ͣ%���A����GI��k���Y�_j��5���:=�'��<�?�?�1���k���)������?8(�>��5?���8����>��>���>vB�����G΍��w�&�?1��?1$c>�'�>)�W?��?�l1��3��}Z��u�$*A�Ye�x�`�sލ�O����
�|���_?��x?voA?�H�<�+z>^��?:�%�ԏ�[�>�/��);�;;=�-�>a1��8�`���Ӿ1�þ=��E�E>�o?w#�?�G?~VV��I�v�!>l�:?��1?h�s?�E6?B??8�Y�'?(h(>��?-c?��4?Ip4?9s?�L>R>s�<�?�<;#��E�����gM۽n�G�&� =?�U={�'��fR�k$=�F=S
��[{8���"�G��c#B<��G=��=���=Ֆ�>��^?=%�>]%O>)�9?pO�BC�$�����??�l�==�h��䐾�gp�A�Ѿ
�/>m?!#�?$$[?�jJ>	D�h.�	)>�?�>�J>@�>9�>a����L���O=4G�=��>^��=��.��i��}��Ε��r�<��;>���>S0|>,����'>Y|���0z�̤d>��Q��̺�\�S�Y�G���1��v�UY�>�K?��?Ɯ�=-_��-��?If�[0)?�]<?�NM?��?�=��۾��9���J�+?�q�>�[�<��������#����:�O�:$�s>�1��٠��Wb>0��v޾�n��J�ɹ��@M=���UV=g�8־o=��d�=�
>~����� ���֪��,J?�kj=�f��LXU�Im����>H��>�֮>=�:�*Zw�n�@�����N�=���>e;>�����w{G�04�L��>�JJ?��e?��X?�F��B-���Y��������\����8�?�>�7�>˨&>�m=�	��w9����9�Z��>���>�G+��!c��侱����'��p�>�!?l=a�V?$Pf?�e?�N?iQ@?��*?���>���<[=��{{,?��?u��=	>��S���*A��^m��M ?�m!?���w�>RC?]� ?�E+?�[V?���>�Q�<�7�i�:�|U�>n3�>R�{�F���%�>�zS?�s ?�l?~�f?%H�=d�<���Ƚp�<Д>��}>��=?8� ?`.?]�>��>�����r�=I��>
c?�&�?6�o?��=�?�|2>(��>��=���>��>???O?_�s?#�J?�p�>iݍ<���C���=!t�F8O���;t�J<��|=�~��+t�^���<l��;w����<����W�C�.���!��;=`�>��s>����0>i�ľM��5�@>�S���N���܊�ׅ:��=)��>��?.��>�W#�%��=y��>�C�>����2(?�?	?B&;�b���ھ߾K�9�>�B?���=S�l�*���+�u�;h=��m?��^?E�W�$��^�b?�^?BJ�Z=���þ��b������O?-�
?�H�Z	�>��~??�q?��>�se�%n����*Eb�$�j�ɶ=�>fx��d�tO�>c�7?��>UMc>���=Xt۾��w�����$??�?���?���?R*>،n�������'����]?9��>."��� #?qx�ڦϾ�������O�U��nF��+�������$��僾HG׽�`�=]�?$�r?nq?Ⱦ_?7 ���c�O�^����.�U����dw�A�E��E�w!C��1n�D��/������T�F=t�ȓA�'��?о'?R0����>ڲ�����%;2C>����o�%A�=;^����?=ƜZ=�mh��o.��[��y ?�!�>Q�>W�<?��[�}2>�I�1���7�&���Yu3>�ʢ>挓>�H�>�:k7-��M�ɾ_���_�ӽ:mw>GKc?yeK?��n?e� ��I0��Q���Q �A>�q����f8>KT>>p�>�Y�� ��X(�?��vr��$�5q���'	��j�=�93?�܁>s��>(��?A(?om
�O����}���0��v<i��>�g?,`�>Tу>��׽��!�B�>�e?e��>�#z>z�O�S��`����Ι<z�>�ޞ=�"4><��N����R��e��V���2@��:=ͨi?V]�mH&�K��>3�?:����=:��>�{�=. H�#�K�������=�@'?�56>a%>��q�,�m�����|)?�2?6��*��C|>�,!?�D�>
��>U΃?��>�'¾sK�;�N? �^?C�J?��@?a��>�=݋��".ʽ��%��*=¦�>xa^>H0v=:0�=�]�\�p��8C=ԁ�=�������`�#<0O��q{k<b�=04>	Oҿ13M�����R��������o�G�	�����x�|������nj[��d���y=8O8���9��X�יe����??�?b�WsȽ�S���.��b�m��q?�����ͼM����h����e�-���j 7�*^��XN�Α>�C�'?+����ǿŰ���;ܾe  ?B ?[�y?���"���8�ͮ >6A�<G6��5��њ����οB���4�^?��>^�2��Y��>a��>��X>�Hq>���1鞾�<�<Y�?C�-?��>��r�_�ɿ;���aͤ<���?:�@}A?��(����mV=��>/�	?J�?>�S1��I������T�>I<�?���?�xM=��W���	��e?�{<�F��ݻ��=�<�='F=���˔J>yU�>���SA�ZAܽ��4>څ>'}"�_��ւ^���<�]>[�սI;��NՄ?_z\�mf���/��T���S>�T?w,�>F/�=n�,?7H��}Ͽ��\�)a?/0�?���?��(?Eֿ��ۚ>��ܾ��M?�F6?���>c&�t�t����=^c�Vऻ����(V���=K��>��>�,����ދO�H������=�_��oǿ!����2��>J��!$�h\3�����M������c��j]S���ɽ�*�=2,>��b>@}>�L>��X>��U?��u?�b�>Ec���H��	��$8ž�g��Y����`i��8|�@�νx����ž�R־�z�O����[�׾�.=��}�=�/R�^����� �"�b���F�[�.?�c$>�˾��M�=.<�aʾ��������	����'̾�1�en��ʟ?�B?��	W�"��������8�W?�y����pାb��=@J��s>=�><`�=����3��zS�͐0?�� ?���ç��.\'>u���&6�<l�,?�P ?ԓ�8^�>&�'?���G�˽+j>'�/>T��>���>��>7�����$�?��W?���K���q@�>Kؿ���q�M̃=�>M�6�Ԗ��t�[>K��<�n���9�����Uü<p(W?4��>[�)�1�,a�����tO==X�x?l�?�,�>�zk?[�B?�Ԥ<h��2�S���]w=u�W?�)i?�>����/	о����5?��e?4�N>�`h����.�.�U��$?C�n?�^?�|���v}�c��n���n6?ݑ�?�{]��r��@<�t5��!�	?V��>�;??�]�d
�>o+Z?�'��������s<�VB�?y�@�N@�||=��`<�t=�#?vͮ>�f��� .��n���8>��6?%��7����;���>�yD?Zʑ?(��>YX�ж���=Nٕ��Z�?y�?P���Cg<z���l��n���}�<̫=d��E"������7�@�ƾ׼
�o���"⿼å�>-Z@�T��)�>D8�G6�TϿ"��a[о�Sq���?��><�Ƚ[�����j�^Pu�L�G�R�H�����gN�>��>��������B�{�)r;�P����>����>��S��%��ՙ���5<%�>��>�>~0��J轾�ę?^b��?@ο?������t�X?&h�?o�?�p?kv9<��v���{�g�n.G?�s?�Z?2i%��9]���7�%�j?�_��wU`���4�tHE��U>�"3?�B�>U�-�V�|=�>���>g>�#/�y�Ŀ�ٶ�?���Y��?��?�o���>r��?ts+?�i�8���[����*�D�+��<A?�2>���I�!�B0=�SҒ���
?V~0?{�f.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?!7�>�2�?|s�=�c�>8��=z�����)�e�D>":>䔜��.?S�R?�X�>zg>1`�m�(��.C��N�� ���A�$�k>5�b?�&X?b�>z
��wuѼF\#�jyy�IH��F$V<(BS�I~(���n�=>��>>&O/>��"�$Vʾv�%?~�����2熿�vپ1d/?�
�>:?��!��H-��X��h?Dd>@����b���)X�:�?e�@��?g���Q�<�?�<��>�?�J�=���A��)��=e�N?lț�l�����j�6��>�=�?��@tU�?d�i��?���\a��m�o�D/-�c��=�T>O�Q?����H>�>pqQ>�{��	��lˀ��V�>J�?DB�?�W?5Xc?QS����-s���Z�>�o?�w�>*Fݼ�`�eX(>~8?�������s7��B�o?M3@��	@{Ӂ?����ۿ���?���@7Ծ�1�=�*>F�Z>63��[�=K����<�>�;U�;>[�>]�>\}x>l,b>~�S>��9>go��_*��蚿$���"3�c�#���A�.�׶��V92�q��&�Ѿ����6�~�;�ּ�f�����7=�-�=KT?!�N?��v??�r�-�>	KȾlB>m=�mF&><Ǿ>s,F?�O?M&.?G��=�����T]�^U��GW��G�|���>��W>غ�>*��>-��>0��<FFR>MX>T�v>A�=/#=v5�<c��:*>bc�>;�>�֤>�C<>2�>6ϴ��1��\�h��
w�t̽0�?X���[�J��1��S9������fi�=Tb.?
|>���?пW����2H?����)���+��>��0?�cW?B�>!����T��9>���=�j�`>z+ �El���)��%Q>sl?|h>'r>�A1�Q88�@0O��奄��>�14?[���	O<�y\t��K�?�޾�W:>���>zmk�y���֕�:%�g�i=�;?Ą?N���8h��l{������R>emH>LQ�<G��=r8L>*&S�tE���tH�RFA=��=�X]>I ?��+>��=u�>9����H��?�>!�A>xW>��>?-$?�hA�o롽V����9�²s>T~�>��|>���=t.I��h�=�?�>��b><{�.u��A���B��S>o����$b��d��r��=p����=�=�=h,���9���/=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�G�>2�N�e-��V�h��葿�g�0q�>��X?����#¼)	��q�?.��>�$��M��!rҿ�Sk���>b��?���?��U��J��*-���>|a�?�B?T::>Ws�?<]�$qA>� B?��I?��=y?O��%n�
-9?.�?]�?�g>�܋?k_t?���>
ҼĨ������l���U���������������7��k��H����₿i�3��!>	.@=�f�>��û
�(�[==_��������[�>�8>\��>�T�>*�>'��>�0�>=� ���xڏ��L?�!�?İ�B�a�S 0:9�3=�<���f?ê(?�v��������>̉d?��w?��d?��>pM�nK���D��mȳ���g<�o/>�Q?@�?ACK;t{�>�b���_=�l�>���>1�7=gК��I\�= =q��>��?q��>���=�� ?`�#?ҝj>U"�>i^E��9��$�E�3��>|��>�C?�~?��?"ӹ�qY3����X桿�[��+N>j�x?3U?`ɕ>h��� ����SF�sFI����r��?tg?HZ�	?�1�?�??��A?�,f>h}�@ؾ������>d�!?i��A��N&��	��~?�O?,��>k����սB-ּ��݀��!�?�\?�<&?h��)a�	þ��<̈#�l�O��5�;��D���>��>b���pu�=�>&�=�Ym��,6�g�f<z�=_w�>���=�,7�Tg���l7?O�޼�}���	��h�V�(�lb�>G�>Ӷ���?Z,�����ci���1���gཹa�??�?'�?�֬=�n��B?���?���>c�?䑄�L羯��YD���5��w"+��Z�>[?�����W�S��:J��������������>�x�>%ߺ>��>�^�>Vj�>�����F�oLԾ�;�u�x��_���Y���Q����lS���5B�-P�穾^)�����>�ĺ���>���>���=�>�=��>�����;*>YE~=�o�>_��>>,�>���= 8�=)�W=��c��KR?�����'���辻���\3B?�qd?a1�>6i�;��������?���?Ps�?L=v> h��,+�rn?�>�>K��Nq
?�T:=�4��<�<V��>��53����3��>�D׽� :��M�2nf�uj
?�/?����̾�;׽�h���*p=�M�?�(?��)��Q���o��W��S�� ���h�↡���$���p�E珿Ml���-����(�?*=*?��?Jt����(���'k��,?��f>�9�>L��>��>��I>��	���1��]�/'�n�����>�A{?v�>n�J?�,?��d?IX?�C>�<%>i�w�_�#?��f�9 ?<�?G�P?��4?�N?�U?n��>Ƥ>�Zv�zF�޾\i)?�2+?1??�� ?{b?��p���c>[^E=��<���J�<�4=�&�d����&5�|�@<m&��vX?|���8������j>6~7?.y�>w��>Z��|/��e�<�>ݱ
?�8�>Z �Rwr�3b�sG�>F��?��$K=|�)>#�=63���κ�r�=�¼Mѐ=U��l^;��<��=^�=�p�������:	�;���<���>1(?Y@�>�\�<��ʽJf���M&���6��>dy,��q����������`��#>j��?�j�?L�<%�=��=3[����<������"�ݽG�??�U?��)?��i?/&?{�&?Z&>�v��'9�ލ���Gվ��G?b,?΂�>���v�ʾ�먿y3�̜?�T?6Ca�^��(<)���¾�$ս:k>�a/��(~�����D�;�������������?ϼ�?�|@�U�6���"���|K��j|C?���>(P�>�>&�)�/�g��!�GM;>���>qR?p�>��O?g9{?z�[?��T>��8��&���ə�c=.���!>u @?鳁?��?.y?O��>��>7�)����h�����т���V=~Z>���>2<�>��>7��=��ǽP[��g�>�咥=�b>�z�>��>k��>�cw>�G�<��G?E��>�]��3��줾�Ń�X=��u?���?��+?9S=X��=�E��G���I�>To�?���?&4*?�S����=��ּJⶾ^�q��%�>�ڹ>�1�>�Ǔ=
{F=�a>��>���>")�a��q8��RM�]�?�F?��=�ƿ�q�Zr��&��"C���e��򮽥}[���N=;l��~�O���	C�����q�����$���&z�h��>Γ�=�I�=�f�=�x=�.��s�-<��+=�.�;;� =��@�ba<�2W�g׃:�O�����{%�<ɉI=u�7P˾z}?�RI?��+?�C?Jy>c�>�2�H�>O��/b?Q�V>KyL���d;��j��|D��l�ؾgv׾�c�H՟���>C�I��b>�n2>t��=t�<s�=S2t=^��=0H�c�=v��=���=,D�=���=��>.>S&�?��v�߸��8O�O}G��K1?g��>�`>Hd��U\?a[>�p���iƿ6�
��sg?=�@3�?P�,?��;Lx>QfT�P�>�P�=�����X=�r><_��;�>�Ҹ>�>�P��Tp�=���?�@Ƿ8?0���*/ο݀>Z:>Ri>��P���1���\�#*T�mML��?�=���Ǿ��>���=�G㾧kϾ��v<O1>bV=��;�^�}�=�7��;F�=��w=�9�>B�C>be�=����ɦ=���<<9�=�b=>0e<�vD�3H��=8�=C�Z>]�%>2��>
�?ua0?Vd?�7�>7n��ϾqE��hE�>_�=�B�>�˅=gB>���>�7?�D?��K?���>m��="�>X�>_�,�7�m�6l�S˧�޲�<했?�Ά?Ѹ>U�Q<ӉA����e>��+Žeu?�Q1?jk?��><��f�翬	��U����:��F��hd���jM;�������wR�s��=?n�>�B?x��>]s:>�9�=�>�h�>Kdu>����M�v�<�O�<a���U���i���c�����wD�@�����9<Y���a�@g�=�ӻ����]~>ps�>[Ε=�I�>�;�=.�o���U>�B_��K]���^>�H;�I�Bn��݆�&�N��z����z>�7>��7�臊���?jSZ>��	>���?�Wh?�/>C�,�!�ƾ��1��z�	�A��=�9<Lw����U�?`u��J��C����>�p�>��>�:k>��+�PK>��gz=��ᾗ�5���>���@b*�� ��q�<������Y�h��t�W�C?�����=�6~?j�I?�ޏ?��>L���8پ�1>����R== ���_q�����r?�&?)�>G��xD��G̾/���ݷ>r@I���O���ί0�d���ͷ���>f�����оD$3��g�����#�B��Lr���>��O?��?�:b��W��UO�r��#��@q?y|g?��>�J?t@?�$���y�s���t�=2�n?߳�?E=�?b>���=���s?�>�/	?j��?n��?B�s?b�?����>�+�;Z� >n����`�=��>���='�=�l?R�
?��
?c����	������^�"V�<>ء=���>.n�>�r>c��=�bg=�u�=-\>Ԟ>>�>��d>K��>P�>
��2�
���%?���=���>y�2?C<�>&�W=��Ͻ���<��R��T�y�0�0�߽�����<���08:=���b��>�ƿ���?a�W>f��9�?	����T�/.S>�<>�1 ��>�2E>�}>��>� >{�>	��>��(>�¾�q*>$�.�F��gg������r���ܼ>�׵���a�_G
�E||��]�:9ƾ���o4x�����p+�k2�=$o�?"c�=8��������ƾ�/�>L�>+Q?��;Q@=ZM=}J?$l>�i;����������p��Nn?Pn�??�~>���>��K?��>�Ix�F��	Z�'���O��Nr��[m�
��N���g^(�9Xf��-?��r?=sL?2yN�v,W>�j�?����?�E�@.�>��1��a��(:���>����a�H6a���׾�*=�l>?)O?�u�?iJ?Xj&���8q>MiM?��r?}t?�N	?�[8?����g?7#?x�;?��?��:?��T?&�?��>�hM�#�|��Sl���J���{�,����iѽH�`�w�b=�Q��Nu�i=������{�wYQ;$x� �<����=r_�=�}>�1�>�]?>��>HÃ>ΰ7?R(��V9�C絾��+?��=H���^ߏ��%���c����=��h?J��?��\?�)Y>N�>�!�:��>��>:~">x2Y>j��>���H�5�C �=��>��>��=�J;�}������А�e��<x#)>i��>_,|>�����'>z���z�¬d>\�Q�dۺ�-�S��G���1���v�wB�>��K?��?�ə=�W�2���Hf�n0)?�Z<? HM?p�?m%�=��۾��9���J��|�m�>!]�<p������'����:���:�s>�G�������b>vu���ݾAjn���I�k�羾�P=߶�&S=�Y���־U~���==	>)���sF!��򖿦̪�P�I?'�n=|���ʘT��s����>z�>�>�>n$5��*w��8@�܆����=PR�>)�:>v���P��}G��X��R�>��V?ǻh?9�?�����o�&QZ�[vX�5騾=�0?�v>�Z
?�|�<�%�;�\ﾕ�A�v�u���@����>���>B��<H��3����ƾ��&�h�i>q�?�	�>W�:?G��?4��>�a�?u�?�G?3��>��߽+����y.?�3�?���=�(Y���i�����W���?�a?���+��>�z*?�,?��+?�=?_J�>=#�=9��z�D��>�@m>�5q�1ٱ���>��Z?O��>��5?�m?�]p=fd;�d�>��c�="�j>��b>x;#?�h.?q�?�D�>��>������=���>c?�0�?G�o?�w�=��?�82>���>(�=��>���>+?�VO?,�s?��J?��>���<�8���;���As��O����;�}H<�y=���K4t��G����<�%�;�T��I�����h�D�����c�;�_�>��s>
��{�0>��ľ5O����@>@����O���ڊ���:��߷=���>��?X��>Y#���=���>"I�>=���6(?+�?�?E$";ȡb���ھa�K���>�B?H��=��l�p���?�u���g=��m?`�^?(�W��%��!�b?[^?{+��
=�:�þ�b���龕�O?��
?v_G���>��~?��q?~��>��e��(n����uDb��Dk���=�Z�>�w�e�D�>-�7?�s�>��b>��=�o۾;�w�s(��#/?���?��?��?�*>:�n���
�來��+�W?�A�>�W��o�)?�,ɼk���,˙�X����Ⱦ�ľ�%���*������%���肾��J�<�z?�o?|�v?��E?�8�`���e�$1y���b������*9�{�8���B���d����e��Ώ?�E��='E|��xA���?�&?��.�S��>�������4ξk�C>f��?���=�=���-7=�f=Yjh��31�����"�?cº>{�>�t:?�TZ���=��2��n7�V!��>p*>$�>�\�>k��>���g-��>� �Ⱦ��~�A!Ž��v>��b?��J?:o?2��.�/�x��L��K�[��b���c6>���=`��>��f������(��@��xq�����)�����}_�=��0?#~>X��>�v�?�?�M�:���h�|��<2����<�;�>q�h?"<�>�>�<� @#�݇�>ΧO?��>O}�>�9b�b�ﾽӍ�K��<�>�O>�ћ>C2�=Y�7�=x��k������g;�N;>�{`?�v�F����>,.^?�L������:�>�~�%z3����$!�����$S?<�b����>�����*��֎�N���)?%�?����0���r>g$?�k�>em�>�?@�>���+Ո=ߟ?W`?��F?�x0?u%�>>j�;]�w�;z�U�	�u_$=�ǋ>*��>��=��>�O�L�5�j�^�Z<h��=�><%����=�+����<�=vW>��ݿWO�\�
���2�1Q �q*�fD;=N�4>x����"�� �˾TE�:�>���&�H�=�#U���g���H��=o�e��?���?6�TLa=�ͮ����-�8���>2g�-�\�Lz���憽�������ǾW�'�w�P�{�J��r�)�'?�����ǿư��g;ܾ�  ?B ? �y?��F�"���8��� >-C�<�0���뾷����ο������^?���>��^0��p��>���>q�X>cIq>x���螾�-�<��?R�-?���>1�r�9�ɿ]����¤<���?7�@�|A?`�(�'����U=���>��	?��?>�N1��H�>����S�>�;�?���?8�M=�W�E�	�e?�P<B�F�W�ݻ6�=�:�=�==�����J>^V�>���SA��Lܽ��4>�م>�l"����H�^��x�<Ǉ]>��սi-����?�����s��q[��>���<��V?'��>��=�S�?&qx��ҿ��q��>P?��@��?Ǵ2?�繾!�x>�;ܾYJ?3�Z??��>���_��s��<B-�C!�=���]�X�9U>1S?��H<�#��!)���ľF+�oP��nM�=̿��$��%,�tk�<+�����W���Y���Ɯ�5����c�$'����=��>�zS>��>�1h>� �>��]?B�q?�8�>���=�EM����9H��?f>����CNZ������~��i�����XӾ���S��6���Ⱦd'=�
�=�>R�M����� ���b��tF���.?�T$>�ʾv�M�S�-<�iʾ2����󃼰��D7̾��1��)n�-ϟ?��A?������V�4����	����W?�����C㬾�=��4=d�>��=U��O3��sS��?0?�!?�_��ʢ��)>�����<�*?_F?eq<ej�>��'?|�������a>�'>զ�>3��>�T> ����0˽%?)�S?W	ܽ����h�>95žOkp�*�=�\�=�G5�>��8�Z>���<iȍ��
��:���V=�W?���>��)���)5���Y�ެ7=�x?Li?6�>�Hk?:�B?�;�<xf����S����w=��W?�!i?�o>����о����ˉ5?�e?�6O>�h�$��u�.�~R���?��n?�.?���M~}�y����Ko6?f�w?�Z_��M��|�.�^�	C�>i��>T��>h(:�UD�>S�??��"��������D�2�Վ�?�q@�/�?��=�����ga=k��>5$�>y<��8¾jo߽Ѧ��@Ɏ=���>\a��4�|�Y�%������<?�Y�?�1�>/%��������=�ٕ��Z�?4�?���ebg<D��%l�o��:~�<ϫ=��=K"�g���7���ƾ��
�Q������ܥ�>Z@�O��(�>C8�6��SϿ���]оVq���?;��>X�Ƚ������j��Ou��G���H�?����M�>e�>���n���<�{��q;��+����>��
�>i�S�L&������ �5<��>î�>#��>,��$轾%ř?~c��
@οc�������X?2h�?�n�?q?�9<��v��{���a.G?��s?_Z?�l%�1=]���7��j?�_��gU`��4�fHE��U>�"3?C�>S�-���|=�>|��>�f>�#/�{�Ŀ�ٶ�6���Y��?��?�o���>g��?�s+?�i�8���[����*��	,��<A?�2>���"�!�C0=�>Ғ���
?<~0?�{�\.�^�_?.�a�P�p���-���ƽ�ۡ>��0��e\�N������Xe����@y����?O^�?k�?Ƶ�� #�e6%?�>b����8Ǿ��<���>�(�> *N>qH_���u>����:�i	>���?�~�?Rj?���� ����U>�}?�T�>kw�?��=Ų�>k>����1�"���)>>�5���F�>�U?��?g<,>M/ս��.�x4���L��O��?�ن>�a?��N?��>�j����h���,�����d��3�߀J���u�Ƚ��E>M|.>�z>x�0�S��� �?W���!ٿ
ލ����7�?R�>��	?kX�d\���P��wh?Ӱ|>,�⹿M��>����?7�?�?6�������^=���>��>�|�3 �����>oEM?���j~���\g����>G�?C
@��?�lO�׫?{�	�?���!p��} ����w+�>�8A?Z$��h�>!z?�3A>Z�q��J����|��L�>��?�v�?I� ?�yk?e�q��M5���Ͻ��?] �?'ʝ>�O><0x�(�>KK?�4�J[��e
;7�}?!�@�@��H?$o��Ῡ⥿�Ҭ���Ǿ�B>x�>
>+>I�k�/(>�P=��=�ED�_��=Ȍ�>r.�>M�b>�e>�2�>�V�>���	4!��H��2���e=�n���a�z�C�����[{�p���W��/��t� ��.[�����k��C��zrǼ��=��W?_�P?
�j?��?xgG�(�>Q��
~K=-�+��b�=��>�U6?N?),?��p=a��M`b�?~{�L7���x���c�>ΒT>��>9��>�3�>���5�L>`�=>�Ʉ>���=��	=�}b��=�V>�"�>T�>P1�>�A<>��>Cϴ��1����h�w��̽�?����,�J��1��s9������h�=2b.??{>����>пl����2H?E����)�ɶ+���>p�0?�cW?��>#����T��9>����j��]>g- �̀l�ގ)��%Q>@l?�"f>�t>L�3�)s7�u�O�!����({>�5?`���>�7��t��@I��޾{CI>!��>�@�K!�:�������h�1u=;?C'?�_��ί��u�9a��|9R>ĉ[>G�'=�F�=��L>�DW�9��FF�\�2=���=�"]>�"?))>�R�=�b�>Q���UuK���>tC>D)>(�??v.%?�#��Ӝ�惾�n.��*x> 9�>��~>�y>SH��&�=y[�>q�]>����&�����N;@�^Q>&��Ӏb�[r���|=�����=tR�=�� ��}6�+o6=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ��>��Z���(�i�hu���A ��?��B?h����V[�9�?�	�>Q^�yிpdοO�{�:��>sv�?o��?�Nj��O���RD��:�>���?�W?���>Lb��)��%�>@?��2?���>�P��ֽ�/2?�u�?%��?\�K>�A�?غr?W��>X��b�*������2x�!{�V�\�C>
�"=�)��_MX��{��5v���P{�yJ��>�(=w^�>�>�c��''�=T~콩͟�1Ȃ9͍�>C{t>?�l>0��>���>8?�>=��>f��=�Ѳ�� ��ҏ����K?�ˏ?_���o��K�<b7�=�d�c�?3?��0��P;�+�>*^?��? @Z?��>�����e[���贾iL�<'B>˃�>%��>�&i��\>��ؾ*8�M �>9�>�-��D!Ѿ��|�g�o:+n�>7� ?6��>���=�� ?�#?��j>�.�>i_E�S9��8�E�E��>��>\I?��~?��?=ʹ��X3�����塿�[�N>Z�x?�U?�ȕ>����Ń��'F��I����W��?�sg?R�I?�4�?ˇ??�A?s)f>�o���׾������>��!?� ��A�CG&�����{?J?��>�n����ս�ּ���F�����?�\?>:&?��� 3a��þ��<�P#�"�M�E <��C���>�>�+��#��=@�>�*�=�gm��B6��>i<*��=$y�>�1�=�7�j���zD,?�YM�E����=|�r�:kD���>�L>�����^?~>���{����0n��XpT�M�?<��?3W�?!ﴽРh��>=?��?;!?�r�>����޾����w�py�
V��G>���>�Yx��|�Ǒ������4F���Qƽ��h��>��N>��?���>3�K>��>���Cj1���Ͼ���^Ao��%�g�K�oK9�/�����̗������Q��T����>�g����>���>�jw>��>w��>5Ω��/�>!&T=M�R>���> ��>�_$>b�>����H�X��KR?����&�'�0��`����3B?�od?b1�>/
i�����o��s�?톒?(s�?V?v>�~h��++��l?�>�>��q
?�Z:=���l�<+T��K��@��j�Ȧ�>�G׽�:��M��kf�Pj
?^.?���G�̾c3׽y���o=�L�?{�(?��)��Q�ռo�q�W�
S��1��rh�萡���$�K�p�g叿,a���,��ܢ(��)=��*?i�?ir�n�����3'k��?��f>��>� �>�>	�I>6�	�\�1���]��7'�����4*�>�M{?��>�\?�y7?ܕ1?6lJ?�>��v>I�ž��?�9���>�A?5�R?]�8?1s:?(s�>~7?�a>DD�� ��;Ӿ��"?�A#?�{?%�>=�>(%ξ $=�	=@
�=����mF����=qВ��!����ż�#�=0�t>Ub?dT��E8����;�j>>�7?�d�>���>	9�������<W��>�H?D�>�����>r����91�>��?�z	�;= �)>M>�=4:b�j�/����=�׼�t�=ꄛ��@�5D<��=H��=�4�(ݥ�v�;��;�]�<p��>Ã?���>K�=��ԽH>Ӿ�=.��"x>䁀=t']�� �� Ÿ�6P��J���X{�3��>���?���?*��=c��=�<	�vF־�Pa�$�v�����:0?�8(?�lG?��?�:?D�?̑�w-'�+��� ���P���/?Y!,?O��>7���ʾ����3�y�?�[?�<a�����;)�u�¾��Խ��>�[/��/~����?D�(������}��!��?���?3A�f�6��x辙����Z��c�C?^"�>cY�>Q�>��)�<�g�%�@1;>-��><R?0�>
�O?�:{?��[?ltT>I�8�J.��ҙ��n1���!>@?鱁?��?Ry?�r�>x�>ݶ)���VM����������� W=�Z>F��>�*�>�>���=�ȽP��}�>��M�=�b>��>���>x��>/�w>�r�<�G?�=�>+��ر�Kأ�9;���o@��qu?��?�*?�G=_���F��J��P�>�d�?P�?x$+?�T����=�0ؼO����q��#�>�u�>R��>.�=�uQ=�^>�m�>$:�>i[��h�v�8�9+M���?rTF?#�=��ſ=�q�	�p�]���c�d<������d�%c��0J[�8$�=Yh���Z�����5\�^���QN���赾n֜���|����>�V�=��=�=/��<��ɼ���<KCK=�݈<�==�"q�˼m<`�7�~�ֻť���P��7[<X�L=}�Rgɾ�x{?��H?�b.?g�C?t�p>� >I��V�>1!j���?u2e>/
�����5��V��gL���)ھ�վ��a�,5��+M>c,9�U�>��+>[��=��c<!�=�q=[��=�O�{;=��=��=�)�=i��=6�>
"
>���?{�������_��)T�iB1?!��>�i:>��Ͼ�>Z?!<>L���~�¿X���9�v?:� @�b�?�
?)N�<?��>qվL�-��\�̳��(8o=�j��z3�U>?�h�>Q������`����?��@z�\?�?����Ŀ�ƅ�Ό7>.�>��R��1��p[��`�rZ�9� ?2`;���˾/9�>���=+c�zBǾ�"=�6>G_=����\���=_y���B=�im=��>]�C>ֹ=݌��[Y�=TB=I��=~9M>b����:1���'�� 3=�[�=/nc>�K$>ɑ�>��?}b0?POd?a:�>�n��Ͼ�5��i4�>Y��=�2�>���=bTB>$��>��7?7�D?A�K?���>���=��>��>f�,��m�Kb��ȧ�9��<&��?�Ά?�Ǹ>��P<yA���ee>��?Ž�t?IR1?�r?*�>v�����%��G9�Q���[O�;B@=4F}��S ��:��W���n��=���>�l�>jȠ>��|>��T>��l>�3�>O�>/�'���&�a���#��t-�=�X>`����3ü���<�Q�<��n��U��M/)�cn<:���#r�<J�>h �>9ƅ=ݽ>M��=坾��%>�컾�eQ�|^>V&���P?�,�f��􀿹8��f�4��=�U�=8"��o��x�?�_>խv>Ƣ�?%-j?��= a$������o�� ����i�n��<á=W=��.�=��zV�RgQ������>�(�>�6�>P�n>8�+�w�>��o=�C��5�E�>4���q'������q������fi�U����C?�����=�,~?�4I?C��?o�>D��]׾ �/>�n���=�P��m������?Ή&?-��>���`NE��G̾P���ܷ>s?I���O���ٮ0���kͷ�Ɏ�>�����о$3��g��5���o�B��Mr����>��O?��??;b��W���UO�������oq?�|g?$�>3K?%A?+%���z�r��w�=n�n?&��?=�?>/��=���6?�>�-	?Y��?���?�s?y�?���>Ŋ;�� >]����U�=��>J��=�+�=�q?�
?[�
?c����	�������D^�ӣ�<࿡=k��>�n�>7�r>���=ޟg=���=�+\>�מ>��>��d>U�>�L�>�ԍ�ʔ�Ug?_T5>��~>�X9?�v>AS�=KM�F!>B��=</��o˓����p��KҘ=���sսdᄾQ��>G$���&�?̀>[W��?n����p�=��>��'>��.��ٸ>� �>V�e>[��>m�>;��=ɳ�>qX>��۾��>�o'��!��k�����	+��}>�Ɇ�1�f�������A8��3ʾO���w��ቿ_��O�.���?)���df�c��Yc�$��>���>�
?{-m�w�����>�?L:�>����A���o��bg����?���?��>��>IK?G`�>�s��ں�a�S�iDF��m��"h�S�Z�5��쁿���>�����\?�[?�W?>�9��X>��?b�ξ(�!�>�-$��� ��
�='m>���b��������Ⱦ����RN>��S?�+?�|s?#r��AC �`��>N�T?��`?\�?=a?!ո>�V'�}�?0['=��@?�+?�8I?eS?m�>�H�;���=�b&�Q�����T��{��Ȼ��F/ǻ�I0=c=3�:=��I��a�=p� >6�9=����F��u�9=<g��i?��>���=f���	U�>�]?z7?�H>�K:?�/���4�Aގ��V?>�,�d��g{���5��D/��f�=n o?p�?�3z?��;>�2��aG��">h�n>T�->�H>h�>�Q��X��3y-=z:�=L�V>`	y=/�ýo3��y��[臾P)�=�&>�V?b:>����tc=P��~if�5$d>Չ��m߾�\�<h,]�Q*.�`���.��>a�I?��%? /U=m���۬���j�j�J?� ?�bc?=$�?? +>]}���FR��"[��v���b�>���=��������6S���I����@�=�8�������b>vu���ݾAjn���I�k�羾�P=߶�&S=�Y���־U~���==	>)���sF!��򖿦̪�P�I?'�n=|���ʘT��s����>z�>�>�>n$5��*w��8@�܆����=PR�>)�:>v���P��}G��X��R�>��V?ǻh?9�?�����o�&QZ�[vX�5騾=�0?�v>�Z
?�|�<�%�;�\ﾕ�A�v�u���@����>���>B��<H��3����ƾ��&�h�i>q�?�	�>W�:?G��?4��>�a�?u�?�G?3��>��߽+����y.?�3�?���=�(Y���i�����W���?�a?���+��>�z*?�,?��+?�=?_J�>=#�=9��z�D��>�@m>�5q�1ٱ���>��Z?O��>��5?�m?�]p=fd;�d�>��c�="�j>��b>x;#?�h.?q�?�D�>��>������=���>c?�0�?G�o?�w�=��?�82>���>(�=��>���>+?�VO?,�s?��J?��>���<�8���;���As��O����;�}H<�y=���K4t��G����<�%�;�T��I�����h�D�����c�;�_�>��s>
��{�0>��ľ5O����@>@����O���ڊ���:��߷=���>��?X��>Y#���=���>"I�>=���6(?+�?�?E$";ȡb���ھa�K���>�B?H��=��l�p���?�u���g=��m?`�^?(�W��%��!�b?[^?{+��
=�:�þ�b���龕�O?��
?v_G���>��~?��q?~��>��e��(n����uDb��Dk���=�Z�>�w�e�D�>-�7?�s�>��b>��=�o۾;�w�s(��#/?���?��?��?�*>:�n���
�來��+�W?�A�>�W��o�)?�,ɼk���,˙�X����Ⱦ�ľ�%���*������%���肾��J�<�z?�o?|�v?��E?�8�`���e�$1y���b������*9�{�8���B���d����e��Ώ?�E��='E|��xA���?�&?��.�S��>�������4ξk�C>f��?���=�=���-7=�f=Yjh��31�����"�?cº>{�>�t:?�TZ���=��2��n7�V!��>p*>$�>�\�>k��>���g-��>� �Ⱦ��~�A!Ž��v>��b?��J?:o?2��.�/�x��L��K�[��b���c6>���=`��>��f������(��@��xq�����)�����}_�=��0?#~>X��>�v�?�?�M�:���h�|��<2����<�;�>q�h?"<�>�>�<� @#�݇�>ΧO?��>O}�>�9b�b�ﾽӍ�K��<�>�O>�ћ>C2�=Y�7�=x��k������g;�N;>�{`?�v�F����>,.^?�L������:�>�~�%z3����$!�����$S?<�b����>�����*��֎�N���)?%�?����0���r>g$?�k�>em�>�?@�>���+Ո=ߟ?W`?��F?�x0?u%�>>j�;]�w�;z�U�	�u_$=�ǋ>*��>��=��>�O�L�5�j�^�Z<h��=�><%����=�+����<�=vW>��ݿWO�\�
���2�1Q �q*�fD;=N�4>x����"�� �˾TE�:�>���&�H�=�#U���g���H��=o�e��?���?6�TLa=�ͮ����-�8���>2g�-�\�Lz���憽�������ǾW�'�w�P�{�J��r�)�'?�����ǿư��g;ܾ�  ?B ? �y?��F�"���8��� >-C�<�0���뾷����ο������^?���>��^0��p��>���>q�X>cIq>x���螾�-�<��?R�-?���>1�r�9�ɿ]����¤<���?7�@�|A?`�(�'����U=���>��	?��?>�N1��H�>����S�>�;�?���?8�M=�W�E�	�e?�P<B�F�W�ݻ6�=�:�=�==�����J>^V�>���SA��Lܽ��4>�م>�l"����H�^��x�<Ǉ]>��սi-����?�����s��q[��>���<��V?'��>��=�S�?&qx��ҿ��q��>P?��@��?Ǵ2?�繾!�x>�;ܾYJ?3�Z??��>���_��s��<B-�C!�=���]�X�9U>1S?��H<�#��!)���ľF+�oP��nM�=̿��$��%,�tk�<+�����W���Y���Ɯ�5����c�$'����=��>�zS>��>�1h>� �>��]?B�q?�8�>���=�EM����9H��?f>����CNZ������~��i�����XӾ���S��6���Ⱦd'=�
�=�>R�M����� ���b��tF���.?�T$>�ʾv�M�S�-<�iʾ2����󃼰��D7̾��1��)n�-ϟ?��A?������V�4����	����W?�����C㬾�=��4=d�>��=U��O3��sS��?0?�!?�_��ʢ��)>�����<�*?_F?eq<ej�>��'?|�������a>�'>զ�>3��>�T> ����0˽%?)�S?W	ܽ����h�>95žOkp�*�=�\�=�G5�>��8�Z>���<iȍ��
��:���V=�W?���>��)���)5���Y�ެ7=�x?Li?6�>�Hk?:�B?�;�<xf����S����w=��W?�!i?�o>����о����ˉ5?�e?�6O>�h�$��u�.�~R���?��n?�.?���M~}�y����Ko6?f�w?�Z_��M��|�.�^�	C�>i��>T��>h(:�UD�>S�??��"��������D�2�Վ�?�q@�/�?��=�����ga=k��>5$�>y<��8¾jo߽Ѧ��@Ɏ=���>\a��4�|�Y�%������<?�Y�?�1�>/%��������=�ٕ��Z�?4�?���ebg<D��%l�o��:~�<ϫ=��=K"�g���7���ƾ��
�Q������ܥ�>Z@�O��(�>C8�6��SϿ���]оVq���?;��>X�Ƚ������j��Ou��G���H�?����M�>e�>���n���<�{��q;��+����>��
�>i�S�L&������ �5<��>î�>#��>,��$轾%ř?~c��
@οc�������X?2h�?�n�?q?�9<��v��{���a.G?��s?_Z?�l%�1=]���7��j?�_��gU`��4�fHE��U>�"3?C�>S�-���|=�>|��>�f>�#/�{�Ŀ�ٶ�6���Y��?��?�o���>g��?�s+?�i�8���[����*��	,��<A?�2>���"�!�C0=�>Ғ���
?<~0?�{�\.�^�_?.�a�P�p���-���ƽ�ۡ>��0��e\�N������Xe����@y����?O^�?k�?Ƶ�� #�e6%?�>b����8Ǿ��<���>�(�> *N>qH_���u>����:�i	>���?�~�?Rj?���� ����U>�}?�T�>kw�?��=Ų�>k>����1�"���)>>�5���F�>�U?��?g<,>M/ս��.�x4���L��O��?�ن>�a?��N?��>�j����h���,�����d��3�߀J���u�Ƚ��E>M|.>�z>x�0�S��� �?W���!ٿ
ލ����7�?R�>��	?kX�d\���P��wh?Ӱ|>,�⹿M��>����?7�?�?6�������^=���>��>�|�3 �����>oEM?���j~���\g����>G�?C
@��?�lO�׫?{�	�?���!p��} ����w+�>�8A?Z$��h�>!z?�3A>Z�q��J����|��L�>��?�v�?I� ?�yk?e�q��M5���Ͻ��?] �?'ʝ>�O><0x�(�>KK?�4�J[��e
;7�}?!�@�@��H?$o��Ῡ⥿�Ҭ���Ǿ�B>x�>
>+>I�k�/(>�P=��=�ED�_��=Ȍ�>r.�>M�b>�e>�2�>�V�>���	4!��H��2���e=�n���a�z�C�����[{�p���W��/��t� ��.[�����k��C��zrǼ��=��W?_�P?
�j?��?xgG�(�>Q��
~K=-�+��b�=��>�U6?N?),?��p=a��M`b�?~{�L7���x���c�>ΒT>��>9��>�3�>���5�L>`�=>�Ʉ>���=��	=�}b��=�V>�"�>T�>P1�>�A<>��>Cϴ��1����h�w��̽�?����,�J��1��s9������h�=2b.??{>����>пl����2H?E����)�ɶ+���>p�0?�cW?��>#����T��9>����j��]>g- �̀l�ގ)��%Q>@l?�"f>�t>L�3�)s7�u�O�!����({>�5?`���>�7��t��@I��޾{CI>!��>�@�K!�:�������h�1u=;?C'?�_��ί��u�9a��|9R>ĉ[>G�'=�F�=��L>�DW�9��FF�\�2=���=�"]>�"?))>�R�=�b�>Q���UuK���>tC>D)>(�??v.%?�#��Ӝ�惾�n.��*x> 9�>��~>�y>SH��&�=y[�>q�]>����&�����N;@�^Q>&��Ӏb�[r���|=�����=tR�=�� ��}6�+o6=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ��>��Z���(�i�hu���A ��?��B?h����V[�9�?�	�>Q^�yிpdοO�{�:��>sv�?o��?�Nj��O���RD��:�>���?�W?���>Lb��)��%�>@?��2?���>�P��ֽ�/2?�u�?%��?\�K>�A�?غr?W��>X��b�*������2x�!{�V�\�C>
�"=�)��_MX��{��5v���P{�yJ��>�(=w^�>�>�c��''�=T~콩͟�1Ȃ9͍�>C{t>?�l>0��>���>8?�>=��>f��=�Ѳ�� ��ҏ����K?�ˏ?_���o��K�<b7�=�d�c�?3?��0��P;�+�>*^?��? @Z?��>�����e[���贾iL�<'B>˃�>%��>�&i��\>��ؾ*8�M �>9�>�-��D!Ѿ��|�g�o:+n�>7� ?6��>���=�� ?�#?��j>�.�>i_E�S9��8�E�E��>��>\I?��~?��?=ʹ��X3�����塿�[�N>Z�x?�U?�ȕ>����Ń��'F��I����W��?�sg?R�I?�4�?ˇ??�A?s)f>�o���׾������>��!?� ��A�CG&�����{?J?��>�n����ս�ּ���F�����?�\?>:&?��� 3a��þ��<�P#�"�M�E <��C���>�>�+��#��=@�>�*�=�gm��B6��>i<*��=$y�>�1�=�7�j���zD,?�YM�E����=|�r�:kD���>�L>�����^?~>���{����0n��XpT�M�?<��?3W�?!ﴽРh��>=?��?;!?�r�>����޾����w�py�
V��G>���>�Yx��|�Ǒ������4F���Qƽ��h��>��N>��?���>3�K>��>���Cj1���Ͼ���^Ao��%�g�K�oK9�/�����̗������Q��T����>�g����>���>�jw>��>w��>5Ω��/�>!&T=M�R>���> ��>�_$>b�>����H�X��KR?����&�'�0��`����3B?�od?b1�>/
i�����o��s�?톒?(s�?V?v>�~h��++��l?�>�>��q
?�Z:=���l�<+T��K��@��j�Ȧ�>�G׽�:��M��kf�Pj
?^.?���G�̾c3׽y���o=�L�?{�(?��)��Q�ռo�q�W�
S��1��rh�萡���$�K�p�g叿,a���,��ܢ(��)=��*?i�?ir�n�����3'k��?��f>��>� �>�>	�I>6�	�\�1���]��7'�����4*�>�M{?��>�\?�y7?ܕ1?6lJ?�>��v>I�ž��?�9���>�A?5�R?]�8?1s:?(s�>~7?�a>DD�� ��;Ӿ��"?�A#?�{?%�>=�>(%ξ $=�	=@
�=����mF����=qВ��!����ż�#�=0�t>Ub?dT��E8����;�j>>�7?�d�>���>	9�������<W��>�H?D�>�����>r����91�>��?�z	�;= �)>M>�=4:b�j�/����=�׼�t�=ꄛ��@�5D<��=H��=�4�(ݥ�v�;��;�]�<p��>Ã?���>K�=��ԽH>Ӿ�=.��"x>䁀=t']�� �� Ÿ�6P��J���X{�3��>���?���?*��=c��=�<	�vF־�Pa�$�v�����:0?�8(?�lG?��?�:?D�?̑�w-'�+��� ���P���/?Y!,?O��>7���ʾ����3�y�?�[?�<a�����;)�u�¾��Խ��>�[/��/~����?D�(������}��!��?���?3A�f�6��x辙����Z��c�C?^"�>cY�>Q�>��)�<�g�%�@1;>-��><R?0�>
�O?�:{?��[?ltT>I�8�J.��ҙ��n1���!>@?鱁?��?Ry?�r�>x�>ݶ)���VM����������� W=�Z>F��>�*�>�>���=�ȽP��}�>��M�=�b>��>���>x��>/�w>�r�<�G?�=�>+��ر�Kأ�9;���o@��qu?��?�*?�G=_���F��J��P�>�d�?P�?x$+?�T����=�0ؼO����q��#�>�u�>R��>.�=�uQ=�^>�m�>$:�>i[��h�v�8�9+M���?rTF?#�=��ſ=�q�	�p�]���c�d<������d�%c��0J[�8$�=Yh���Z�����5\�^���QN���赾n֜���|����>�V�=��=�=/��<��ɼ���<KCK=�݈<�==�"q�˼m<`�7�~�ֻť���P��7[<X�L=}�Rgɾ�x{?��H?�b.?g�C?t�p>� >I��V�>1!j���?u2e>/
�����5��V��gL���)ھ�վ��a�,5��+M>c,9�U�>��+>[��=��c<!�=�q=[��=�O�{;=��=��=�)�=i��=6�>
"
>���?{�������_��)T�iB1?!��>�i:>��Ͼ�>Z?!<>L���~�¿X���9�v?:� @�b�?�
?)N�<?��>qվL�-��\�̳��(8o=�j��z3�U>?�h�>Q������`����?��@z�\?�?����Ŀ�ƅ�Ό7>.�>��R��1��p[��`�rZ�9� ?2`;���˾/9�>���=+c�zBǾ�"=�6>G_=����\���=_y���B=�im=��>]�C>ֹ=݌��[Y�=TB=I��=~9M>b����:1���'�� 3=�[�=/nc>�K$>ɑ�>��?}b0?POd?a:�>�n��Ͼ�5��i4�>Y��=�2�>���=bTB>$��>��7?7�D?A�K?���>���=��>��>f�,��m�Kb��ȧ�9��<&��?�Ά?�Ǹ>��P<yA���ee>��?Ž�t?IR1?�r?*�>v�����%��G9�Q���[O�;B@=4F}��S ��:��W���n��=���>�l�>jȠ>��|>��T>��l>�3�>O�>/�'���&�a���#��t-�=�X>`����3ü���<�Q�<��n��U��M/)�cn<:���#r�<J�>h �>9ƅ=ݽ>M��=坾��%>�컾�eQ�|^>V&���P?�,�f��􀿹8��f�4��=�U�=8"��o��x�?�_>խv>Ƣ�?%-j?��= a$������o�� ����i�n��<á=W=��.�=��zV�RgQ������>�(�>�6�>P�n>8�+�w�>��o=�C��5�E�>4���q'������q������fi�U����C?�����=�,~?�4I?C��?o�>D��]׾ �/>�n���=�P��m������?Ή&?-��>���`NE��G̾P���ܷ>s?I���O���ٮ0���kͷ�Ɏ�>�����о$3��g��5���o�B��Mr����>��O?��??;b��W���UO�������oq?�|g?$�>3K?%A?+%���z�r��w�=n�n?&��?=�?>/��=���6?�>�-	?Y��?���?�s?y�?���>Ŋ;�� >]����U�=��>J��=�+�=�q?�
?[�
?c����	�������D^�ӣ�<࿡=k��>�n�>7�r>���=ޟg=���=�+\>�מ>��>��d>U�>�L�>�ԍ�ʔ�Ug?_T5>��~>�X9?�v>AS�=KM�F!>B��=</��o˓����p��KҘ=���sսdᄾQ��>G$���&�?̀>[W��?n����p�=��>��'>��.��ٸ>� �>V�e>[��>m�>;��=ɳ�>qX>��۾��>�o'��!��k�����	+��}>�Ɇ�1�f�������A8��3ʾO���w��ቿ_��O�.���?)���df�c��Yc�$��>���>�
?{-m�w�����>�?L:�>����A���o��bg����?���?��>��>IK?G`�>�s��ں�a�S�iDF��m��"h�S�Z�5��쁿���>�����\?�[?�W?>�9��X>��?b�ξ(�!�>�-$��� ��
�='m>���b��������Ⱦ����RN>��S?�+?�|s?#r��AC �`��>N�T?��`?\�?=a?!ո>�V'�}�?0['=��@?�+?�8I?eS?m�>�H�;���=�b&�Q�����T��{��Ȼ��F/ǻ�I0=c=3�:=��I��a�=p� >6�9=����F��u�9=<g��i?��>���=f���	U�>�]?z7?�H>�K:?�/���4�Aގ��V?>�,�d��g{���5��D/��f�=n o?p�?�3z?��;>�2��aG��">h�n>T�->�H>h�>�Q��X��3y-=z:�=L�V>`	y=/�ýo3��y��[臾P)�=�&>�V?b:>����tc=P��~if�5$d>Չ��m߾�\�<h,]�Q*.�`���.��>a�I?��%? /U=m���۬���j�j�J?� ?�bc?=$�?? +>]}���FR��"[��v���b�>���=��������6S���I����@�=�8��qؠ�G[b>����g޾E�n�*J����N�M=���n[V=���־(*���=r
>����E� �i��yԪ��-J?8�j=�t��r^U�k����>龘>n֮>�:��w���@�z���4;�=8��>7	;>N���]��+~G��6���>��Q?&�g?��q?dژ�Yf�|_Z�,�ξڂ���m��H
?�A�>Uo?;O>�X�=t��aU!��Ӌ��0_���>�]�>�.M��e��(�����J��8�>l`$?\�>353?wke?��+? �?߃Q?4"?���>�=���.�.?�&�?\R�;��}�pB:��&l���?̮?��I�Ҕ�>�?�`1?G ?�Y?���>N�=`���Y�Y��>��d>T�~�Gɩ��~�>�@J?�>l�C?�Wq?O?>f�I��}d�;�'=�]>n�9>�.:?��?A�'?�y�>q��>R���q<�=��>c?X)�?c�o?;��=?v$2>T �>ni�=]��>���>�#?�IO?J�s?[�J?�r�>U��<�﬽�<����s���O�D:�;@�F<��y=!Z� Us��f��B�<�պ;������|�,�[D������y�;_\�>t>����L�0>��ľ�0��p�@>�5��0>��s�p]:���=`��>G?K��>FW#����=ˣ�> ?�>��:)(?��??�+;ʣb���ھ��K��)�>�B?"�={�l�����_�u�HBg=�m?��^?xW��(����b?A�]?fJ��=�#ľ'c����O?��
?��G�+�>��~?� r?���>@6e��0n�$���Yb� �k�`B�=�D�>ۥ���d��@�>�7?��>�3c>�=d۾A�w��/��4?���?]��?��?�A*>�un�࿄�������]?)�>>��I="?U����ξ[8����֢�����������;����s%�ߑ����׽�þ=^�?iUs?9
q?6D_?|D �l_c�P�]�� ��f�V�����.��OE�0�D��/C��n��I�d����lQ=��}�tIA�aM�?��'?`�/��>����9!���;:�E>�'��b����=Ҷ����9=�V=�g��F.�������?9��>>��>��<?�#[���=�rS1���7���rP0>|)�>䞓>�K�>��;�4+�e����ɾ`��	ν��u>�Jc?�L?bo?����/�?Z��b �|v9�8�����>> >Ϯ�>�AY�s����'��h?�s����×������=Ҳ1?���>���>ڗ?�?�O	�q��8�z���0�ffr<��>ȋh?!-�> ҄>8<۽�"�l�>�;f?�J?�5�>cT��C~�v��Et�>5s�=B�=9n�=���:�c��V[�ʝ�����? ]���=1�?�O}���M��|�>�u?����H�:Q��>�{����(龺���m��=��?��h<= �>#�^%�����`n)?R.?�����*��d}>d�"?�F�>�2�>t��?���>��þ&��;�>?'_?Z�J?�z??���>&v=����"WϽ��#��S=�L�>�]>�7�=��=�6 �$�X�^�$�H.X=O˶=�=��MȬ�VQ<�����H<��	=�6>��ֿ�sP�K	վ>M��5��n@���/�����%N�<��<�V�������n�&�߽��0=�i���F�U�C���བ��?���?5z׾�'��qK������Gn����>�����;�����dؽ�UھZ���ﾆ]B���U�F�S��i�P�'?�����ǿ򰡿�:ܾ4! ?�A ?8�y?��7�"���8�� >�C�<�,����뾬����οB�����^?���>��/��n��>ू>�X>�Hq>����螾\1�<��?7�-?��>��r�0�ɿb����¤<���?0�@}A?�(���쾍V=E��>H�	?��?>7S1��H����=R�>Q<�?s��?ىM=h�W���	��~e?
P<��F��޻��=/F�=�H=�����J>X�>����QA��Fܽ)�4>�م>�r"�D��v^�z}�<�]>��սw0��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=�h��bȿ.��\	���#޽]E��t���p�h��K���n������=Sw>ش\>@��>Y�r>�'�>��V?�"u?Q;�>7c> H�@ڣ�a���~���@������b�S���������ʾ*��+)�L��H�Ⱦ =���=�7R����1� ��b�v�F���.?�s$>/�ʾ��M�d-<+rʾ����oل����-̾}�1�n�+П?K�A?m���^�V����L�A��C�W?j�ѻ��嬾D��=�걼r=�>�e�=���c3��}S��0?�o?B���`����o)>#8:�<�)?�?�<���>+o&?â�Rѽ��b>�.>���>��>a
>�i��O�ӽ�?�S?,��uM���ѕ>z¾|�u���==��>45��3ȼW�a>3b�<�U���[U�1ń�@N�<�&W?m��>��)���@Z���c�<=�x?X�?�-�>�qk?p�B?i��<�k��1�S���Ew=D�W?�+i?U�> ~��8 о;z��Ļ5?��e?{�N>MPh�_��*�.��R�%?r�n?^?�r��|u}��������q6?��?6r��R��
�@�T~E�|H�>%?��?�A(���?"�2?�cJ�E����W����/����?��@��?5�>�d��\qz=���>M�?L<�{V��������=Ľۍ;?�8��	P����	�]�����%?q�?���>0�ҾpN߾C��=ϕ��V�?`�?����e<k��V
l����Y?�<�f�=7��>g"�����7���ƾ,�
�뮜�]���蟆>X@�B轧�> '8��)⿓JϿ���zо%�q���?V��>Y�Ƚ	����j�
Hu���G���H�L����L�>�>d���������{�(u;������>��M�>7�S��$�������g5<L�>��>��>/��w轾ƙ?�]���@ο����	��k�X?2h�?�n�?Km?sD9<H�v���{�Js��)G?ׄs?Z?Ef%��3]���7�$�j?�_��tU`��4�tHE��U>�"3?�B�>T�-�K�|=�>���>g>�#/�x�Ŀ�ٶ�B���X��?��?�o���>r��?vs+?�i�8���[����*���+��<A?�2>���F�!�B0=�NҒ���
?S~0?&{�i.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>iH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?� �>F��?� �=��>���=2������>�� >�������>��O?�?7�>a�����,�6]C��O���h.C�zn�> h?O?Io>������4%�@�� �Q���<�VH���T�7���x�E><�8>��>`�'�*˾s ?���ؿݷ��ߨD���1?���>�G?����co��R1�w{c?0^�>ē��l��=���	��Ȭ?��?�?mQᾊ������=���>
�>A꽯כ��;����,>|�E?�� ��Q��L�p��Ń>}p�??@���?�Bd�i�"?��0���t���+��&��C�>d
2?�����|e>�>��>���������E�?˦>�J�?*7�?*�?��j?�Յ�&�#��3�3�%?*e�?(?�>]*=�:��f�D>��"?��������̾u\?3@��@y&d?Ij����ӿ�o���g����Ⱦu�>�X>�Q>�$���z=^
Q���U<��<S�+>Z��>�I>��>�>x�>�`>���Ӫ$������H��6@���u>���}L��@%��Ⱦ�"� h���־�3��N�����i��^6��r��"�=�J?�-R?�c?�		?D����=�]�B�>��>�ɞ>�8?VjZ?6B-?h=�E��%ZV��̀������O��a^�>��K>���>�M�>7�>i�27>��D>�X�>��=�x�����`<�C>+�>�X�>��>�f<>�>�˴�.����h��w��̽�?^y����J��+��B ��H��쒟=�f.?�j>~��<<п���@*H?w���T4���+�x>��0?`eW?K{>�����T�,�>;��mtj�3�>�% �3Zl�X�)��JQ>Z}?��f>�&u>��3��`8���P�fv��Z|>�/6?�춾:+9��u��H��^ݾm/M>���>#�C�Ie��������vi�K�{=wy:?Y�?����հ�
�u�
A��nGR>:!\>�[=mq�=8`M>[c���ƽ�H��s.=���=Y�^>�O�>'> �Z=X��>A����Py����>+��>��;=�O?��?'/B�m��i��*|��o>�0�>��r>Z��=�Z'��i�=?�?���>o��:T�ὐ�=�r4$�.'�=�o� "��������>�0���P>Ԋ;���$���A���=�~?���'䈿��e���lD?N+?Z �=O�F<��"�D ���H��G�?q�@m�?��	�ޢV�<�?�@�?)��R��=}�>׫>�ξ�L��?�Ž2Ǣ�ʔ	�&)#�hS�?��?m�/�Wʋ�;l�6>�^%?��Ӿ.��>�Sͽ����'e��4w����S�q�?�@?�����=�>����?@�>Q�
��E����ȿ��Z��t�>��?��?v`�������`�\�>��?�Af?ӄ>�Q�@���D��>�fs?��5?[��<��F��`���*,?��?!�|?�lJ>A�?܂�?p�?�����@Ԫ��Bu���]�M������=\�u<׮��[�K�I{��}����i��6UA��?8>�n
=!��>�⼽TFѾ��=�U�S����{+��,�>l�>k�r>�!�>��>\��>�Ϧ>"$7=��<����$�޾�<N?�R�?0���i��v<wO�=����%�>ZO#?�����K޾�k�>��{?ކz?�`?(�[>�:
������D��v"��y�g=��>�2�>'��>��=��>N�a<��~�>Uih>/�<<�ʅ�N	�����<�	�>�?m��>�Ô>�� ?�#?�j>�&�>_E�9��y�E�{��>q��>1H?��~?��?cԹ��Z3����桿A�[�!?N>��x?�U?Sɕ>S���ʂ���E�=9I�v������?�tg?�\�b?2�?��??�A?�&f>���9	ؾ�����>��!?�����A��K&����}?�R?��>����ґս�CԼ���(�����?n\?�F&?N���!a�P�¾h��<s3%�H�H����;��A��>�m>\��B��=�>RF�=,>m��86�*�f<,��=K{�>�6�=g�6�:F���e;?���+Ծ��ս��y���A�Cu>��=�V��A�?�Ҭ��q��>J���M���ԾS�?���?�?��-��g�6�O?Ʌ?�%?I��>hľ��־.�����A���c�7�?�=J*?y0���!��ͭ��i���ś��-P�����ܗ?�?r>�b�>u��>�_>���>1򩾧 /�Z�����׾�}m�./�O�C���D�8��P�x�_�&�ऱ�V&ľ�#d��?�>�e��X�>Q�?�^1>KM�>���>�	�M�>7E>X�?>�;�>��>�8>��>Fo�=[���^IR??�����'����a����;B?DLd?�	�>>�h�򆅿;����?���?gq�?�v>�sh�%'+�aU?x4�>�,���k
?$�<=k��z��<���7�A��V���p�>�ֽz:�:�L��f��n
?� ?�/���`̾��ֽ�S��QYo=,B�?5)?�)���Q��o�S�W�C*S�*����h�������$�:�p�)����U��m����(��X,=�o*?G&�?nw���ڬ�x�j���>�ZNe>�K�>d��>���>K�I>��	��1�+�]��4'�����{0�>�h{?k��>��S?F�0?#R;?fH?�d�>�U@>O}�Z�?�q�4��>��?+�[?��B?B�H?y��>�[�>a�>*������s�%?V�-?1�?߰�>�-�>(-@�(z>߬�<y(�=��d�o<��RL�<����`��)�<���=�<1Y?���8�����k>��7?Fz�>���>���9.�����<��>�
? I�>�����|r�xb��R�>ڡ�?b�َ=��)>���=6e��vκ�l�=�$¼��=1n���d;�T<��=��=�s�K������:BF�;ࢯ<���>]-?�z�>�>��ؽ�о��'�.H�<Q�F=�TT>�3��!#��[���u��Rv��Sj>M�|?1��?��p>^��=T��=#k��Գ�BZ���q���02�A51?,E?0�.?CB�?G8?��?~.3>m7������^��eN����+?a!,?$��>U���ʾ�񨿔�3���?�[?�<a����;)�'�¾E�Խǰ>�[/�e/~����0D��养�����'��?ۿ�?�A�O�6��x�ɿ���[��>�C?g!�>�X�>z�>*�)�	�g��%��0;>F��>R?��>��N?��z?��[?Y>�78��ܬ�|[�����&�>�@?|��?(��?�vy?r��>��>b'+�ZZ߾�W���������㽂�w6=��S>{j�>��>���>Z �=��ݽ�m����?��y�=>,m>At�>��>+��>6u>�}�<׸G?d1�>�!��\��E���E���y8��#u?�E�?��+?�t=j���IF������>og�?�۫?��)?�xS�Q��=Ցݼ����q��v�> ��>۠�>W�=DH=�|>߯�>ni�>��0��7�eL�*�?.<F?���=Q�ſԺq���p�0����a<�D��@�d�1���S/[���=Fј����E���'�[�a����o������q���+{���>�X�=��=�A�=���<V̼.�<�H=R��<�=�q���i<*�7�3λ�����"���\<��H=��fʾt|?]�I?�+,?�C?wHz>�,>�O�,��>FW��c�?�(W>M�8�����7�Y֧�u�����ؾq ھj(c��`��M�>�1A�2�>Gr0>�m�=��q<�1�=xw=�F�=#*�_=��=�Z�=��=��=T�>��>U8w?ƛ�������6Q�/V�(�:?�;�>���=�ƾ@?|�>>A2�����+c�b*?$��?IW�?�?ji�@c�>���jގ�\��=�k*2>ݶ�=�2�웹>w�J>����M���y���2�?��@��??����s�Ͽ�`/>��6>ǻ>�HW��20���e�kP��@�c�?� <�=m���/�>t�U=J��c�о���;MO>yk�=J��P�V����=sL��KS�=�;�=��>c�=>���=�BS�[��=V�g=O�>�eL>~揻�79��t���G<=���=T�z>1�'>���>y�?�^0?TRd?@C�>I�m�MϾ>O��?�>��=A@�>�օ=�|B>֊�>�7?d�D?
�K?Ʌ�>(։=���>��>%�,�F�m��Q��ӧ�ح�<]��?�І?�ո>5�P<A�A�Š��^>���Ž1s?�L1?9k?�מ>���o$����+�m�������	Q=^-S>�ŽY�y�l>���ǂ=���[�>{�>�7�>��\>��>L��>i�>���=ƌ�<!�>��H�~��2Yڽ?k�<� I=|hL>�/,�A
�Z�1=D����<��G=ң�=��>J�d>��#>'1�>����H�>��7�qȮ��^>�Bʾ0d�.�>�S�{�Y�*�c�ZA����W����X�F>��=�'�>m.,?a'�=��U>�f�?��r?�,Q>����_$���$��3�<�aݽ�J2:be.>�|"��^3���O���,��3��_��>���>
*�>kp>��+�ZW>�;6n=)�6�5�M��>|���Q'����Kq�I���3���i��*���SD?���C�=T�}?S_I?h��?��>�ߔ���پ�	/>d ��Ô=���c�q�S���?hD&?��>]�pE��?̾#羽χ�> TI��1P�1ە��u0�k���Ƿ����>�1���о�$3��a���񏿙�B�Ur����>g�O?\�?�a�uh���VO����������?Ayg?���>�*?�C?�E���v�)����,�=��n?��?b4�?��
>���=�����6�>
*	?���?��?4�s?�?��t�>I��;�� >�͘��4�=q�>/u�=6�=�q?6�
?L�
?�j��m�	������>^�a]�<��=3��>n�>��r>5��=��g=�z�=@0\>מ>�>��d>	�>�O�>������MC?u�=�N~>��*?y��>���=;6�[;�=��'=�+��|���949��
A�ػ�=�q=t��=W�����>8�ȿ��?S>ų��n�>�A	��Z=�3>(%~>u�G�m��>�c�>�]]>�O�>��f>Y- >EI�>�>">Ӿw�>��b��ddb��w�����\m>����D���������;j�0���������q�Kz�{F+���"=�W�?��3�<���^*���x�pR?�Y�>�S8?�ƾN	˽f�'>��?ԧi>�$�+͡�#掿fѾ4��?�Z�?��w>�7�>�F=?b?�|y���.dF�av�dn�2�C��Ac�!���p�p��h$�
GQ���A?ޔb?"�1?�cA>�CS>��?�9��b�k��>���~�L���Ͻ��p>�6��6���-!��F���6��0�;�2a?��b?m 0?�B���μV�> 
G?�J?�Jg?�?�l�>�꾩��?,2ڽgN?��?9]?"�a?�� ?�^�=S���J=�7}���nt��Q�h�Ž�T����W��=�� >�y8=�G�;�a�=L؆��E@�� ��G=��=�3"=f��<!=^�=��>_^?���>�L�>}S8?;f�z�8�E_���*?��?=�w���Ď�Co��`Q��o��=��i?��?�Z?��l>��?���?�_u>Y��>vS)>��Z>;�>
�ݽ�y8�@Ȇ=�>��>ki�=�:�FJ�����g��<�<�A%>\��>�|>~���q)>�ꢾ�{���c>�XQ�X�����R���G��42��w��J�>�K?�3?�ߙ=$����a�e���)?��;?�L?�?O�=�۾z�:��K�B���T�>��<q���e��6Ρ��:�h��:�nt>/��_����a>��ܾn���I���{7=�5���T=����W־�:�����=6�>5���~#!��얿����5I?)�b=�⣾��S������F>%��>,w�>�k$�0����?��	���
�=n0�>B9>���2�F��h���>�aL?F:V?(U�?�D~�~w�(�H�4*��`v�b���Y�?X ^>�F�>!]�;��b>������E�J�����?�@ ?����h�緯��t�z�G����>�p?rZj>�?Yn?�$�>�`S?�P)?@�?��>=����s����9?}�?I� =)o���~��$
��:Y��?6�"?��	�ޮ>l�?�?�??Bf?f{�>�vV=�V%�@I���>�w>, ]�˵��X<p>/l?���>��J?�i?)R>�7G��%*�Ph�=�}�>���=<0?��9?*?�9�>y��>I�����=ƞ�>�c?�0�?�o?��==�?�:2>N��>(��=���>d��>�?QXO?=�s?��J?���>H��<�7���8��Ds���O�vǂ;�uH<��y=���3t��J�0��<~�;�g��5I�������D�P������;�[�>��s>����t�0>W�ľ^A����@>Qۣ�I��ۊ�d�:��޷=���>?���>�g#�*��=���>�I�>���3(?J�?�?��#;ңb�C�ھ��K���>bB?���=��l�D����u��#h=��m?�^?=�W�u%���e?��b?ښ�I8�eɾ��k�w+�h�N?87?�Z>�t��>4x?$Gj?���>�4�q�i�Kޜ�<�o��q�Q��=|4�>��U`x��ю>�wF?���>G��>���=Zk����p���|�.�?\:�?���?Dt�?�	_>�ua�H�޿Wc��^���N
^?y��>����8�?ꆻc ��V݈�CI�����uг�^\���8��i����+��F��	����ډ=��?�/{?#�j?7�R?�xܾd�a���[�!a��I�Y���
�j~�'�;���7��0A��|]��A	��ݾX�s����=�E���>�aw�?�*?�B0�I}�>*�-���Q̾o5>�ɟ��$�'��=hX���7=��=�s�� 2�O����?�7�>.)�>`;?B�W��?���.�K
8�����2>�*�>���>��>�^�������A:˾[��օ˽�uu>�`c?n�K?h4o?A���0�7Y��B$!�6
3�vӨ��hB>?]>���>�IX�>��&�&���>���r�
h�=��[i	�yd~=s�2?�Q�>�m�>c9�?&l?w	��>��ʹx�I@1���<R��>Qi?���>B�>��Խ�!�ʑ�>�L^?�#�>mL�>w�K�8�ܾ�v���J�>�>0��>��=M�(���J�JL|�}َ��|*��3 >�{?��b�g���`�>�1^?�-�6�x��>oY��p��U�������<'?zn=L܈>��羇	6�ˁ�n0оEo6?1#?�C���)J��>��O?�G�>W<�>�@|?&�>�۾�>�f8?Z#r?��D?��?�o�>ӊ��l<`�r��p��>�>F\�>O{�>�ʬ=��0>p����6��F�,x��*g�=�$�=��=F{������J��<�!>L��>5jۿ�?K��پ<���p?
��ֈ������o��	���d�����afx�\��'��V��<c�����A�l���?�;�?ڀ��*/��k���ڑ��V���盽>�q��4��o櫾��$.����ྲǬ��d!���O��i���e�P�'?�����ǿ򰡿�:ܾ4! ?�A ?8�y?��7�"���8�� >gC�<-����뾭����οA�����^?���>��/��o��>ޥ�>�X>�Hq>����螾h1�<��?7�-?��>Ŏr�1�ɿc����¤<���?0�@X}A?��(���쾲�U=���>I�	?��?>�N1��E������L�>�;�?I��?;�M=��W���	��}e?��<��F�-�޻�=pZ�=�t=�����J>�X�>����PA�Dܽ÷4>�օ>�c"�����^��T�<��]>�սP(��*�?p�k��yb��x(���v���=�'[?@��>�
K=�s_?A�V���ɿBST��M?���?���?r�4?,���!��>�)�PW?E?�ɺ>3�v7k��K$>���H ��ü��JV��sP>+�?Ϭ>0�P�Б�|ϝ�aJ���<g�8�ƿ��$�9z��?=G�޺/�[��p�ӱ��-U�!&��qlo�e���h=���=��Q>j�>�W>�*Z>RfW?��k?uN�>z>佬���\ξ9X��L���������(��|裾�R���߾��	�?�������ɾ�6=��=�0R�9����� ���b�[�F�T�.?�^$>
�ʾ5�M�{?1<�TʾS���ԏ�������:̾w�1��#n�K��?��A?B����V�t �rE��
���W?e�����!��9��=kǲ�a�=1��>���=���	3�
eS��j0?�%?ו���M��@h-> $�^��<�*?��?�@<���>��%? ���}˽�]><�.>�9�>���>e>������۽�?�XU?���ʔ�����>���ʍx�X[=l�
>�6�x��6_>��<���9���Fꁽc��<�&W?	��>��)��m\�����:==�x?�?Q&�>�xk?��B?���<�e����S����}w=l�W?�,i?��>z���о�x���5?΢e??�N>oVh�)����.��R��#?Z�n?�_?DN��fw}��������n6?wU�?�u��f��D�� ̈́�Ŭ>?x7?1:�\z�>��/?۽f����D���0��h�?��@�)�?¡=���<{�X=��>�^�>�D̽�߸�~�B����=>�H?~N���d����3�j`<�	�O?�A�?#.
?���� ��M�=b���jR�?4%�?�q��0yg<|��_�k��g��3�<u�=Op�|"������7��#Ǿ��
�򽜾}ľ���>�K@*^��>�Q8�E.�J?Ͽ"
���о:�p���?���>�Ƚø��'�j�/-u���G�(�H�;����O�>�>���������{�Gq;��k��u�>9�8	�>��S��$��:���X�5<��>B��>L��>$A���罾�ę?sa���?οE�������X?Dg�?�n�?+p?>�9<��v���{�9��/G?�s?�Z?�P%��:]���7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�a�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�^�_?*�a�N�p���-���ƽ�ۡ> �0��e\�N�����Xe����@y����?M^�?i�?ϵ�� #�f6%?�>a����8Ǿ��<���>�(�>*N>zH_���u>����:�i	>���?�~�?Oj?���������U>	�}?�W�>6�?�=ݽ�>4��=�D��D�P�8!>H;�=�A�i�?6�M?6e�>���=�5��/�M�E���Q�����C��>ӈb?�`M?�c>&�����#���!���Ƚd�0��oɼ�#A���7���ڽ:�5>]=>EN>��?�:JҾa#?u�3���ٿ�͚��J��R�&?7.�>^u?���	�f����dm?7�f>� �|���_��������?p�?��?U9㾧��9w�<L;�>+��>>���Ϻ�^�d��nt>��J?�D<�)����wb�N2x>#\�?<�@��?�Z�n�?u%�?+���p��{�����I>&??+��;�>EM�>�&>yAv�让�w�o�>�ٯ?t��?o?8�m?�Nh���9��Q�<ּ�>Bpj?A�>a��:��ľ��>Fl
?�s"�����/��&�g?�&@��@DZU?�������=��g���~U��L=K�<<=U>c^��N>�7�=��>��=��A>���>���>Iln>!0�=�B>��)=y�z�21�/n�������o�%�@�����ǜ齳�(��TO��O*�Pq�����H����߽M~K�K��̝���NI��W�=�V?�R?�@o?��?g�e��>�0 �c[+=R�"�1E�=S^�>�3?5O?+?�{�=R�����b����r����AG�>�yP>�L�>E?�>x)�>�Q}��oR>%>>cŃ>w��= v=�0�=`�R>i{�>�>�>�,�>�T<>�>|ʹ�X2����h�N�v�S9̽�?�|����J�V/��{0��g���Yy�=�d.?y{>$���>п@���n0H?{���2*�~�+���>��0?dW?k�>�����T��><��Ōj�v>�3 �/xl���)��0Q>�k?Of>�u>�3��R8���P�9���ߨ|>
6?r���29���u���H�1zݾW�L>xg�>�xF��n�������/ui�a�{=n:?�z?}��������u�kF���R>��[>+B==�M>WYc��ǽ�H��.=���=kd^>L??W',>o��=kL�>WD��K�O�6K�>7�B>��+>i�??;%?��횗�����~�-��!v>���>�>R�>0/J�n�=�N�>>b>���r����*���?���W>�|��_��yu��oy=)������=ܮ�=+j���=��#=�~?���䈿�뾤d���lD?:+?e �=��F<��"�@ ��bH��J�?p�@m�?��	�͢V�(�?�@�?i��#��=4}�>#׫>�ξ�L��?x�Ž)Ǣ�Ĕ	�)#�ZS�?��?��/�Oʋ�3l�W6>_%?ܰӾ���>,���ZH|���A���# ?�Z\?�=�Pw��07���i?'Y�>`d��頿h�˿��s����>$	�?�ԡ?�u��}����P���>���?��l?ib�>}���8hm�;6�>:97?�\)?W�>i�.���ƽ�T#?�'�?��?��<>Z��?��r?��>��j�$�'�.A��������8=v~��s�>��=e����hF�J����ފ��%q�L��gd>pv?=��>����歾ʁ�=!�ܽXn����Pټ>�\�>fB>bl�>�l�>uD�>��>�S=i ս���������ZR?�4�?�@��mw����<�2>C���"�?�>2?a��Ͼ�ھ>A�c?wJ�?|e[?>��>��ꉛ�/۸�戯��_<L�A>�R�>LD�>�����Wk>��ܾ�&/��$p>#QX>�9����$�G�/�r�>d"?�=�>C�>Ԙ ?��#?ӡj>�9�>x\E��:��*�E����>���>�@?P�~?��?�й��[3������塿ǚ[�U�M>Z�x?!Z?kӕ>v������B�F�"�H�}_��̛�?�rg?�:
?�3�?G�??ѩA?@9f>Le��׾�ꭽZ׀>��!?�����A� U&�N�+�?�D?���>i��P�ս0�ּ���e��?�)\?�<&?����/a��þ��<*�"���W��K�;MB�:�>4�>����ו�=
�>Et�=�9m��6���i<f3�=Qy�>�4�=�7�)0��%�,?H���;��T�=|[p���C�JR�>j�S>¾�/g?�W�	{�pL���u��a�8����?J�?Ww�?�U��53k�K�??���?k�?�!�>�K��"վ���;���̀������ >�R�>���`ﾘQ��z������<�ā�)��>yI�>zq?C��>?�>��>���4�4�A�ᾧ��=\�o��G�A�n]C���6�̾Јm��f2�� ����z����>eRL�k�<>�?�>gf_>�>�ʃ��h�>v��=>�,>�u�>��B>�>�&Q=J���m�:�NHR?���%�'�j������NB?#Sd?��>�Fh����?��K�?��?oz�?�_v>#yh�+��Z?�A�>�)���b
?F<=�����<a��m�g쇽2��#��>��ֽ�:�RM��#f�d
?< ?�]��QN̾S׽����r�q=8�?�r)?¨)�s�Q��[o��aW�	�R�u���Th�����$��p����,d��J?����(��q*=1e*?i�?<e��0���8k��?�t�d>��>��>�̾>�J>o�	���1�2]]��&��������>��z?u��>�U?i>?5�&?��O?~�>��]>��Ѿ�5?U�S�-�>z?��^?�`?�3?�#�>�A?�b3>
����	�ɾ��*?�;?��?Y�}>�.?�Ŵ��!=��5�t>[��2 O�?ڒ="�m=b�7�ڡ׽.	7>�e>5c?c��֟8����(k>�7?7/�>���>Cߏ��#����<?2�>�
?���>,����lr��I�#�>���?2��RS==*>�k�=&���Y�ʺ��=/ ż^א=�����w;��<�5�=��=��v�qJ��LX�:���;~�<��>lG?V��>ȿO>TС�	�˾�6+�a6U< ~>�y<O։=� f���$����i�eA�>�"�?��?�V->1�>�_�=Ćj�6�G���r2b�(*;>4)?��?�RG?�.�?er@?�v?�pG>u�6 �������׾�vE?t!,?��>�����ʾ��ŉ3�ԝ?b[?�<a����;)�ѐ¾��Խ�>�[/�f/~����<D�;텻���V��4��?�?1A�U�6��x�ۿ���[��s�C?	"�>Y�>�>M�)�v�g�p%��1;>���>eR?{�>�O?�={?Q�[?�T>��8��-���ә���0���!>�@?Ѱ�?q�?!y?S{�>l�>�)�|ྒྷI������Ղ�ƁW=�Z>Cz�>K'�>��>o�=�ǽD����>���=Wwb>��>u��>/��>ۊw>Ӯ<��G?M��>�]��X���뤾8Ń�&=�ݜu?Û�?q�+?�Q=5���E�~G��KJ�>So�?���?	4*?�S�A��=X�ּ_ⶾ�q��%�>J۹>�1�>�Ǔ=SyF=1b>9�>���>s(��`��q8��QM��?�F?6��=�]��/3s�1&*��<w���u�#w����=�±���G�<�A=2���_Z�zq��qJU���Ⱦ�������y���p%����?Q��=��L>H�=i��=��{�B�_�]=J=]@��ݪ7������c<�k�;~�<!��;�'��wc=Q�=6�=��˾O}?�mI?��+?��C?�y>�C>��9�Jt�>���,�?�^W>sJ�#����;������^����ؾ=k׾sc�p���4�>��E��>"�2>��=J�<&�=�ru=0U�=�_G�/P=i�=1�=��=�t�=&>n|>��?M������l2V�g�5��H*?�>�+�>"x���0\?���=폆�j�5��=�w?�� @@��?-?��Iv�>S*\��4�=j>����R.�=|5�=Vd�#��>��>��)�bp��
�m=���?��@*�>?i���Ɉ˿I��=:�6><>�R�'i1��m\��b��Y�	(!?�\;��4̾���>N�=�^߾��ƾ�(=J6>��`=���x\��_�=�z���;=��k=�n�>OtD>��=鼰��O�=E�E="��=F�N>����7��.�,�2=wa�=,Sb>�s%>��>p�?�a0?PXd?�6�>n�NϾ�?��)I�>��=�E�>Z߅= rB>Ǐ�>�7?9�D?��K?y��>���=/	�>��>�,���m�m往̧����<z��?�Ά?�Ѹ>��Q<��A�Ġ�}g>�..Ž�v?�R1?�k?j�>�U����8Y&���.�'����u4��+=�mr��QU�P���Hm�5�㽮�=�p�>���>��>8Ty>�9>��N>��>��>�6�<yp�=ጻ���<� �����='�����<�vż����ju&�7�+�&�����;���;S�]<���;3��<i��>A�s=���>i�=��Ⱦm��>)���B�c���6>�ž�B�.�3l\�\y��3=��J���>��>�f*�)폿�g?��>I#->�v�?�^?L��=�Ŕ��վ���Iam���P�@%B�!¼�:ľR�N�v�g�}�H�BX�����>wߎ>�>�l>�,� "?���w=,��b5���>|������*��9q��?������^i�~�Ӻ�D?�E��]��=q ~?o�I?���?���>��m�ؾa<0>�I����=Z��*q�s��s�?�'?��>f�'�D��I̾v$���޷>�9I�>�O�������0�@;�Lз�'��>)�����о
#3�f��������B��Hr���>вO?w�?�b��V��TO�q���-���o?"tg?z�>eC?�;?q���v��x��t��=��n?T��?�=�?>���=���>�>A,	?��?���?gxs? v?�t�>@y�;�� >�ؘ�H7�=M�>�x�=W�=Qr?ʒ
?y�
?fc����	��������!^�B��<��=q��>�j�>�r>��=Šg=V��=b/\>[ޞ>gݏ>/�d>��>$R�>�$ھ4�~�?�>>�>�*?�C�>	�S=VtȽ�I<�{���Ҏ��ȋ�v��������<Dz9��z"���+��>Kſ7��?��G>�#�6I?�D�a�">���>C�>���ҫ>}�\>��>9�>f��>2D>�|�>�`>'W�-�*=DQ��n	��a�&F}��1��P�>aM�� ޽���	�<ئ�����i�ܾ�r�N������2ސ;[;�?Ho��}�����'��ǧ�Վ�>U�?�kO?�Z꾮�(��򈽂"?1�3>���~L��0��2�о4��?���?T�=0ߔ>5wF?�>ų�;� ��Y>��t��-6�.6|�+�e��ߋ�A�t����+&�,�G?�z?�O?�ϰ��]�>�D~?���p���-��>�����I�aB�QHj>d{ᾩ?u�yԾ�ƾP����'>վY?�}?2JN?j4� M���>
W^?�&?�M�? M�>I�>���Fv�?��4>b�f?A�"?�O?K�d?���>YV>�-�,�:un(�vI��社.>��p����O�6��Ir>���<Qt=�>�E5>V �<�����gҽ��=,&<᧼p}����>��I?�)�>��G>6�C?��ԽI�J�y�˾C�?{I�J?�������1þ9���:C<�Z?)`�?��l?��>����s0��>4��>��=7"�>�r�>܈A<!�A��Z�=K.K>||>p��=�����Xb���1{����e���>T��>�**>_X���7/>�љ�����0!�>���H�ؾ�J>��oT��:)��m���>��C?�3'?���=9���ҽ�p�$0;?�/?�H?>�z?�Ii=����f�>��^[�7Ɨ�r-�>��=�Q�$��Xa����N����}7>*,���]m�Y'�>#w�C�y���z��v�1J�?�=��V����=��[��5޾
�<l��=�w>�H������iǧ��^?a&��Z���\���*ƾ���=�X�>O�z>^�;։��L��K���� ~�>?�>����rþ@�4�����>�Z.?HAT?��v?پזT�F�=����0�վ��&�>'?V>���>�T>���=7Ă�)��<N`���B�u?���>�B�i�N���c����)��G�>���>�X|>>?��e?���>�yb?P?���>�>�J~=)���0?p?��=������V���I���>C�*?B�潐��>S�*?`]?V�0?�B?8m(?b��=�i���J'���>lŗ>)�f�&񭿌�>2�D?��>�&O?�*�?�&>�k7���v�SO�<3��=J��=J�0?="�> �>��>���>����v�=�j�>Wc?x4�?�o?Za�=n?J32>+��>��=���>���>��?�WO?��s?��J?���>���<�-��,=��Y�s�4oO��1�;ڴH<�ty=x��%t���Z�<!=�;Q�񀀼1��G�C��^��!�;�p�>t>���Y�0>��ľB8��Ln@>�;���D���Ȋ��X:��6�=��>��?^ɔ>��"�D�=s;�>�B�>E���)(?� ?[?=�$;nhb�A�ھqhL����> �A?��=��l�)Q��S�u���g=��m?��^?�CW��l����^?�X?G ߾��1�F���+,��EW�^sJ?�)?��2���>-�?��[?$?Z�E�N^�Lʕ�*�Y��6����=QG�><z��\��>�,?gK�>��:>�ǹ=Nݾ�#|� x��{�#?n�?�ǧ?�ܗ?0cN>��x�a����ԑ�ݍ^?���>�G��z�"?�N�c�Ͼ2���3����ᾥQ��4���J���;���$�낾��ս�#�=��?�br?^+q?9�_?2| ��gc�^�K�� �U�F����E�?=E�C.D�#n�������&��=O=�q�3��@�?��/?+M9�:\�>���@���e#׾�O>�x��0��W�=�>齆�=��=�qV���K�5c���&?cB�>��>N1>?��^�W�5�N�&��d2��5����%>'B�>Nq>���>�����-��+"��ӾԄ�����~-]>�[O?��u?�ڌ?<Τ�����p��1L�ٽyV�*yY=�\�=Q��>mü�g#���Ѿ�(�A��� ��C���*���>ޑ?8�ǽ�m�>"Ϙ?#��>b̾"y�n{�V�g�F�ٽ�>K�0?�t>��=�7[��2�Z��> �l?��>e�>g���P!���{��ʽ��>���>���>�o>e-��\��e�����!%9����=W�h?Ӓ����`�%�>8�Q?X̆:��F<�~�>XKu��!�����'���>�|?�>�=ء;>X`ž^
�5�{��X����D?!�? i��4m���?Y�T?O#W>h�y>���?�v>X�u�w�=S�?��n?���>C�M?bH�>^�������F��e�ֽ�r:�(�=�c>�h=B.�=���g=��:���[=t0;�v����<<�C��5��,�=?=ѼUY�=��Ϳ�v2�'���?�ܾ��ݾ���w
��xy=̾����B�F����1߽�h��! =�@V�2Fƽ��8ӆ�1��?���?w��ɂ������f��(��G�>�|Ⱦp���Gӆ�\o⽺��b'���j��o����p��bn���L���3?x���t��a_����Y!-?�5?Dߎ?A��qM�T]_���=ڈ`<�5��E��-���I̿��=���2?�F�>���G.ϼxV�>�U{>@��=Ɋw�ξ�繾��=��:?��?�k>�٠�����O��B ����?�@IdA?�(�����[= ��>>2	?Q�=>y	3��&�8����>sN�?��?g�J=�iW�_���)Ae?-��;&�F��������= ��=�6=x>��"K>[��>�I��'B���۽�;3>{��>L���d�^��u�<7�\>y)׽dY��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=s6�鉤�{���&V�}��=[��>c�>,������O��I��U��=#A����ǿdc�N� ��D[<�9=Qμ��k���㽞�	=�1M��ӊ�g@��$���K>+W>��>}:�>P�>(e?k��?���>�Y>t�5��zɾu?���>�D������"�\�8�����8�ξ����A� �p>��;�4hӾ�<��=P�Q�����ڬ ��2c�֣F���.?ff>�`ʾ�L�Y�<��Ⱦ4�����H��4�˾��1�C�m���?�0B?�ㅿ�4V��P���������V?���c����c��=�����=�Ŝ>���=qF��O3�_RS�Z7?e�?)վd-��C�q>���|	��E?h:�>��ݼG�>m?�	���C�=�5>1!�>�n>�}�>��=����߳���?f9x?����Ҿ�!�>�w�-�ξ�i�=>��==�r�P���>���������<�"��}�L4W?*��>\�)�e������!�`�:=p�x?��?73�>vdk?zC?���<
�����S�Ǽ
��u=��W?�h?�	>o����Bоe⧾��5?8�e?��N>�+h��龭�.�Tf���?s�n?A?<,���7}�������E6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>��������=Օ��[�?��?�{���$g<J��Ll��e�����<�ʫ=���l�"�����7���ƾ)�
�����Q�����>�W@�l�(�>nG8�2�@SϿz��iQо�8q���?$��>p�Ƚ����G�j��Ru��G�-�H�4������>��=��2�Hʴ��(���BG��;Ǽo��>��+�X�s>��ͽ3T¾
Z�7di>ю�>ײ>��f>5����c���?j�Y���g��Y�޾"�?��?K��?J�^?�R#��B���d�_�1�'�2?�Ĉ?!A?5�۽�:&��~��nl?`ʩ�m`��`?�z�N��>4t?P�>|1�sC=\�o>���>D��:` �Q�Ϳ\ѳ�õ?�梟?'��?6��;
?���?WF??���z���UҾ��:�	h�%�R?yN>����]]� � ���Ӿ`�2?F+?gy9�Χ־�_?��a��p�0�-�CKǽ�ϡ>$j0���[�I�������\e�������x�+��?za�?�	�?���
#�]%?i�>n����8Ǿ!��<Xr�>ek�>��N>�o]��Nv>z��;�Mg	>Ҥ�?h�?+�?-���< ��"�>7�}?�H�>���?�n�=�.�>��=氾��0���">��=Y�=��?�xM?)��>Z�=
0:���.��\F�yR�����C��o�>|�a?\�L?�Rb>(鸽�<0�s� �Wν+2�^��k�@��,�ж�aa5>U�=>mC>wD���Ӿ��?Lp�8�ؿ j��'p'��54?.��>�?����t�����;_?Mz�>�6� ,���%���B�`��?�G�?<�?��׾�R̼�>;�>�I�>I�Խ����]�����7>0�B?W��D��t�o�v�>���?
�@�ծ?hi��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?pQo���i�B>��?"������L��f?�
@u@a�^?*Eɿ����E��a���߷g=kEԼ�>�m��?¤�*s�>������<�8V=ԯ�>��>�/>-�?o�>'�V>��t�t�!�E���Pw�:gK��M&�']��9H�����N߼��ԾB�j���'���J�UZf�!c���z7B�T�=�[?�G?/2y?�?5�A���[>i)����T=�^�.DּN��>�23?Ѥ??�A;?ud/=�����MP�~�z�/�����^�N��>�W�=��>��>�~�>%[@=�Hv>��H>��m>�W>�->��=�v=��T>���>�D�>���>��~>���=!���&��� n�ys8���s=���?��V��~T�"���،��qp��->2`?���=�#����ɿWp��U<?2j��Y�	���I���=ݲQ?u h?d�u>��۽��M��Rk��v���|U��޺Ļ��4�k�	�B��á>��%?�xh>X�u>E�3��8���O������)z>p5?ۀ��1�9�ɯt�<H�BQ޾�lQ>/z�>M���5��򖿑�~�5oj���~=e:?��?�˸�����f[t�g-��ђM>+ ]>�`=׆�=��M>�n�C�ɽ7}H�]�==1=�='W[>`1?��->�N�=�|�>�Q����P�.�>��5>�&>Q@?S�#?�H�A\��	���(�-�-~>F��>�py>?�>��N����=;c�>��l>q&"�<N���w�&�A��S>z���xe��֎�6�~=� ��R��=��=uy���=���!=�~?���(䈿��e���lD?T+?i �=B�F<��"�E ���H��G�?r�@m�?��	��V�?�?�@�?��J��=}�>׫>�ξ�L��?��Ž5Ǣ�ɔ	�-)#�jS�?��?��/�Zʋ�=l�}6>�^%?��ӾWh�>x��Z�������u���#=Q��>�8H?�V���O�V>��v
?�?�^�ᩤ���ȿ<|v����>W�?���?_�m��A���@����>1��?�gY?Foi>�g۾�_Z��>ϻ@?�R?	�>�9�g�'���?�޶?ٯ�?oI>^��?x�s?)t�>�,y��R/�g1��b���#�=�7X;�g�>�D>s����eF�ӓ�c��Ʒj�_����a>��$=#�>�g�\A��T�=�苽�C��`Wf�]��>�q>��I>XO�>� ?y�>���>��=^W���݀�W�����K?��?����n�,y�<{��=�Y_���?�94?ÈY�]^Ͼ1�>>\?�Ȁ?>�Z?�>����2��ƿ��y��욗<�L>Q��>���>u���s4K>gSվ�,E��~�>�r�>px��a�پ�j���㪻�"�>�a!?)3�>�D�=�?�$?��>t��>5���,��e�c�h�>d?�?44�?M:?	�3��(U���w�i��>R�1'�>-��?F�?)�>�f���〿E
�H���bfW��[?[:M?�7��ּ#?gC�?l{-?5�h?Y�>\8	>�d�����,9>�["?��VA�E�&��	�T(	?0�?(��>Y6��ȷԽ��ϼ�����dz?�
[?i�&?��� �`�d7¾N�<2��B
����~;����>4!>�f��*��=��>���=Y�p�K�1��=d<�۵=�;�>8��=��5�:���#=,?ۼG�ۃ���=k�r�/xD���>�HL>0����^?al=���{�}���x���U��?��?4k�?���A�h��$=?�?	?�!�>�J��y}޾(���Pw�J~x��w�B�>���>r�l���S���˙���F���Ž�c�f�?���>�&?�.�>��>���>4��bP��8���`k��<+�k�6����oh�v�����Tʱ��Ҿ�&2���>A���h�>/Q�>w0�>���>B�>[	�͋/>6�N>#˛>D�>e?�>)a�=�>Y>6mk<�V��(LR?P���g�'����2���a3B?�pd?|2�>��h�Ӊ��]���?⅒?�s�?�?v>�|h�g,+��l?�;�>���Bp
?�L:=���P�<V��k��6.����q��>�H׽�:��M��mf�Ij
?�.?�=��ӊ̾h9׽g����;a=&��?�/"?�(���8�]ud��;L�� 8����\�w��z;/�K�z�&���RY��Gp�~H�_R�=�20?m�|?������V��/�Z���Q�gVI>��>�η>���>5�w>ɐ��}<�s�<���0�'F����?J}?{�E>E~O?өO?�DJ?�R?�c�>�R�>�ѾY��>��m���=|5?.�Y?)� ?� .?�?�?�W>�̡���n�1?�D�>���>?��?.r���<��k�=���M%��pϷ�-���y�&�̽�o��G_=\�>ǁ?����8������l>�7?��>���>$���R�����<®�>��
?I��>c �)�q�JS�;��>�m�?&���,=v�)>��=�ʁ��0>��e�=�ȼ�=�=ޡ��d4;�;�<�<�=枕=ׇ������n;��;3]�<:��>Ý?�s�>F�>�������_��m�=	\>ppP>��>=u־Y��(���h�j>,�?>t�?J(�=�O >v��=Q������Z��
C��ٸM<�\?~#?�U?q��?��=?��?�]�=�� �������w7��~Z?�&,?�a�>'����ʾb㨿1`3��?Xv?�	a�vK�O)��¾�ս�~>��/��O~�{��`�C�:M�����3����?Գ�?'8A���6�����5�����C?�z�>;]�>H��>B�)�Ah���C);>X�>�-R?���>l�??��q?W7??_>>��N���5���F��=k.9>�};?7k�?�'�?Z+s?8��>ר�>w��� ������ܵ�����2�����=0`>X��>��>zW�=��
����EM�J
���H�>�M>*�><-?)�>"��=��:���G?���>�\�����դ�K���)]=���u?8��?�+?Qx=�w�"�E��1��E�>o�?��?m,*?@�S�@��=`ּ�嶾�q��4�>��>�0�>���=�G=�U>���>���>B�|\�Gp8��NM���?�F?`��=��ſ
�q��p�g^��v<O<�В��lc�����w[����=�������ͼ��˕[�G �uj���<������kT{�Gm�>0<�=���=n��=͑�<�Jü�3�<�I==��<��=p4m��d<$�:�9Oû�)���9���W<�:N=����˾��}?t;I?��+?>�C?��y><>}�3�.��>㍂�@?�V>k�P�ψ����;�֬��y!��m�ؾ�w׾��c��ɟ��I>�dI�M�>�83>�H�=�Y�<�=-s=�=�R��=�&�=EO�=�f�=���=��>�T>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�8>OA><�R�G�1��\��Cb�Y�Z�?�!?�;��0̾�9�>��=�߾jMƾ�t.=��6>`a=p��@\��#�=�Pz�s�:=^1j=�>}5D>ӕ�=�U���ɷ=�I=�(�=�jO>��N�7�F�,�L�3=���=K�b>"�%>%�>]L?$0?��]?���>��W�	AԾ�j����>n��=��>�=&�.>��>ξ2?[C?l�E?J��>K�x=���>Á�>wR;���o����f&��p���6�?��?�5�> e�<ӎѽ�����1��;���j?�*?��	?�¥>%����
�:��]����<�Υ�sȲ>�!����g�uƓ>��c�U9%����=b4t>���>�R >3�"?b{?K��>a�>���=�r�=�cG<9*�;�=`�l�ن*>>�弳!���>�;ɵ�G<�<
Ҽb��=杢=q�=P�>���k�>K��>;��={X�>.4=�b��.>g���q+C�5�ż��ľ�9�if�� w��=���g�A׶=���>y���01��? }y>j�V>�s�?I�g?Y�h>+J��?���[��iN���ǂ�Kz�<��=�N}�k[E�x<O��;+�_��B��>��> �>�@b>W!0�Q8�WF=Rw־��1�t��>�����۳�t-�i�MW���=��q�l�/J=wuQ?���x�=>ǌ?ŽM?��?}��>�0$������ >W٭��^�X�z�|�5���er?#�?��?xξ��S�/ʾ����׻>k+E��*P��B��!0�`�J����t�>�U���pҾ13�����W�����A�l�p�\0�>�M?7��?��a�ĥ���'O����>���_ ?k)g?Jb�>ǖ?�^?�S��9���~����=�m??��?]��?��>�|o<j�<��?EM?`à?��?�v�?�ח�A�>*T���=����C�<@�o�쩉=��=��?�+ ?�5?�⾽�/��Z����R��7!�=�E�=�s�=��
>�>M��=�!��&����t�<Z��>�)�>k��>���=���>�����߾�'6?D��=�n�>�;!?d�>u
>mSʼ�Q��0���Z�mf1���x�����f�tP;KZ�=�z��t��>�����?��W>���C?g����9��Q>���>�C��)�>�>�+�=\�>���>�O�>�>6KX>�4Ӿ�v>���GO!�C=C��eR��Ѿ�,z>����`=&�����L���SI�g���f��i��)���E=��6�<F�?����d�k���)�����?E9�>+6?wˌ��ш�� >���>���>P#��ℕ������Fᾞ�?���?yb>�ݜ>^q[?�!?g&I��� ���W�8 v�?��ne�/�\�D@�����j���5ɽ�-^?�s?A:?`O�;���>�|?�C)����L&�>��,�ZR;��r=�1�>1s���I��xɾU�ƾ\_
��!H>�yk?Ƙ�?�?`N�H7x��`0>�=;?�J1?��t?*e2?��<?���$y%?�5,>��?�_?+F7?�/?�f?(�/>�V�=R�:p�+=�䚽NЊ�h����6ֽ�輇�M=���=�����~6<;W'=���<�H������_���[���û<5<:=�z�=;��=v��>��\?Ƃ�>�$�>P�6?m<��8�� ����,?VfZ=���Ua���5������>t"l?��?�W?��_>�F�Z�@�
� >���>�>��\>5г>�����H�`��=��>S�
>�ĥ=�rv������d�1E�����<��>ё ?�g�>�ƽ%^>�����g�@�#>�H��p�ž�8&��52��4�����£�>�#%?,F ?�U�=��6%���c���%?��5?<�o?��b?[o=����mUF�b-A�}�/�=>s�ܽ��־&����L���ZC�|P>�}>s̳��Ќ��Ɲ>�%6��*L��t�"���`��*��>�N�4ߚ=mMc�r%龗�Q<��:>��>�1���<�F��|x��Qy?�~�%Yx����b> ��>S��>�׽��g��K�H���%>�]�>>��>���1���3����ᆍ> �=?)�Z?:u?���Ib���H�s����L��@<C�(?1O�>`&�>1�J>�G�=������VW�q7���>�Q�> #�eI�>\P�͞��T�,�I�>o�?v�>>��?ަh?�"?�h?d�+?K?(۰>ۣ��$�˾DF1?�n?��Y=;�0�r�.�1&&�:�C�)�?��4?�l0�1̛>��)?,�	?��6?)*D?�#?��=؎��@���>t��>��j��|��Uռ>~hB?"N�>�bG?�(�?�/5>K<+��	X��Z�Lj9>��]>B�5?c�?��?�>�9�>�y��0��=��>�h?N�?��q?h�=+x�>'�N>;�>�f�=�=�>�>B�?��I?Տt?��K?�h�>��k<+g��w����ӂ�`��5��~�6_=�ռ�^�3u�T#=�^<TBȼ�Dռ���8�C��꒻7��;[��>��s>���->�þ�l���,A>�.ȼ�l��!���X0�/�=(~>��?�u�>��~(�=�>�1�>!K��'?�?�1?(�@��8c� �پ��V��;�>1�@?���=�sm�T����v���U=S�k?�o^?%�[�y����b?Y�]?�T�=�.�þf�b������O?��
?K�G����>��~?�q?d��>��e��n�,	���6b�y k��<�=�v�>5m��d��s�>��7?�2�>r�b>���=t^۾�w� 9��/?��?��?@��?*>H�n��'�u��Ґ�|c?H7�>�`��g|?�e��	>ž2��c�����ê�>���=���l����$��Zq��ˊ����=\&?_b?2ks?�)W?ǉ�h�\�c����4XT��޾�V��r@��6K�H�I�))c�AB��=��A��$}Y=��r�u�A�ࡶ?�G*?X7K��7�>~����H�z�ƾ�)6>�o����%����<����K��b?=}W�M��}n��B�!?T��>��>U�/?OV��4��A;��L�R��$t>��>g��>���>�I����ýyE��fW��bcg>�P?�=V?���?z�y��B�������!�4!u��������=��I>���>ř����w��)ܾܤ��mt�_������	�}�>��5?�_n�#%�>$��?���>۶2�(�W�4�l�z�<��9>�??�u�>R՘<����t��Ʒ�>��l?���>@�>����JZ!���{���ʽ�&�>�ܭ>���>��o>B�,��!\��j��=���(9��y�=T�h?����m�`���>�R?��:^�G<�}�>��v��!����Z�'�1�>/|?V��=e�;>B~ž5$���{��7���EM?�,�>}�����e�oH�>6C?5ߟ>���>J��?��G>��@���>v4�>lT�?�!?�Ed?'�>�E<��V�����fP�G̻���	>v�8>=��=��J>�*X��Ʉ�x�޽i ,>�M����N<.���B�<F⭽3�,�I|4=�]�>�տ@��о��A�޾� �� ��}�-���o���E��;��>�w�q���x�<w�$������V�<��?���?��y���ͽ���� ���+��G�>�Cɾ�w���`�8 D�����}�c���f������_�U/|���Y��f>?�ξ8ɿ뇭��\��5�>`	?�L�?�� �S�E�^f�6G�=�l���ê�l��ܨ�a|ڿ�\R���x?���>�ﾖ�v=y۷>Z�>6�>��>�t�k0���Xv�UG�>e	?�q�>��@<ܿ6οZ��<5��?�@|A?��(�.��^"V=���>Q�	?u�?>�I1�"9��밾L[�>�>�?��?�#N=-�W�Jb	��~e?�<��F��ݻ��=)(�=�s=r��D�J>+c�>���:�A�68ܽ�u4>I��>{�"�٧�ze^����<cg]>�ֽoG��4Մ?�z\��f���/��T���T>��T?8*�>�9�=��,?�6H�2}Ͽү\�&+a?�0�?ئ�?��(?Rۿ��ؚ>��ܾ^�M?MD6?���>�d&�=�t����=�I��Ť�2���&V����=��>��>P�,���K�O��R�����=�����ο��#���&�k���y6i:e�s��&�Ϸ����x�Ӛ���ND���J�t�	�!��=�b>[-�>�Y�>�?>=�`?{,�?�۵>��.>��:�Q�ؾ8��\N>[7��DG���P��-.����\PԾM�̾�˾����L'�⳺��<��~�=_�O�gV���5 �P;i�n�H�`/?�Q�=D¾��C��g�� ežN���V�3>���;��4�'�k�B֠?�lC?P
��`#L�?5��7���Ͻg;V?[��0E�\���i�=W3�;"\�=�Y�>g�=�����.���T�y*;?o�?/a۾~�þE>~h�1�D=��?:Q?
��<�4�>�+?S�%��ʅ=4S�>G��>mu>�ɸ>��>����ݽ0?%Ef?�`z�C�ھ��>����þ6�=�$>�jy���N��f@>�z�<C��ƛ=�������*W?痍>��)�	�W�����G==U�x?��?�(�>�vk?��B?0��<�L����S�G��Bw=��W?i?>�>q���о�����5?��e?�N>z^h�n��M�.��R� #?��n?f_?;��*l}����0��?l6?��v?s^�ws�����W�V�^=�>�[�>���>��9��k�>�>?�#��G�� ���}Y4�"Þ?��@���?Y�;<7 �j��=�;?l\�> �O��>ƾ�z������
�q=�"�>
���~ev����R,�g�8?ݠ�?���>������3*�=f*��N�?���?�x��!�<�W���r��+���XT=>q�=R�<��1��s��s>� �Ⱦr������!��;c�>��@J#�R|�>d�0�u7ֿ"ѿp���>��0i#�/�,?�ܴ>�?6�e��� �M�k�i��TY��R��4J��S�>9��=dYu;��x���y��/$���4����>=��;/�Z>k�%��ĳ�A��X�R=y*|><�>8>cM��ɾ�r�?up㾪jҿs���N���`HA?"_�?'ǁ?�s!?FL�<0f<�5	����k�bD?G�e?�gR?s�#�Os��t=_�t?`��#R\�Q6�0e<��@�<N!?��#?�	�#��=��P>pΦ>�_��_�2��ֿ}ǿ����Ҽ?���?��j �>�E�?١1?M�H0���d��f>����=��Q?���=c���E�,?�*�Q7?)�R?�r���0�^�_?*�a�M�p���-�}�ƽ�ۡ>�0��e\��M�����Xe����@y����?M^�?i�?ֵ�� #�e6%?�>b����8Ǿ��<���>�(�>*N>kH_���u>����:�i	>���?�~�?Pj?���� ����U>
�}?y%�>��?�h�=:`�>�b�=����,�yg#>n!�=�>�š?`�M?K�>~b�=��8��/��ZF��GR�-$�]�C���>"�a?�L?|Fb>�#���2��	!�	�ͽ�c1�pl鼢\@���,�f�߽�%5>��=>�>n�D�EӾ�	?�����ؿAm��͞'��4?���>W@?����u�Շ�?_?�X�>�-��>���K��X�?��?]�?��?ş׾7~Ƽ��>���>0�>�(Խ���� 
���8>��B?�4�p'����o�-�>���?`�@�?��h��	?���P��Ia~����7�v��=��7?�0���z>���>��=�nv�ۻ��^�s����>�B�?�{�?��>�l?��o�<�B���1=)M�>Ŝk?�s?Zo���{�B>��?������L��f?
�
@{u@S�^?)WտRߟ�I*��>���=���=�U>�\½�y/=㶬<��r���t<E>��>��>т>?"�>0~i>�C,>4����%�/j������F��z�����^����z+�����-�� ��<����Qӽ7QŽa?^��t+�)u�~p	=n�^?��V?h�?w��>l��<���>a���X�<�=��h�l��^>,sY?�i ?�=?�[>
���ūn��+��������n�?q6=Jk�>[	?��>w>���>��>�l>��M>��+>�JV>�?>���=�e�>gN�>�1�>ߕ�>[K�=ʣ�����=:w�gǾ�k��ʢ?�0��M�;�3�z��fh������>N�7?)Y�=���xͿ;����3L?m�ƾ�2��&���;�=�t@?Tg?��>]p�1�%����<���Nƾ�k=�J����ʾjN-��>�5?��f>s5u>i�3��T8��P��p���{|>�"6?�㶾�q9��u��H�5^ݾF5M>s��>N{B��e�������+�i���{=�v:?]�?�C��;ڰ�&�u�:���IR>^\>2�=���=�qM>�c�]�ƽ�G�.H.=E��=�^>2d?��+>�Ӎ=H��>c���RP��q�>��A>��+>� @?�-%?��5H���;���-��6w>S=�>}݀>@%>��J��k�=4w�>��b>"�X9��ߋ�u�@�=�V>B���&`�7�x��~w=}0���u�=�=����<�=�"=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ5z�>;���Z��+��T�u�-�#=��>�DH?�X��4�P��=�|r
?[?}]򾟮��g�ȿ��v����>>�?�?��m��5��F�?�B��>f��?�bY?�i>�I۾�+Z�x��>��@?� R?��>'A�I�'��?b�?!��?��I>�/�?�s?���>vz|���.�I>��4��Dr�=$@�;�g�>B>�ľ�JF��;��E눿>k�Rr��e>�&=��>w��N����=+"����h�^�:K�>Xs>��Q>�9�>��?���>���>��(=�����@��(���L?j��?,��<n���<\!�=�r^�?�?4?�4Z��6ϾY��>&�\?1Ҁ?��Z?���>I��(-���ǿ����\�<�K>��>���>"ߊ��DK>�eվ_E��x�><ė>�/���0ھW/�������>�i!?�1�>i�=`�?�X?��>:§>08�������X��<�=�� ?@�?M�?vh?w���9�#҅�8���j���>9m}? �?���>@-��aB�����=������<"j?@��?6�ݼ��??��?+d?�`?x��>#�:�ڕ��Dw���E>E�#?z�
�� A�R�(�B}���	?P�?���>�O��%ؽoӴ�B�����]?݊Z?{�(?��cT_�'r¾|�<9����9�aD�:�Ё��#>�W>@������=I>娳=�xr���2�(�u<�߷=���>}[�=H4���y��<,?�H�l؃��Ϙ=��r��zD�v�>�BL>[���\�^?�s=���{�����~���XU�H��?���?�h�?v���h�-=?��?&?1�>���fk޾N���}w�y�*���>4��>�Hj����{������"G��I�ƽs&��?�.�>F??��>�8N>��>�����N�F�����Nd��'�Wa�9�.���)�[F�s���j�d��㾙�T�x��>��=�\�>���>���>���>��>�{ֽ��%>(Q�>ҥ�>)��>R�V>��m>W�>��<W��MR?O����'���ج��3B?Wod?c/�>��h�X�������~?k��?4t�?�Av>Cxh�x,+��k?!=�>��o
?�G:=%��<��<.^��V��G]��Ki�/��>3׽� :��M��jf�ji
?d,?轍��̾�Q׽&_��lh=��?��*?��*�zTK��[l�+q^��M���{��{`��Ý��}5�a y�mݏ���,'���$"�+.}=�o)?��?lg�Ϋ�����d���I�B}> ��>���>�(�>կ`>e@�z*�kL�AC#�/ޞ����>x�{?>GZ>Z�T?8E?SS?8yN?۲�>�U�>殾�!�>��٬>>��>��J?&�9?x`;?Z?�`)?��2>�&*�C�����Y?x9�>��?��?�+?i":��l
���=UZ��Z폾P�&���<��E��:I��>�=7�4=��e>ӿ?����8��q��t�l>��7?���>g5�>A5��dM��Z��<i��>Ll
?�*�>z���)�q�Ǭ�\N�>���?�WP=^�(>l��=�;��p���R�=mü���=��x�x�2�(�<C�=za�=��\��譺w�!;�r�;W1�<qs�>|�?���>�E�>LB��9� �޵��X�=?
Y>MS>�>�Eپ�~��>%���g��Yy>�v�?�y�?��f=[#�=���=�|��U��u��c���W��<��?'I#?;YT?���?��=?�e#?ܮ>�(��L���_��>��d�?�",?6��>��)�ʾ����3�C�?@]?�;a�%���8)���¾D�ԽO�>^/��1~�����D��u��������G��?ٿ�?�A���6�7u�e���GX����C?R!�>�U�>x�>��)���g�{%�:;>��>�R?�п>�3P?�(_?��<?>_/E�+�¿Cs�����>m�>�<t?��?��?/}?!��>��c>� �;@��_,꾖�3����@�IZ2>}
y>��=a`�>]e�>�Ƅ������ ��&�M�I��>�~�>Nc�>��>H^
?S>��)���G?���>=I�����ꤾ?����u=�=�u?���?q�+?Х=_o���E�����>�>n�?��?k'*?��S��7�=�%ּp���r�uP�>Bй>S�>��=�MG=g>��>���>A�M�}^8��L�P�?�F?ĝ�=�ſ��q��n�%��}�T<H���yd�����Z���=߹�����3���[����^ ������O��{�
�>��=[��=�0�=.S�<[�¼*
�<�O=��<ZH=k���r<��:��wѻ}���x��0mf<9N=����=̾�2}?<I?�I+?tzD?u�z>K@>��9��%�>�Zu� u?'�U>R�L�d�����9�3�������w�־�F־�9c�'͟��9	>��O���>l�1>��=O��<�N�=l�v=���=�κ�=�I�=ł�=\�=��=>��>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=J����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�8>�>f�R���1�X\��bb�X�Z�¢!?h;�S?̾v5�>wѻ=�(߾_>ƾ2�.=7�6>��a=�u��Q\���=rz�OC:=��j=��>G/D>/��=�8��m��=�yI=��=��O>mї�7��+��]4=�M�=��b>�'&>~��>�V?�[7?��^?kÕ>ć<�eɾӹ��C�>���=˝�>a8�<0�K>䙹>�9)?vTF?�CD?L��>�>=���>׭�>�?��tv��i��������׼���?α�?BY�>�\E=�_��Z��>�.�H��??�.*?�I?���>������[���'/�H�0=.��=��=�_ʾ"��#�<tR �2��#(>���=J̭>��c>�2�>�š>�`<>���>� 4>���:{��<���G'�6����:=S��<�0a==w�;�g5=��P]r�j�P=�h�<z���!N<�;>���>7��=��>��ϼ�����H>�z���K:�Yᦽ�7¾4�^�#r��tp�3|7�?͈���n>zU>iyd�?͖�t�?Blu>�{�>��?�wx?�C{>?�̽A���8N����t�M�=��U>�屽�q7�O�-���:���	��>z��>��>�Oc>k�.��`@��<�=�'ھ�A1�?��>�)��VE�`�)��w��[��>A��]_�6��<�F?q���
>fL|?ƇG?_��?���>d��]�羥;>�3����F;�����~��2x���?o�%?:��>(���:I��)̾L����> I�5P�宕�}�0�$G������g�>�᪾��о,3�,Z�������nB��(r�h̺>G�O?��?�*b�'b���cO�����d��0U?�|g?U!�>�F?zG?�~�7^���V�=,�n?���?�=�?M�
>�B���=_�?e��>q��?�O�?X��?�!?���^>~�>�����g/��W�=Is�;yp>?���2�V?��>J2�>݅��������#̾kV���nn���<K�>���=/"�>�O->P���̰����<3F>nm>rD>J��>[ӻ>HY��^��K5?7o�>\5>�?��>V�A>둼�=���｀~��W\=��r��!���T�ż:q�=L*�=d����I�>�Hſ�M�?��	>F�徨f?�g���p�]�E>�>��}���>��= ,=n�i>ɵ�>��=���>�O�=��Ҿg>Z��J|!��AC�b�R�f�Ѿ �z>�᜾�K&�������WI��B���J��i�&6���S=��Y�<�?�?yz���k�t�)��#��L�?m��>`6?����N"��UP>0��>m�>�]��L���6ۍ�u�ᾁ�?��?�;c>͞>��W?<�?/�2��92��LZ�4lu���@�e�͏`�퍿�x��"l
�@Z��z�_?��x?mA?�
�<W�z>���?�&��9�����>��.��);�V�?=`E�>����_�zӾW�þ����E>�uo?>�?`�?�&V�̍>�&TJ>�46?U�&?3|�?�Y:?B�P?� L��]?�>���>i��>�P(?��?L?ö>�3e>?��=��=���������������=�[���˽_����L=(�{=c�=��=�q�U���ֽ��ż�I=�q$>{��=�b�>@�]?�p�>���>j�7?xS�N�8�L®�\5/?rfA=�H�������á����{>|�j?q��?�Z?uwc>�A�HC�F�>��>6�$>6][>���>�`�X�G���=0�>�>1��=��O����	��l��4}�<�>}�?x��>��
���>�ɔ�Ab}�e-`>������ӟ�����9���w����>��:?!?kD�="���E���l�Kg#?��<?N�k?'\?~1�����xK���M�D-a�ޓ�=p���>�%���zx����9��,�==.�=�ؾ#��7-�>c�M���*�h�[�	∿z�5��~�=�s0���<�N��~&���$���1>PI�>���o=�=m���s��^�y?����_����N�_	���>�מ>IK�>d=�����wH��v�i>y��>!>m��=���[�#�(Z�M��>��=?TW^?��?�w���n��.A�8��gP����м��?�z�>�q?h7>��s=c
�����#_��D�/��>� �>�$�FBL�1R��5+��x2%��n�>�O
?�u&>��
?��Z?:?ּe?��*?��?��>@���-���t7?Oc?�����h��p���"�c2<�b�	?�=?0G6��Đ>��?Ps?�5A?��"?|~,?k��=������1����>̥>[�]�VW�����>��^?�̱>�<?�P�?�Y7>�z-��*�����=��V>���=NHP?��?O��>��>"��>������=c�>�Tc?�!�?U�o?���=��?�3>�>lϖ=�{�>��>?O?|�s?��J?#��>}r�<�ޭ�����r��qD�a{`;�e><�Y{={���,Rp���J#�<��;�/���(������3A�B��~�;j�>'�s>���7�0>#�ľ�g��޼@>���C��_����$:��Y�=^]�>��?�~�>�a#�{��=P��>�s�>����,(?��?R'?f�;k�b���ھ٩K�I�>s�A?��=d�l�v����u�16g=��m?��^?�yW�58����b?*�]?�a�0
=���þlc�����O?��
?�G�H�>x�~?��q?o�>!^f�{�m��蜿�b�^Kk����=Ϣ�>z��3e�I�>�7?r0�>� c>E#�=`D۾>�w�����V*?��?=ܯ?��?��)>�n��߿�����䐿��`?^�>Y�����!?�T1;��׾���ӌ�b4�`⪾�,���J���䫾��/�#��䙷�l��=/m?�]i?�~o?��^?ӥ��U�a���d�A݁��P��~��f��/�B�$	J��uI���n�[U��=��n=���Gj=��|�w+A����?'?��3����>sҕ������mξ�B>Y�������v�=TN���=SlA=i�h���(��m���� ?���>S-�>�n<?=WZ���=�oY4�XR9�X���g;>ƀ�>�v�>C��>�J���2��M�˾���[ɽ��u>�.a?�,L?qp?�gV/�����c#���y�9����+?>,t�=���>�a�,�%�+�%��<�Uzt�n��&C���	��K�=�p2?�y>$��>|K�?r�?

�TƲ��:���5����<��>��f?��>=�>���|P#��a�>�N?{��>�=�>发��H�K����f�y��>,�?�A?��>�#��"�������}��A��((>+p�?�b���t��ek�>�_?&��b��=�K�>���d�C�Ƙ����4�$�?H=����=���'���t�h�Ӿ�DC?�?�ȿ��������>kRT?��>T7�>٣?ʪ�>��r�t_K:q�C?���?S��>�c}?j�?&sM��Ķ��{���彎|T=b?D>h�'> ˗=ޘ6>E^����Q��6��j�=�H=��2�d���n�>�gu����=f9{�tx�=$�ҿGm3���Ͼ�C �p��o���Ծ��V��f���I���m��!���匾�C��������� X� M����J5�?D+@@2u��L��ٓ��:䍿%�SE�>�;���Q��X�X��|F]�,���D��[��C�Z��L���XV�c;;?~���¿*x��=&ݾ��?�?��?R��~�(�\d��|�>FH)=vy�<\�y�&O��/ۿ�ݽ��Z?F�>>6���ӭ�i8�>��z>i�l>� �>9���6�1��3�<�i?�?��>E���ſ䝲�����:��?�@��A?��'�L�t4=u��>��	?��;>I�,��i��Ү�ģ�>P��?�? �m=��W���Ӽ��d?cN�;T�E�8���1�=��=��	=d���N>꽓>|(��	@�۽M�2>�!�>�1�{����_���<�_>_�۽����5Մ?�z\�Kf�\�/��T���T>��T?�*�>�:�="�,?�6H��|Ͽ�\�Z+a?�0�?ߦ�?�(?ܿ��ך>��ܾ0�M?XD6?E��>Ve&�,�t����= QἛƤ���㾲&V����=���>܃>�,�����O�tO����=��M�пn�$��\$�w^�<��<=O���#���[ü�!'������v��$����<��>�+�>�M�>��>��F>�zh?]��?ˁ�>܆,>TI/��ƾuj����Ə�����ݔ��� �Y씾q?���߭�"�"����:㹾>T<�z2�=�Q��ڌ����|�f�J��,-?�D>�Yʾ�F�,��;�oǾQ������Fb���k; �1�h�l�Ze�?��C?]f���2P�Ⱥ�f'C����ZUT?��!��������=�*,�D=���>�l�=��ʋ7�,8Q�^??��?r�˾�?;:|�>^��]�=;�:?�f?Ά�vս>4g!?��x�B>(g�>v�>d��>�l>r �=����=����?�q�?���	q��u�>]侂JѾ��w��2>�N��Q��>،>Ga��!y���ɬ�'��?ZW?�X�>L	*��{� ���H�Z�7=�x?�5?Oȟ>xk?7�B?���<0�򾆵S�_�	�ڃt=yW?��h?�)>��|��'о����X6?�f?�O><h�6��T/.�����?�o?w[?�����{�O������?a6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?r�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>�������i�=v����V�?N��?;Ӫ�f�e<�����l��O��|T�<ګ=����1�O8��%8��*Ⱦ��
�@N��h과2�>:@���v~�><�7����9[Ͽ 煿M�ξj�p���?�w�>��ͽ�����j�D�u�ػG�(�H�&o��8�>V,�=��|��܃�*dq�R8��暽���>D�<���>����g���Pà�k�1=2�M>��>;Pm>����ȾE?
�վ�ֿ�����g���=?mю?A�?!.?*�<�օ�圛�����	\?�o?�s?��ji��e��Nl?�i˾xtl��1��XI�@6�=�!?�h�>B��u�>�͗>,A?�B�<I�� V��PT�����I�?���?%�
�l�>l
�?�~C?��(�3���b4����H�	׽��E?t�5>����!c#��5J�K����>�qe?��(����]�_?*�a�O�p���-���ƽ�ۡ> �0��e\�N�����Xe����@y����?M^�?h�?��� #�f6%?�>d����8Ǿ��<���>�(�>*N>FH_���u>����:�i	>���?�~�?Oj?���� ����U>�}?.!�>��?as�=\k�>�[�=W찾{�+��`#>�,�=>�?�y�?��M?�N�><<�=6�8��/�(VF�BR�(���C�D�>��a?�~L?IHb>���Z 2��!�Ekͽ�[1����gK@�2(,���߽�/5>m�=>>�D�]Ӿ��?Kp�7�ؿ�i��"p'��54?%��>�?��r�t�D���;_?Kz�>�6��+���%���B�_��?�G�?;�?��׾�R̼�>8�>�I�>]�Խ����^�����7>1�B?S��D��q�o�x�>���?
�@�ծ?gi��	?���P��Ta~����7�l��=��7?�0�6�z>���>��=�nv�ݻ��Q�s����>�B�?�{�?��> �l?��o�K�B�M�1=6M�>Μk?�s?�Lo���h�B>��?������L��f?
�
@~u@b�^?(�hֿ����^N��O�����=���=ن2>
�ٽ(_�=��7=�8�F=�����=s�>��d>!q>?(O>a;>��)>���P�!�r��[���R�C�������Z�A��Xv�Vz��3�������?���3ýy���Q�2&�%?`���=�Z?�I?�2|?g�>LW��a>���pI=7�u��2��(�p>��E??6?�-0?��=䐊�m�P�a?��3�˾�Yq�"��>�>��>���>[E�>n�μ1W,>�i>�d>u<>�>$S�=�?�=|�>�{�>��>׭�>T�>���=,��1=��G�p�V٧��M*��'�?oM��T�+��2|���ս�TS�r&*=~s=?=�a>r1��NW̿sͪ�zI?� ��DY׾�J����>�H?�c?��>}�m��d���n=������DQ>=н5��H9�dӇ>3�M?3�f>�u>A�3��Z8���P�zy��bw|>(6?0ڶ��W9�Ϭu�ɥH�fݾF�M>Ծ>��?�U\���������i��{=w:?Ж?�⳽	�%�u��o��ZR>L\> �=Q�=H@M>�d�}ǽ�@H���.=Ԍ�=�E^>aR?��+>��=+Σ>UC��d�Q���>�zB>�,>:O@?x�%?���Y��ׂ�I.�R�v>K�>�(�>.5>)�J��~�=7n�>*�b>�Q��C���m�?��(V>�����_�Іw��~=�ϗ�}�=!*�=�t��) =�d�!=�~?���(䈿��e���lD?S+?a �=(�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>׫>�ξ�L��?��Ž6Ǣ�ɔ	�-)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ\h�>�x��Z�������u���#=T��>�8H?�V���O�O>��v
?�?�^�٩����ȿ?|v����>U�?���?e�m��A���@����>1��?�gY?oi>�g۾`Z����>˻@?�R?�>�9���'���?�޶?د�?�J>��?��r?�c�>�}��Vi.����� ����=��;�œ>�
>�Qɾ�nG�$�������j�:p�y�i>��$=M��>ͼ��n���I�=ݑ�e㩾��G�J׶>w�s>T�T>�?�>A� ?g!�>}�>�4=����邾����L?���?�����n�\��<��=�e^�[W?L�4?�V��%ϾZר>�\?4�?�pZ?Ǫ�>�q�%������q���y�<��K>���>I��><���.�K>��Ծ(�C�U2�>i��>�l��r�پˁ�xC���.�>�H!?6��>N&�=� ?��?��u>��P>�+4�k�{��*\��ڐ=�]	?_D?��?�?��6���-��0��XȮ��aT�,�>'�?OC�>���>����w郿�S�=��������̊�?�y/?���=r9?�?\Q?�q?�x�>�_>7�+�͊$��E�>V"?&`�7�A���'���
��	?�t?J��>%���Fӽ{aм���k��G"?�_Z?�y'?���x�`�v¾�>�<����s�R�;���v!>��>�{�����=Xy>ң�=��n�CH0����<ˉ�=�e�>�^�=A)9�	Ӌ��<,?�G�Mۃ���=|�r��xD�_�>�IL>D��e�^?Li=���{�����x���U���?���?9k�?+�ܠh��%=?I�?r
?O$�>�I���w޾ڏ��Mw�a�x�Mz���>L��>�l�5�L�������gE��ƽ����,�>ң ?��9?SCz>wC~>�[?�)Ͼ]"��3�N�!���|��ξr{@�ٶ�-
�պl��4���J?��#�*U�\1�>� ���%w>��?�f�>=�]>R��>b�ؼ�=��=���>|�>�>B�>Ň׼��>�o&�`xR?^5���L(����Ǵ��>�A?,<d?�}�>�qa��c�����w?�%�?�1�?X�u>`\h�,���?��>�O��Z�	?�9=�P��
j<�Q���Q�r����u��H�>!нz�9�M�Âf�ͤ?B�?�Nz��̾��Ͻ�=�� ��N��?`/.?k�1�����C�a}��5���?�c�^��-��5�F'���푿aى��p�}�־/��=Ue2?z-Z?���Pྂ+e���Y��Wg�W�G>4w.?� �>q�0?��>J7�m��A�J�xI1�`U��d�?[{p?�E>�n]?��O?��W?�#H?��>��>�tȾ�d�>5�~|]���>+Hu?�?7�D?jK�>s�+?H�>�͈����-��cQ ?{�>əK?��?���>��r�����E.M>K��4���w�L��=��=�����OR>#�:�� �>�f?"����8���ɩj>m7?&��>�j�>�����o��~��<=�>̦
?�J�>s����nr����9��>z��?1\��	=�)>+��=�_��`�պ���=�ʼ6�=,�|�&69��J<���=P+�=�'��ISF�v��:�֖;�!�<$t�>��?7��>E�>�C���� ���� �=�Y>�S>�>�Cپ����V&��y�g�,<y>t�?�z�?�f=�%�=���=I���W���������B5�<9�?�M#?cUT?���?"�=?�b#?}�>@+��N��@^������?��,?ͪ�>���(�;x���1�4�?Ʈ?�j^������&�+����ս-Z>[#.���}�DŰ�!C@����;��c���k�?D�?WLa��7����cH��Qح�7`E?��>�v�>Y��>2G)���j��~�oB>�D�>v
S?�Z�>�xL?Ҟu?��X?ZfL>?���v��7J�:$zF><J?ʅ?�'�?�x?���>�I>����_վ�1߾��9�����Ft��3�=�TF>��>{��>ú�>ѓ=$<ݽ����9I�h��=�o^>P��>ĵ�>
��>5/l>,�q:B�H?�*�>\,���)����-H}��UF�{ku?mc�?��*?��=ɂ�vfB�U��@�>���?V��?��'?Q����=�ϲ�����8I|�"�>��>���>p�=fSi=�>���>Z��>���jM�	k9�I�/�5M?YC?~��=�ſ��q���p�����d<K��be��ɔ��2[����=l���;���é���[����ɀ���󵾬���;�{���>Q��=JY�=��=7��<*�ɼY��<%K=��<E=��o�gon<x�8��˻�r��fP��kZ<E:I=V����޾.�z?]�??��!?.Z?Lz>,�M>�۞���>o�b=>�>@�:>8�e���ƾ�S�+b���G0��aƾc�����a�IU����0>��n�Ȋ0>T#3>s,h=rt7=.�="��=δ�=��<�I�<j��=�u�= ^�=��B>�:>#�=�6w?X�������4Q��Z罥�:?�8�>f{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��7>v%>\�R�t�1��t\�P�b���Z�4�!?p.;�[@̾�5�>@�=�߾^ƾM/.=��6>M�a=؀��M\���=8Sz�k�:=��j=��>�3D>���=�!��`j�=��I=���=T�O> �"�6�OW,�)�4=���=�b>�.&>ܖ�>]�?�`0?�Rd?>%�>n
n�<Ͼ�/��D�>
�=N�>���=_B>	��>Q�7?�D?G�K?��>1��=��>��>��,��m�J�է��ʫ<X��?�φ?Ѹ>��Q<;A�K��uO>�P�Ľ?�?�M1?�f?�ܞ>�S�U �h�_�+��!<��u>Ox7>�͖��[=�pY93�i�;���2�=Ӛ>$?UC�>`�>6��>�7>|7�>�%>�t����<����$�<�b�a1=�=�lN:8��<�7���}���
��q�����=��S��=+�s�o��=��>��>���>�/˼X�׾T�a>4s�`/<�{�	��1����0�U�Y���y���=�&x���N2>���>���<�1����?6s�>��Q>Ա?6_]?�m�>�W˽�ח�=z����ο��� >��J>�R��9�E}X�3r8�uW����>b A>�!�>ㇲ>i�A�Q�7��0S�i����L���>�������H0��w���Ȏ���C��r#�^IL?����=��='Z�?1�W?i2Q?�� ?��>4��U�R�c���"갾�:_�R>��􌾞O�>��>`��>{W���q���yd�4��>���& P�L���?�+�.� ���/�>�ۑ�,�Q�,�𿅿������B�V<v����>ԸD?��?�:V��~��.U��e����ye�>�l?���>V�?��
?�7< ���`�<�V��=��s?E��?x)�?;>�!����=&�?�h�>.��?O��?��w?��F��2g=납>�~����R��ʁ=���m�>�6�;��\?���><��>�b�3r��ھw���a��*�7=_=Hʩ>�C_>�z�>�=[F�=��=e�>LD�>�I�>R�V>�ΰ>���>ں��&]پR3?]g�=�u�>��.?��>�M<ѽvc.�̻R�r|+���!��Ș���ٽ���D`=�W>O�<���>�Nǿ,k�?�K>�4�Ϫ?"��B/�Dd�=1��>Sn����>�=�L�=뀜>^�>��I>դ>IP>lӾ�\>y��Bi!�j+C��vR�z�Ѿ�{>�����&�ɗ����6*I�4b�� O���i�n4��k;=�[�<�A�?����1�k�G�)�6��N�?�y�>�6?>���腉�֣>���>E��>;.������Lʍ��ᾡ�?d��?�Ac>��>�W?�?5�1��3��rZ���u��&A�Oe�	�`�<㍿������
��3��?�_?��x?vA?� �<�Kz>렀?��%��ݏ��/�>`!/��';��<==7�>�!����`�'�Ӿd�þ�� NF>��o?!#�?BZ?OV�V�����:>�.7?{5-?F�z?�b0?d5=?����?��V>�	�>R@?� 1?��'?�?�'>��>���O�N=�_��i����qϽ����i �@�<�/=e^<`�
=F~w=�7=��¼�^�5A����;�8�;0�=+��=#�=L��>��]?�>$��>��8?
���6�Ō��-N.?f�L=�⃾7���ѯ��x#񾮢>��i?��?�=Y?wd>�C�	�C��>0ǉ>��'>=Z>z�>E����C�y�=��>M>��=J�Q�J���t	�&Ï����<��>�w	?ع�>zv�3�x>ɽ�������>qF���w������K�!��#��X�����>�c??W?Ҩ.>
�2�����y�g ?Q�,?*�k?�a8?1�q=m璾^�7��w)�����ڜU=Ha�W�Ⱦ6ޯ�nJ��V�K�!��b��>ɾIî�^�>,XC�kލ�A������
7�Ґ> �j���<=��׾b��.G<�=뇮>��b�mf/��!��Ӧ��O?�>4|��!����c=j΂>B�_=�k�<�J�f����*��Ŏ>�و>��>�=b=��v^'�U�|�>R�5?�`?���?Fr��Ec��=�I���Myľ8�q���?��N>D��>��0>߷=Tm�����f*a���C�$M�>���>|&��H�ѝb�: �������>�?���>�H!?�s?Yg?V�f?��7?�f?�Sz>\(?=�CN���.?A�y?`�C="���(�?�=�1��D?����>��)?��ѽ��>��$?��?o4?}F?�B?�e�=�u꾙�"�8��>>@�>nr��d��x�+>l�A?\��>k-9?���?rR>�;���Q�&r �3>V>{�.?��?w+?�#�>�ƕ>����s�e>�`>���?ȭ�?�l?N'Z>�� ?�Mg>\�>Ry>z�>3�>��#?�Q?f��?��;?L�>��p;��ϽT�ܽf�<�y�����8�޺n��=G3=��
��Fd<�i�<���<�$\<�y���c
=BA�M�V<��<&W�>tWr>L��$�">"q¾qX��̇>>�q��{�������3,����=apv>p�	?��>��K�=Jr�>���><�r�'?h_?T�??;�Ja��оc�N��h�>[X<?��=Jn��e��n�o�̏H=2p?��Z?]Z���
c?��]?�����<�*pþM+b�a�龀�N??k�D��ϳ>�>?�;q?��>�e�Vm��ǜ��&b�[)h����=�y�>��He��Ü>e�7?���>nQ\>���=��ھMax�n����?N~�?�,�?�a�?D�)>�uo��߿K���K���8b?���>�o��� ?���#Ͼ�Ò�=c���d�C6���#��Ex��J����9�葃�E^���$�=a�?I)i?Sp?jK\?>O�z�[�60h�2-����O��m��0(�G�A��/Q��
G�5j^�z�=.��֝�	�=��p���C�`��?�$?iA���>�<��� �t�ԾX]>`V���%�z�<�ٽ>J<�;<�j�i!��㪾�f#?eϪ>�	�>;k8?j�]�x�4��DF�B�@��2꾽=V>��>�W�> �>�JU�%\ýZ�ܑ�좈��J���|>�Z?�NK?�o?��-��!�*�~�+�|��W�����E>W�3=�x>܅�UW*�
��nv0�l�p�F0����Xv��U>�8?�=Q>O��>��?���>q�u��'��xM��7p;C��>��D?4d�>��>Se��[1����>��i?ۆ�>�c�>&�����#�SM��ö�����>p��>�?�}>�-���Q�|B��������7��$>Ǟd?a���O]g�w��>��R?QvD�j�=뱪>j<��V)�[���y�g��X=}�
?&ł<��>�̾������_����??��?�
����D�8|4>�I(?�o>��	�dʟ?��>��̾�Bc><U?f I?i�?��?��>,6s�m.=����BJ��ܤ=Y6>�>��	��p�=Q�߽tT��)�9�w"8>{*�=����"->/���3:=�Z�=�>V׿h1G���&���6Ҿ��{龯�>�Oc��\0��\���ۖ��2����8���>%P,�ɧ���l��1���E(�?O��?˰m���Z��������<,�L�u>�����ͽ~؟�O`����������t���_�=�G�#�g��(T���9?X�پ�"ÿ�.��.[���+?��?8km?�F��S=�8��L+�=�[>�0�_��$֤�OοZA�P�}?º�>j	�%/�<׎�>�4�>G�J>���>2ٴ�bL@�8h�)��>Z?��>�����οb���/��=�U�?X
�? �H?6�վ��u���>a(?;W>o�p����KE��5��>-�?"�?e
>��N��B<$�N?��0�.�F��>ֽм!��7�5?�>C-z>�H��!��W�ٽ�L=�>W>E#�B&7�[8���B�*�}>&n�NH̽5Մ?'{\��f���/��T���T>��T?�*�>H:�=��,?R7H�[}Ͽ�\��*a?�0�?���? �(?@ۿ��ؚ>��ܾ��M?dD6?���>�d&��t����=�6ἠ���~���&V�G��=Q��>m�>ɂ,�Ջ���O�J����=�~�K�ڿ�^(���%���_=	��O���s>Z��Xa<�{��C���p2���J>G\�>��~>:M>�˂>�y>#i?��{?�|>��!>u&��Ǭ���D)�Q����e��
 ��� �㺽�-���弾�!��i��iED��w��S���<�d�=�?R������ �R&c�*�G���.?��>�ɾ��L��G<�Jɾ�慨��N��w����̾Պ1���m���?�B?b�q�T��!��M
�K����T?k
�@��.�����=M�-J=�S�>��=�K⾆53��R��6?�?7ȾӃ���
>�z���j��"?�+?���>I� ?/�]?�ꑾ���>�^�>+X�>���=�b�>wus>�'����ѽM]?�gL?�T�~Ǿ�>�a������p���#�=�؟�I�@=᫐>��=�w�F��<C%�>	)��[?h:�><%�b��v)��ҵ̽v���h?�s?|��>�Au?eqY?A�����39���Ҿ}o��G?�:i?6D>
>-��3�3�ɾ�/?��^?d>潾I�ξ����9!�2� ?��e?ן?䮣�x8k��$����"��� ?��v?{s^�p�������V��0�>�]�>��>��9�Yp�>	�>?�#�G�� ���*`4���?\�@��?p)=<�`��ǎ=�;?�]�>�O��6ƾz��&����Kq=n�>�����av�7���Z,��8?.��?F��>����p��	Y�=
����?z9�?�z��
\�<�����k�������P<��=&	$�Wy��A,���6���;8��Х���¼\�>�@�P�0^�>�a7��߿:�пk�����ƾ"b�3�?ը>�x����}�d��s���K���F�]̇����>��>����"����ku���8���7��>:�����>�40��®�Eɠ����<=ƍ>�=�>".�>hQ�����Fv�?����Ͽ>���A��R?�T�?%8�?��#?�=��p��jD��hf;!�G?�r?�Z?�8`���L�@�L�<�s?�����;�B|-�[=�:�=WX6?B??�Ծ�@��y�>?�>�>l
�	⿊�ÿ���1 �?�$�?oݾ9��>pΝ?^�S?�4��3�����z����&N?��>Ia���e������_�Gt9?�(i?x�r�հ(�]�_?*�a�N�p���-���ƽ�ۡ>�0��e\�	N�����Xe����@y����?M^�?i�?ֵ�� #�g6%?�>c����8Ǿ��<���>�(�>*N>|H_���u>����:�	i	>���?�~�?Pj?���� ����U>	�}?3+�>��?�H�=�U�>�V�=���TR-��Q#>�!�=��>�.�?��M?�D�>��=��8�P/��XF��HR�"���C���>\�a?_�L?�Gb>����1��!���ͽQm1�C�鼟h@�:�,���߽,5>�=>�>��D�?Ӿ��?
x�q�ؿ:k��Rp'�Q44?Tă>/?h����t����36_?��>3�b/���,���d����?�I�?�?��׾9eʼPG>��>�-�>y�Խ�̟�����d�7>��B?*"�rE���o���>���?͵@Xخ?;�h�[	?m ��O���_~�0��B7����=Y�7?-�w�z>���>s�=�nv�l�����s�c��>�A�?�{�?���>��l?�~o�o�B�&�1=�I�>%�k?�r?��q��󾆮B>Z�?�������/L�5!f?��
@u@��^?.{+�ˠ��%צ��پ�x�=���=��>��=�;>�}=ռTď�/�O=���>q��>@��>֬�>��>F>�4��� &�?���'��E�d��*�CGݾH�����L�a��]��iʾLݾ�%y��C�WC��q=i�����L��O�a=�{?!�Q?iK�?.��>�<=ߓ�>ʽ�,�=�J���o�6>P�G?Z5?��*?t��>R���i�5,���ʾ�QF��
�>ׂ�=?m�>yc�>��=Nܿ=��>_�>�w�>S�u=&T)>Y��>
�d���>x��>���>ܙ>>U�>�贿E֯�Oi�Ԛ}��Hݽ���?Dݞ�״I������;�������[�=9�-?�J>wґ�ьϿ:8��v*H?�������<4��D>��1?�W?S] >�-��J�V�C�>i����l����=�'��ds�[G*�ҳP>�*?�bg>��u>�3��&8��P�ʨ��u�z> t5?����q8��~u�{H���ܾ�M>�u�>_6�1O����y�~�Z�h�e�}=�	:???z���j��gVu�G���"�R>5w[>%�=�Ъ=��M>F!h��lȽ�RH���2=ʐ�=+�]>�?G�1>_�x=��>���Q"h��?�>B{E>9>��C?�*?_y��Fζ��`�Ƶ(�U�z>N��>�ф>��>�I���=��>9�b>�)�l�d����R�I�=>^Ԋ���m��Ɲ��k�=�*��V��=$j�=�ҽ�Q�7��<�~?���(䈿��e���lD?P+?A �=��F<��"�D ���H��E�?q�@m�?��	�ߢV�;�?�@�?��U��=}�>׫>�ξ�L��?�Ž1Ǣ�Ȕ	�@)#�gS�?��?��/�Zʋ�>l��6>�^%?��Ӿz��>���L��� �����x��ZJ=��>��D?��L���3���?��?3������D
ǿ�7{�<i�>�
�?.�?�;k����]�H�'u�>��?{Ca?�6k>x�Ⱦhkl��{�>�9?L?�ַ>K-���4��+	?h��?-��?�I>M��?7�s?�d�>�Gx��X/��5��T���T�=�xb;�v�>�q> ����aF�Xԓ��e��ۼj������a>ޞ$=�>�|佪2���S�=�#���G��Nif�M��>�<q> �I>�\�>�� ?�j�>�>��=Kt���܀�L����L?aێ?;�:gn���<��=��`���>��4?)'�l�ξ�=�>+�Z?p%�?��X?��>X���`��4ý�#ǳ�/9�<(XM>&��>&��>+����K>��վWD��H�>�|�>��żm[ؾ񮀾�D���>�� ?l	�>%��=3`? �?�:�>��|>9~"���q�r�Y����>�
?�%?`�?m�'?g�<��k	�'o�ő���g���>%�h?!�?��>m����G��/>��ܢA<�֌?k?|p{>$8?�/�?9�Q?�v?��>��u>��־LY�=���>�:$?�*���D��B(�����K?�� ?�`�>g�W��Ȯ��&��� )��#�?ܪT?Bl$?ú�%6d�������<0�<�x5`��O��w�g�(>�r>��E��=sd>���=�On��0'���9���=5\�>�<�=�kE�mm���@,?/�_�~��x�=s��TD�,z�>�M>=���W^?�G<��m{��묿�T���X��s�?e5�?A��?J����h���=?��?}�?�A�>����ݾ��:z�Ҟ}��"�?�>��>/�i�!8⾺_��� ��rI��Z_ʽ�u۽��>���>E,?"��>��>���>5�˾:��P��]�_v���\
��m*�xLD�4����^���&�ؒ8���þ��{�X�>jƼ<�m�>}P�>��b>R��>ݜ>r׼��OW>7�Y>r��>Wj>�>�]a>x��=Uo=�Ž�R?����H(��v��t��*^A?j�b?ѐ�>�OF�����%���j ?	�?b�?�v>,4g�AN*���?}_�>���T	? �H=&9軘֊<�M���j�g�{���5����>��ͽGl9���M���]��?? 3����ʾ��ܽ\�_�>7�/��?u,?��(���,��[n��X�hrJ�����-9��y˾X�X�6�}�@`���[���|�/���;�5.?Ֆ�?��QC�(�[���W�N4_��wi>�%?]��>5@?��>�	)��4�J�+�q����Ͼ��>5}z?g3>>^[W?PcK?�W[?8�W?�ӽ>i��>>���ʻ>���<R�:>3��>W�1?�_*?YB?O�	?{N9?�'>������w?OQ�>��:?�?�?E:D��U��=�i�5��4�T���<]��{�P�i����">�R�>��?�q�� 9�������i>��7?���> U�>n��������<��>��
?�Q�>p �1�q�������>�z�?p�W =��)>�i�=��q�Uͷ���=�Ǽ�v�=d����4�)u$<�?�=��=&��Y�Ji;c��;�ܰ<�t�>��?@��>�C�>�@���� ����$d�=]Y>�S>>�Eپ(~���$��K�g�-\y>ww�?�z�?�f=��=_��=v}���U��W��B���u��<�?mJ#?>XT?{��?{�=?�i#?�>�*�*M���^��{��ڮ?Z!,?{��>���&�ʾ�憎f�3�/�?�Y?J9a�ˤ�'3)��¾Bս~�>iX/��*~�n��D�t��l��2���X��?D��?�WA��6��q辭���e����C?��>H�>��>&�)�P�g�z$�JG;>Wz�>oR?:f�>d�O?�Dz?��Z?��S>�9�-��嘿9����'>[�A?��?%
�?��y?��>s�>0C-��Nݾ ����^�{��)'��k\=��W>�ڒ>P.�>ɧ>_@�=8�ɽ%���9�B�f�=Zb_>i�>n�>�X�>nqr>B&�<��G?2��>�n����:餾�����{=�t�u?��?��+?j<=ik���E����7�>�j�?8�?f *?�S�:��=�ּ:���<�q��>f�>�!�>��=��F=X>���>Ə�>�2a��r8���M��?0�E?x��=�iĿ��m�R {�#b���qr9 U���yw����:)~��	�=���u���S��� a�ۃ���.���n���;������� ?L/�=j�=T��=�n)<���es=��=�x*<4� =W�y�EL<���ث�������$]�;��,=�lл{�;�t~?�6K?�1/?:M?�z�>�H>h�|��#�>L���"?��=>��?��^ƾ�:��������վT˾�j�!˛�cl�=T�j��">�>���=�*�;�	>4��=E�=��<�/Y=|�=���=�q�=/#�=�_>��>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>R�2>��5>>2e�������+���D��vr?� @� �Ⱦ�<�>�3>�����̾�2�=�+M>j�[<D6H�$�o�-�=Rrq���u===%�>��X>c�=.�w����=��=A�>��[>�;T;Խ�'��(�<��=x�Y>�J>)�>�?��/?�c?ჸ>:�o�t(ϾP���^�>6v�=��>�%�=�7>v`�>I�4?ԂC?�I?D$�>Ӓ=�ݿ>�U�>k2�o�R�߾W���ߧ<$��?�R�?(<�>��<=��(��)6� ���w8?��*?aF?}t�>e��g�d�#�8~0�����ċ]�7ӵ=�)��м����` ����8֛=���>Y��>�ί>ׅ�>�6a>��I>6и>e:�=����z2�=��Ż	��l��/��=>�2�i�==�퓻%�r��m��)�R`�<&뼲򽖝�����*>"�>$_>ޭ�>4�������g>����*H��-��X;��5�R���a��5n�ʾF��ƥ�T:E>��>s������P	?`�>>=I>֎�?�)q?ʓb>򝛾�W�*����þ�嶾��';��6>���+jT��A��K�J�L��>ML�>':�>�H}>�]*�?	9�6��r�ܾ�1�@?�M-��H�W��|e�����z�����\��4<��8?ĳ��j��=���?��O?AWn?t
?}=۱���4=�l������V9�*�=��EQ�~@�>�?�?�<���V�3�˾k)����>�+H��O�̥���0���-���<�>�k���ZѾ�(3��O����sB��q���>�sO?e�?�a�'b���WO�}��+f��M?��g? ��>f�?�?�`��e-�K��w�=��n?���?�L�?+�>��7���=��*?�m�>
��?/�?H�?2:˽ʩ>uWX>��s��:k�Yĥ>�_ؽ�l>;H?>��h?Ł�>���>%�½۝��vʾP�ؾ؋�OHZ�kw!�v*�>�z�>��K>�-�=���=�\%>N�>�q>ͼ�>�ވ>i��>�-Z>�\���m	��c1?�O�=1Cq>�]%?�t�>���=�O ��P𽔱��rH�=�S��t��Z�{�Ƞ���<ĺ6>�S<���>�4ÿ�Ϛ?�M;>9>
���?أ�~4˽
� >��>���d�>���=A�=���>�ǹ>�Fn=,�8>0�j=Z�A��J�=�C;��r��`��=L�������>����W-�gா��F���T=���W��'�P����9G�.��<9�?Ȣ�K�%�T;c�p����f=?Z[?�i?k��>�ǽ#��=��u>9�=w�Ծ�/������K��jj?7Q�?�sc>R��>��W?��?=�1�=�2�!WZ�4�u��kA�m(e�Re`����d���ۍ
�K½�j_?ؾx?��@?h$�<7�z>k��?
�%�?ꏾ�ދ>�)/�r;�L�C=�f�>̏��P�^���Ҿ��þ��� �F>�o?���?[�?t�T��hZ�٪k>"�C?:�?4�?�f<?�K?�J����?�g�>G��>�9 ?]�A?�7&?q�?���>_J�>/y;��g=ƞ��\9���0��x��F��_=R\���>tG�<�3�<0�|=� ��� �jh��m��<$�<Z+�=d�	>
|= ��>Ts]?�}�>Z��>`V8?�9���5�(î�K�-?�92=����:j���P��@���>�j?�ǫ?e�X?��`>�C��A�J>�Ǌ>D;'>��Y>闰>��ｷPB��0�=��>t�>,Q�=";W�Rf���#	�����O�<��>3?9��>%[a�D�l>�x[�~���y�z>���a6����X�9�$�*�[��}�?,!?�pH?��}=��~�����g���4?*�F?�Ɂ?c�D?s�>%�@����.�����0�������ܨ��Ű��{��5��/^d=�j%>��#ن��4}>K:�`��͉�
,z�J-���>i0�o.�#����Xɾ�w0=B=���>��ǽv�*��2���Ѡ���V?u֎������Z���O���� >$e�>���>��ּ�m��s�s�
��/=��>�~w>�=���UB(�)W��e�>%�-?�Ng?���?}�|��S_��"6�ɋ��ݦ���!�?e?�]�>��?��>��w�����Ϯ����Q�2�>�$�>�y�>��,��Z��)�����u!����>�e?8h[>��?�u?���>�5{?�I;?*,?���> 6���K����3?��j?�=I�)��ý��!�:�=���>��4?��'�3��>��-?MP?��??f0?vG,?b�$>���5��B�>[>�>�s��N��>ߧ>�K?SH�>	�0?��?���=r;����%���&G>�G�=ed??Y�>t?�>���>��>����<6�=��>$c?�1�?_�o?�`�=��?I�2>?��>�'�=���>A��>2?rPO?#�s?n�J?,��>�V�<.���)e����s��VP�˅�;�H<c�z=����us��#�?��<�A�;*����h{�`��b
D�-��,��;V��>��t>�����0>��þ�f��lVB>���S>��H���@q:����=hŀ>�?���>��!�+��=���>]J�>k3�(?k?�?s]�9-Xb��+ھ�K�[P�>xEA?	m�=-�l�^����u�a�h=�Nm?�D^?wUV�@�����b?��]?g`��=�8�þ5�b����O?g�
?�G��>��~?��q?4��>l�e�/n�$��@?b���j���=�u�>�_���d�_E�>�7?uH�>a�b>[V�=bp۾7�w�g��?g�?V �?=��?�*>��n�70�a~羷����e?�	?&T��c?��<�hྦ���q���J�*���s��������ȀN������/5����={�?�^I?(�n?�T?"5�_L�?4O���{���R�N�� ,��FT��IB���Y�];x��y�τ	�鸯���`���|�S�A�~��?�X(?�5����>�[�����;c>>����� �<;�=�I���=�4=�=i�{3�Nv��d ?]��>\�>F�;?��Z��.=��#3���8�����a,2>��>���>��>
�*��5��꽎�ʾ����۴ֽ��s>�M\?Y�L?�ut?���oh.�05����"���c���{�� p>2�=Aa�>��6�o�%�$F!�:�0�2;g�~m��q��n���o�=L�4?�5>O׹>Wz�?��>I���Ͼ�C���N�&�><��~>�X?�@�>��M>kA���4�O��>�tj?�4�>��>dp���!�g�|��ٽ���>g�>-�?�*u>|����U�S��H��|C4����=�,h?����;g�5r�>�hR? �v�}-=�=�>���&w%�ki����M�Η�=k�?�c=��3>�;���~�Ի��<IF?�X?)����yt�dw�>��j?޸�>pB���?M��>g ���|>�?R9�?G0�>�I?�p�>rE���U�I�0���"R\�7�>�w=A�=�3>��R�6����!=k�|=--o=L6н2+Y>�wʽ_�=�N��Z�=��ڿ��L���ɾJ{	�����V�����

<������9�WZ���G���F��9����=G���j�rl,�6Qe����?��@K��B23�/���"-���S)�8��>wo��a�?��˝��η�U�z��3��칕��� �9L�����X}�{�3?�K���uĿ١��WX����"?��?J�x?�9���:������=��=�3�F��	�v��ٿ������_?�v�>b�� ����N�>TG>٘>e>����~�_���=�#?	\?ϧ�>�5�oͿ}��H
�=5��?T��?|�A?Χ'����^�I=7i�>J�	?�;>	�4�0C���� �>��?�Ҋ?�Sa=b�W�	u��Ke?��<��E�F���X�=_��=N�=���WN>y�>��!�� C���ؽ�A1>f�>�y�_��{�Z����<`^>yMڽ�2��5Մ?,{\��f���/��T��U>��T?�*�>R:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=s6�쉤�{���&V�|��=[��>b�>,������O��I��T��=���vѿ}:��m �H �=2��<J��;��,�Q�1��L�����Q*��M���
 �=�A>���>-|s><I�>)7[>�h?��?j��>ĕ>J�X��G��M�ྂq�^�>��H��4���m��U��aT�_W��=��)!����؛;�<�t�=unP�vȈ���.�`�o��rL�Gk6?vJ/>��߾�mB���ڻ�����m����5=i�i�B�о8;���q���?�1P?:�����@�����k��e�2���Z?����T�D@���^�='3<��=�ơ>��=�ܾ�D�/[�ES3?��?'�ȾOo��=�W>h �h��=j�?���>f!�;[�>��)?oP�����>rX>.��>��>6�=����ۙڽ��3?�f?�y�� ���.�>S7��4T�����
�=��H��Ϲ��>]�)=�r���@/=�r�2螽�*W?��>�)���PN���O�� ==��x?�?��>�mk?8�B?�E�<�>����S�	�Ǧv=��W?bi?�>Є���о����3�5?Ϧe?��N>��h��龎�.��M�?(�n?U?�-��Ys}�_������i6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>�������U�=�\���i�?n��?�����tp<� ��3l�!����<��=?��ſ0�n��C8�xrȾ
�
�]���ݳ��O�>3/@������>�i6�}��jϿ�����Ͼ��o�{w?���>э̽T�����j��u�Y�G�t�G�c
���&�>��
>t�{����\'x���9���μ�;�>���χ>�HD��"���Ț�L�<oh�>p��>��>�d��a콾:��?�X�=Sο���> �̲T?^�?��?A�#?�-�<,�t�<xW�Qᑼ�K?��t?��[?�����W�Q'�/oj?���A�j�/�<�-e>��h�=��?�/�>�,�k�=�B�>;��>���x��o�ƿdŪ�Xr�W�?���?� �{��>��?	K?�P�5y���誾$!�pȡ���R?�O>����O-� �0��@�n.�>~�b?�V��qӾ]�_?'�a�R�p���-���ƽ�ۡ>��0��e\��M��Z���Xe����@y����?E^�?e�?L��� #�e6%?�>e����8ǾH�<���>�(�>P*N>I_�۲u>����:��h	>���?�~�?;j?��������1V>�}?�M�>C�?���=�G�>�A�=�尾H��R�!>y��=�S@�#Z?��M?�j�>j�=(7�?�.��E�u�Q����	�C��0�>�b?Y�L?=]`>������1��� �q̽f�1�W���@��u(���4><=>��>�FD�u%Ӿ��?Qp�8�ؿj��5p'��54?0��>�?����t�u���;_?Az�>�6��+���%���B�[��?�G�?4�?��׾�Q̼>8�>�I�>��Խ
���d����7>5�B?F��D��l�o�E�>���?	�@�ծ?Ui��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?hQo���i�B>��?"������L��f?�
@u@a�^?*�hֿ����_N��P�����=���=Ն2>�ٽ*_�=��7=��8�B=�����=t�>��d>"q>=(O>a;>��)>���Q�!�r��\���S�C�������Z�C��Xv�Xz��3�������?���3ýy���Q�2&�(?`��k�=�([?�N?�2q?#�?����6>t����=i/9�wX4<6I�>8�9?�y>?T�0?/�e=�䀾%�Z�}B��Ϸ��~����>L)C>,@�>s.�>/�>L#;%�O>Z]=>�g>N�="S=V/"��jG<�)*>�ѝ>V5�>	��>�Ŕ>/��<X����	����i��n���'c��ʫ?˲���N�i�}�` ��(���#���>?1$�>�����ο{�����:?䶾F��rľ��>%�H?�.e?��B>�
���=�R�z=�i����K	>��.��ZL��CD��>wF?�L>�W�>d�3�TT.�>W�������>>��>?�A����R��m��L�W�ξ��J>^&�>�3&<�R�ږ�C�~��BZ�� [=��0?�?�E���ɡ�mz�I���u>nh>��8= �u=�f>�ȶ�b��57<�	�/=ȹ�=�s>(+?��1>�=AC�>�(yO��>X�9>��%>��=?o7#?�!
�UԊ�������#�� y>R�>u�>��=R���=l��>vUk>�m)�\�x����>�� _>�І��b�w끽���=��ծ�=4f�=1~��7<�� #=�~?���(䈿��e���lD?S+?b �=+�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��I��=}�>	׫>�ξ�L��?��Ž5Ǣ�ɔ	�,)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾOh�>x��Z�������u�ͷ#=`��>�8H?�V����O�j>��v
?�?�^�ܩ����ȿ9|v����>T�?���?i�m��A���@����>5��?�gY?8oi>�g۾`Z����>˻@?�R?�>�9���'���?�޶?կ�?KI>ˇ�?[�s?�k�>�4x��X/�r6�������=�e;�~�>�s>�����jF�9ד�yh��;�j�E���b>v{$=^ �>����+��R�=�S���V���tf����>&>q>J>#j�>�� ?!|�>Ǩ�>u�=�Y���Ӏ�����(2O?@�?�K��u��\�=��#>��6��'�>j�6?��<*þ�h�>	W?�p�?�U?�ͧ>[��7���񵿿�����R���~>�6?1"�>�0�x8m>V���"��?#E>�T�>�R�^Iξ�苾�]�=߮�>�8?�9�>\��;�j?�h?���>YЬ>����{��d��",>��?`X*?G��?�(?�9��C����d����C_�a�?�]�?��>99�>͉���9{���=u����v��Gf?�5?��W=��X?�G�?�
M?���?��>s�>����䗼�~�>T�#?�<���D�/�,��e��? ?�;�>�O�x�����bY�P�?��Y?�5'?�O��`�1�����<<���k2����9&����h0>{8>>[ǽ!�=��>��=�]v��<�|k�<��a=T��>)�=a�	�'T�r<,?};G�|ك�n��=�r��vD�O�>7?L>���b�^?pn=�\�{�K��fw��\�T����?���?j�?�#��{�h��$=?��?�?D�>�F��}}޾���Aw�f�x�Ox���>���>�>m��
�>�������E��`�ŽmC��e�>��?_ ?غ>I�2>���>+ꂾ�03�-!��8�~����^�J���J��|5�!>��wч�L��#�����q�>�A5�5��>��?�6>�z>�ߦ>(�NR{>�&`>$Oz>2{>��>��K>�ߣ=X��:�D�4NR?K���(�'����c���L=B?jd?��>��g�=���;��,{?鄒?�q�?�v>�oh��%+��d?�1�>��Qm
?^w9=V��2�<oI��2��
����K�x��>X
׽�:��M��df��r
?U"?~׌���̾0׽�}��������?�Z*?��,���#��Z�f�[�4�1�Ro1������;L=��G���*��v苿�*r��*��>��0?΂r?��C;u^��:l�e�b��q�=�r	?#մ>Z_?��z>���0d,�D[Z���i����?��h?L">�Zp?�@,?�L?0�M?��>s��>�ԾĽ�>���������>��a?!o�>9lS?0n�>��I?ӻ0>5
վ�>0��Q���7?��>o�&?��>���>�����L����;`̽dBS�d+��~��(��C��{��:U�;�"�>��?����9�����$�h>ݗ7?���>���>�����G��|��<:n�>�
?���>2����q��?�,��>���?���ػ�<I1(>_K�=(ˈ�׏���u�=7�޼5��=�my��A4��<9[�=T%�=w��<�:���(;��;��<�t�>��?	��>D�>~@��ة �����a�=\Y>KS>Z>�Eپ]~��
%����g��Wy>3w�?�z�?G�f=`�=���=�}��vU�����?������<ƣ?BJ#?XT?���?��=?�i#?H�>�*��L���^�������?�Z,?3��>����<̾鮨�U�2�ff?�?�`�+r�m(�F8¾�F׽̹>�/�L�}�\%���(C��9��g���)��LM�?Ʊ�?pt>��7��JИ��ʬ�BD?�8�>�[�>���>ZZ)�\�h����_?>�p�>U9R?�x�>%�<?k�k?��\?�T@>��Z�����v���J�=^��>b�?�9�?�Mt?��?iȍ>��>�䑽��C��J6�ث��x|��8Y��^6>�(>i��>t��>'��>�v��8[��M�g��é�פ�>�ZG>�Y�>�k>�?�V=�A��H?���>3P�������؂���?�Ou?Ϻ�?P+?=�7��E�����"N�>�j�??«? �)?�T�o��=;�Ӽ�R��A�r�R	�>E��>�J�>��=V�I=��>���>g��>����F��e8�'�P�L�?+�E?�˻=	�ſW�p��Rr�6���6W4<���g�Y$����]��Ԣ=�:��x�{��� �\��D��٥��t ���?���{|����>�w�=ֽ�=_��=���<�μ��<��F=���<�Q=�fk�E߀<ճ0��}��7���h����B<��L=�w�־m`~?-'M?o�+?T?�&�>:?b>̭��9X~>��P���>c�<>9.��伾l*2�Hw��F�S��Ѿ��оUat�؊���P�=�L"�w�>��'>�=��0�v��=�J>fP�=�K��V�99��=�6=�"�=��=�g>��9>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>2^�=�4>\�T����Y��x�����Ǿ�D??�>J�rvվ�t>C,��.I���Ⱦ�2�=�h>�i�:�ـ��U�l�=��˽y�d�^��=��u>�#7>�=ܰ۽�����=�>��A>��=o��(���=��=��=�Y�>z	L> ��>�?�1?�a?V��>`l�gY;i�����>���=�?�>�Š=U�@>�ʻ>KE1?g�B?9�K?A�>}{=\$�>z��>A4�fts��Ҿ?y��iU<�)�?���?�*�>�6<h#�R�ޓ/��/�?��.?s�?k�>cS�M�������+�D�7<��c=�[>�s����N�KId<����	�TBI=�!�>���>{�>N��>�5�>Sb>�6�>�=>�e��X�9=K)��י:���<�!�4>�>a��μ<k�<4۽\⼽U=կ>�:�==VZ�Sb�>}h�<��='�>͍[>cD�>iHj=t�۾q�>�J��3:��:i����>A�	�c�n�f�z=�)���Q�4>��|>��=Е��OB�>�g�>�_>^�?Wl?d�>b�����M����𾉮��朼oӖ<�#��K�c�T��[Y�	3��4�>`>r�>�Xy>�"��G���={�Ѿ��"��k�>�9�U���>���f�5f��Z#��x�Q��]�=f�U?Ͱ���B>O5�?��T?'��?��>B��<����U�=�)���-�i	�Ҁx�.M�_p?s&	?8�?Jݾ�HS������T�>����K��P��w)������ž���>�阾9*�r'��`��$Ƒ��:���b��x�>�>?H_�?�;��"��GV�y�vH���=�>��l?b��>��?�?�y5=��龃��[�>��j?z%�?�U�?$-2>𢍽�@�<Ƚ?5>?�-�?�W�?�k�?�퀾)�>^8�>��	��rg��NJ=+>���=߳{<�>?�/�>�x? |޽�5"�%w美�?x��[#=ʈS=�L�>��w>���>��>@o�=̦�=r�>$Y�>���>{��>���>tW�>���^���΂4?E��=?�R>��<?���>>�=����Ž'�K�6�0��j���$�.`�u=�.� ���C=��=i�>��̿�#�?h0>�����&?�]��l��A}>��>:���8p�>>�~=WX�>�ϯ>��=$�p>��t>DӾ!�>����`!�j/C�8�R���Ѿ��z>࢜�!&�7�����6I�uo���b�j��-��w==����<�E�?������k���)����/�?Y[�>�6?�ތ�H���j�>m��>Hύ>^K������wō��gᾷ�?t��?oBc>���>� X?@�?�	2�S~2��;Z���u��FA�N	e�ho`����n���
��5ýǊ_?��x?�A?�r�<%{>H��?(�%�Q��׋>/��;���A=�ȧ>p���_��,Ҿ�þ���m_G>�so?]=�?פ?%U��{��+>�;?��1?'lu?�Q2?�d<?1��'�#?��0>�B?Y�
?[W4?��-?��
?��->}��=�ûW�"=�&�����Qmѽ�ŽV�e�4=g�=����!7<^�*=�Ҳ<���}��m؞:�Լx��<��9=]��=Ұ�=���>�w]?L��>�Ѓ>�:8? ����7�u���80? (9=g���퉾@������9�=_�j?c�?�X?��`>wC��sA�>`��>[�%>-�_>��>	~���C�S�=��>x�>�{�=��S�����
�����,�<��>2��>r_�>�n��h;>*��1�v��Y�>cP�x�;�}[���A���$���C�R�>�(Q?�?��>�ھ��"���j��0&?��A?�NY?�U^?5�=�Ӿ�1��5��X;��q�>������ݔ���a��v5�c���Kuf>g���H�z�5OG>y�$���澎�u�xS:�� 쾻�$>���~n��8��c�Gq��Է�=�3�=�4���� �5H��ݜ��!4>?��=HE�T@��xݾaSL=&Y�>w��>$����o��o:�؍о:
=l8�>��>=f�=�e	���B�):�l�>��C?�`T?�`�?S�Z�KȖ�F}Q���ϾjN��b����%
?�>(�>s8r>-)�1�վ9�۾<Od��C�y��>��?]=��S~����"*��U�D���Y=�l/?5^W>�>�`?��>Z=&?n��>�?ķ?�pE�$L��=�1?7X�?j�>I����?�����pT�!�>0�?�@�{��>�o=?��-?�?�� ?��?4�>mq�m��ꌃ>��n>��K�ְ����I=��?��>�6?-�U?�:>�G�𞾾#ʽ�@�=>K�>>J?X��>�	?z��>�6�>���+��=�	+>��$?nu&?(�r?E+� !�>TY�>s95?�?*��>K��>�C?�R?<�p?��h?�y?`�;(����$���^� �~=�;:��x�=U��;������9P��%>�^>�W������u����(0�-�-�_�p;���>j�s>���ը0>��ľr���>@>�����&���P���8�4(�=��|>h{?4�>fn!��F�=�>��>�D�HE'?�?ɢ?n{��d]b�B�ؾ��G�."�>%�@?�8�=�l��Q����u�P
b=�wm?7+]?@W��e��7�b?�^?E!�Y=�ܣþ\�b�I�� �O?��
?*[G��˳>�~?��q?���>�e�;0n�l���Fb�d�j����=x�> \���d�0�>�7?�4�>�Qb>E��=
�ھ��w����Q?��?�?>�?I�)>A�n�c"���𾖋��Z_?��>�F��� ?���,I��.��ȼ���վ桧�P��������􌾐	6��H����̽�y�=T}?��r?�4s?�?`?&��c��Kb����ږX�6\
��2�YQE���F�E�>�n�w����������t=��d�oK��2�?��)?�����>K���
�����־��u>2Հ��.�?y�=�TǺR�>D�I;�w�]�,Ʈ�R?�3�>���>D�B?�}D�=�=�*�9���6�aX	�x��=�j�>��]>2��>o�<h�'��D��{˾����BHjt>�LW?��>?�K�?���>&(�������2��[������(>^�'=Ҳ�>d�=�d��x?��Y��c����)Ty�p)���Ի=nN?@D�>�֋�Q��?C1?]8���������.�8?�\�Z>-�2?}7�>[/Q>�Y7>������>
�l?r��>��>�����Y!��{��ʽ�"�>�ݭ>��>��o>̯,��"\�bj��&���9��u�=�h?�����`�b�>�R?��:ݡG<H{�>Ыv�A�!�o��a�'���>�{?R��=֚;>a~ž�#���{�7���u*?ܮ?�|��Q{6� �*>�'(?ҍ�>�6�>,:y?�Ւ>�=���"�=IX?��U?9U<?c�M?���>a�_<�0/���˽ѣ8� ���%�a>�x7>�Z�=�>/>bս\lh���J��x�<҂�<�1U�ȤٽI��;��`����<�cX=p�>V�ۿ�I�9?�Q���a�g���B���%�.W1���
�`�~蟾�����k���j���x�
�e���P�<ʃ��P�?CZ@���X���G����P��h.� ͳ>Z`�t#�;��þǉ�X����"�ܾin"����O�Q��'s�Q�'?�����ǿ𰡿�:ܾ9! ?�A ?=�y?��=�"���8�� >C�<i-����뾨����ο=�����^?���>��/��p��>ݥ�>��X>�Hq>����螾�0�<��?2�-?��>��r�-�ɿ]������<���?.�@}VD?������(>)��=�>��?�@>�%��w�C&��xn�>.��?�Ň?f�a=f�U��-+=Ff?4m/��.�L��
7�=�i�<o�<*R���z>RO�>@uͽ �G������=g�>bi���7�'�S�j�<�C>0┽����Ԅ?Mr\�df�(�/��S���>y�T?m/�>7�=`�,?@H��|Ͽֲ\��a?�*�?��?-�(?�ܿ�Fܚ>��ܾ��M?2A6?��>l[&���t�0��=/d��������(V�i��=��>$`>�n,���\�O�+������=���pͿ�o6�z?$��к��\=�p�<p*��}�;�,�VX��B��5�V��ٷ<��=�p>&{>l�>v�E>`�^?�}?��>*E�>�ֽ^���́��K��Ԃ�Ft�豬�����Xp;]p�f�Ǿ�G�~�6��D<����9�)2&>a�c��.���'��a���6���?>(�>.	g�JL�u u�V�ɾ��-�-Z����J�wt�􀇿��?��Y?4Ֆ��W�2��ͨ���@��br?�P�<g^��Ez��\=�b>�\�=x>�Bo>��{��i�u���0?��?�I��%��w%>:����4=p�+?	c�>�
�׸�>��"?�4�����V>�50>sc�>��>�w
>%����`
?0PV?���/��@��>e}��~���H;P=�X>��*�f�+�T>�-<�<���u[��r^��p�<DS?�э>�O���!�������=tq弣ւ?,��>��E>�a?�:-?H =Q����zJ���R�>'
J?�pZ?u�5>���#�˾p����1?��\?l%>��$�����"3��4��.	?�3?C�?��}���n��ܝ�<���
P?��v?pr^��s�������V�K>�>[�>���>��9�Mi�>��>?#��G�������Y4�Þ?3�@܍�?��;<$����=�;?A\�>ѬO��?ƾ�v��-�����q=�!�>�����ev����R,�ه8?ˠ�?��>C������> ���=��?�?�$��۹��z�m=���"�ϲ9��ɀ=�	���_��ɞ��7�X� ��������BһC�d>��@x�ֽB�>F����˿�xڿ���cǦ�����i�>es�>Vt��= ��6���`j���B�z�Z��-0�S�>Zl�>w;�&پ����(������?�w}>��>��v�wҾ����L�>��>�5?T�=m'�mM�?�,�@ο��~�:�����r?oxs?i��?ᖪ>�M<���'���N����N�.?��f?_�F?��ɽ�Ɨ�dIv>!�j?�K���`�?�4��^E�]�U>9�2?���>c�-�D�t=�>��>�>�/��wĿP��������ɦ?]Z�?�&��d�>T��?�O+?R���:�� ۩�ق*�>|�`�@?��1>������!�O�<������
?,�/?���Y�M�_?�a�+�p�y�-���ƽpۡ>��0�f\��J������Xe�����@y����?K^�?]�?���� #�u6%?�>U����8Ǿ[�<���>�(�>�)N>	H_���u>����:�i	>���?�~�?dj?񕏿���� V>�}?�"�>6�?ڌ�=Au�>x��=a���i�,�1f#>���=|�>�i�?�M?~F�>�~�=d�8�� /��]F�,DR�W���C���>��a?�~L?�@b>@,��2��!�upͽ�S1����T@��,�x�߽z5>��=>j>�D���Ҿ��?Gp�?�ؿ�i��Jp'��54?��>�?��Դt����;_?1z�>�6��+���%���B�W��?�G�?;�?��׾4Q̼�>(�>�I�>�Խk���{�����7>*�B?v��D��f�o�b�>���?��@�ծ?hi��	?���P��>a~����U7�x��=��7?�0���z>���>��= ov�һ��E�s����>�B�?�{�?��>�l?��o�G�B���1=�L�>��k?�s?�.o�D󾅲B>q�?!������ L��f?�
@ou@B�^?��Կ�=���w��Z�����=V�=� [>1t��w�=dKe=S����+<�b>i��>��W>�h>�W>y�R>�p>���nO#�U���$J��qA������b�[�P��`%p����Ȱ��Ǿ�>���B��������C��N��W���A�=�)I?j�I?Wa�?]2?�T/��>>d�޾������	;!>[��==�'?o�M?�d?7�����̾s`Y�weh��Ο�Z$����>�R>A[�>�/�>�ٴ>	�='{ >U>9��>��=ò=�����;A�L>qL�>fz�>���>\-?>M>bk��h˰���h�Z�r�B�ҽQ�?�)���L��!���ҍ��/����=˕,?If>�x��_Ͽ�1����G?������r	*��(>_�.?�V?o�>�a���X�׃>���$%o�B�>c��"Ze��+� 
M>��?_�>Ϯi>/�9��Z3�]�p�_Iu����>� h?�쾷оr~��cj��s�����bB>Y k>P�l���(th�򊋾(3+=��d?8�.?,����������N����)>��Y>��Լ=i�=�Mm>��W����S�;�����e�k*�<�\�>�R.>N-6>́�>ي��a���D��>��=��c>x�P?�%?#���ݱ���h�>TP�2�H>��>(�>f�P>��[�4
y=���>W��=�5:�Ə��LF��-߽�>}�;�N��V�μ�ܻ=ё�=�п>��r��;}�m��^o>�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿfh�>'x��Z�������u���#=Ψ�>9H?]V��V�O��>��v
?�?�^�ɩ��y�ȿ�{v����>0�?���?u�m�wA���@����>!��?UgY?�oi>�h۾�`Z�͋�>��@?;R?�>�9���'���?�޶?���?�O>��?��r?�$�>զz=N*$�~t�������_&<L�ứbB>Ps�=b������𾆿�D����s��a ���T>po=a�>D4��羲)�=�?���־�&m��n�>!�>��>�@F>�:�>I��>���> r=-��<������؃K?⭏?����om�)��<wߛ=4�f�B�?�4?
���gо��>��[?xw�?��[?�\�>V��or��d���.��X��<0K>��>m��>F_��F�I>�վT�B��K�>���>����=پ�o��h���Λ>�� ?�>Ʋ�=�� ?��#?��l>k�>��D�~璿�F��>m��>а?�~?�?������2����Ip���Y��xI>x?� ?ז>� ���
���_����@�y4����?�h?*n�Ty?���?̈́??^�@?�_>P���Ҿ�뱽j�~>�Y'?�h̽;VR�;e/��}S���!?���>��?I۽�c����X� ���� ��>,0=?}l"?sE뾝KT�����s��<�X�sB!=��=̅<0�V=�;F>7w<��;��=��;Q��-���nR�Yv�=��>�B¼w�_�����@,?b�D��܃�^D�=/�r�QID��>OnL>)�����^?��=�L�{����Iz���U����?U��?!^�?I���~�h�^=?��?1?./�>ok���f޾�`��@w�b�x������>���>�hq�����&����E���ƽ����[�>�m�>�@?���>��`>T�>�i��0����澈�̾�'4��$6��zT�$#5���'�-.����=X�ݐ̾9HV����>����Я�>#W�>%�p>5`-=�?�>C��>�p>9>��w>]C�>�@�=��w>$�2>��=>Ɛ�NIR?Գ��K�'�i���ڰ�.NB?Od?�T�>�~i������X?rd�?WU�?�u>0Lh��+�+U?ZG�>����F
?�:=W���<	L��[2�$T�����0c�><nؽq5:�I1M���f�+S
?�?����̈́̾�׽�j��)js=uC�?.})?Y!(�B�Q��,p��W�US�&%�ˏh�ٍ��$�aSo�늏���������(���1=!�)?�k�?������I����Jj��Z@��y^>���>��>uҼ>�I>����I1��^�9�&�̋���O�>%=z?>�;B?N�>?pFJ?�??�y>��>�t��D�?�_�=Չ>'�>��7?�"?�8?f�?O?�E�>\b������lӾK�?}�?A?�?s|�>�m�u'm��w�;㋽�n�Upɽ���=>��=�>�10潅�Z=��Y>�\?�?�\�8�������j>+�7?���> ��>+���B���
�<���>W{
?9�>����Ir��6�t*�>���?
3���=��)>�"�=�[���g���=Fm�����=�=�� �=�J<�%�=�;�=P�b���)�Cǿ:a`;	��<<��>K+?�;�>cs�>�톾�z ��	��t�=�qU>^�Y>V&>�!پ�r��hė� �g���v>�?��?�W=1��=z��=����G�����#k�����<se?�!&?�V?��?Y�<?�%?��>����k���$���օ?�c-?PR�>���>-��@����=�Y?dD"?Hh�E�b�=�&�Z� ��8�{��=c�1���8���A�	���F�������?� �?��=�F+��ꦾO�����r���J?���>���>�L?�,�1	O����bB>���>�Y+?o��>J�[?�i?3Y8?���>l�pq���饿{�=���>�d ?�w?{o?��?��? �C������	5� x����'���CU���&>��y>�`�>���>2�V>הU=�OS���(�U/ν�%0><�>���>��>7�>�w=��=3J?�|�>ҕ���'���ɾJE�Dw<M:c?���?,�?	H�<�7�b{>���?��>^٤?���?��?O�׽ګ�=���!xѾ�`3�pA�>gs�>,�>	P(>���<�I�=��->Ӧ">p=��q*,���!�c����>�~A?�Q=��ſ��q���p�h����h<�Ւ�P�d����T�Z�\q�=���bu��詾(�[����������뵾sZ���W{����>E��=/ �=��=���<�}ɼ<�<&HK=�"�<�7=��n��o<8�w�һm�����_<��I=����4�þq�u?�AE?�E%?�=?&�}>ѢE>�^���E�>&��a<?�/G>�������dKO�����G��οϾǫ�i"m�xD��`�>�����@>��0>��=�j(=&��=�3�=�� >n5^=dz=X	�=���=��6=���=��.>W�>#5w?���S���|3Q�V�<�:?�#�>W�=7�ƾ�??3�>>@3��n���G`��?���?{D�?��?��i�Z�>� ������8��=<m����1>��=��2�G��>��J>���M������+�?f~@��??�䋿ښϿl />�Q>�|�=jNg�x�0�b�~��#!�u}�a.?��9�����a�>��=�a��Ǿ��<]fD>�	�=�M�#M��Y�=׍ǽ�H�=�ҋ=���>7�>*8�=�������;��c<��=]�9>�ֱ�7ݽ��=����=�ʻ��1>p�$>�q�>R�?�S0?�t?� �>ɺ��
KľOz���E>���=J��>�[�<��4>���>�!.?�1?�8?�l�>��=�n�>:�>l�#��xm����B뫾�'*�"��?I�?||�>��
�nG��^��o�I�����?7�D?���>7b�>P��6����&9��?��C��xv�=���=�b �u�P=�Ƚ�M#�EŜ���~=���=���>���>���={0�>C��>z��>�>������럱�)}>�c�:]�=�6)<4Oo=Љ�~��6��=v�<2�ǽ{�<��U�
<�<z��6�=~��>��(>^g�>�Sw=I朾O�F>�M��N�=� �=M[����A���c��,z�{�!�>�G�/2>��_>z�	�L������>$>G>k.>��?�t?Ut<>���=�Ҿl⛿���9�i���= ��=��J�UQ>��\���H�]پ'a�>��>Lx�>�r>Q=*�ѐ>�=/:��W6�r	�>�k���+�����r�m���B�����e�c��`~B?�/���p�=u�~?cOJ?<�?9�>YE��JG�}�'>|�y��=7=���+Lr�lח��q? #?\��>/jܾ��D��;Cຽ��>P�K��O�����>0�k4.�=紾�w�>+0��7�о�l2�jY��f���UB�xFo�[U�>n#N?�P�?8$Z�������O�TG��1��E1?��g?�&�>V�?r�? ��������~��m�=��n?��?��?*>��:=o�1�.��>���>1�o?m?�u[?�:n����>U>�m>�>P.��R���m�=�`=&�	?0<?+��>v�k��1����v��������7=<'�=z�>ˎ�>�0�>��=l�=A��=�0�>U��>���>&�q>���>��>�+��o��U?�=� �>Z"-?��>�4H>e��D>�@��Y��je�zu�we�<MBN�n�@�ɝ#>�_ɽ��>,jɿ|��?M��>è��Ԣ�>��	�Xb��Ȍ=q�>^m��ִ>q��=���>[��>B=>���=�2>�Ve>�EӾ�>����d!��,C���R���Ѿjz>����$&�����x���AI��n��Cg�j��-���;=�ν<H�?������k���)� ���0�?[[�>�6?�ی����z�>g��>�ō>J��.���'ȍ�Ki�:�?*��?�@c>D�>��W?��?;�1�B"3�)dZ��u�$A� �d�1�`��ݍ�2�����
��?��d�_?��x?�wA?��<c+z>��?��%�$׏���>k /�v#;��_<=�D�>	���a�q�Ӿ��þ���[uF>��o?b �?AU?�%V�cuR���>xw7?G�'?�Sl?�*?x^A?
��M"?�`I>�H?��?�:?B�%?� ?ɾI>�>>��:�Db=����و�V���ѽ�]���/=�)�=J�<m q<���<o(���U�����g�;k���3: 0=��^=ө�=`n�>W�X?��>�&�>"�0?��!��C.�cx��aW4?H�=�ތ��놾�[���R�O�4>� _?�ͥ?�|[?PZ�>�qH�sDB� %>q�q>��7>�Aw>J�>��߽�P-��-=u��=v�>S$7={G`�]i��!��\���,}<��>7�>��>�㻢�g>-���舾9��>��
��a���L��i�K��B$�|ʒ����=eD?gn?ؖ�<��v_���o�u?�JI?�&R?��?��=�A����R���g�ٽ��?:d>��Ͼ�T���1���cF��?>i)�>}t��Y�~�@�c>u�2�Ot�>#~�,�;�����=�k�����;�[���*���_��՜=��=[[׾ ��������MG?G��;:̖��Q��'��+4�=�q�> �>�L}��^��y@������;z�>��!>xg��!2�gJ��Yپ툤>��=?yQ?��?�U2�0��C�9�����侔[�=�?�>v��>P�={��<�Ӿ�t��g�P���H�l��>�5�>;S7�*�d����-����O�q��=�f5?b^<���>P�?�<?�N+?�@�>�?�m�>�ց����-5??+�����`��^��!+=�Q:K�܌�>�?�4�����>y�<?�h6?�?UM ? [E?�	�>��7��uB��7�>��>��W��{���3Z>��z?�g�>!�A?ڌd?���=�iE��Bξ�}����>�e�:~-D?wM?�-�>���><��>P�����=�l�>��\?1w?�+w?�}�<���>b�>���>��>s�t>V�>f�?
N.?/�n?4�P?�`?��:������J�����D���=|o=	}����V���j�=��X<�H�=ս8=�m��P�,�#u1�w~�=S��>��s>ؖ��Ku2>�
ž����f@>3���jٜ�_J��� :�j�=~>��?tD�>un%�Ў=�Ż>m��>���E�'?�t?�?��j;: b��eپ�hH��>��A?<��=��l�:~����t��9_=�m?&�]?�,V�E�����b?M�]?�g�<=���þ�b�&��?�O?A�
?��G� �>?�~?��q?���>�f��5n�d���Eb�a�j��Զ=*s�>�X�c�d��>�>�7?jM�>��b>�&�=at۾&�w�:s���?I�?q �?���?�)*>��n��2�0����U��&�]?�[�>2���c	#?�]���ξԱ��+�����몾\����U��a-���$�����Խ���=;�?O�r?�|q?q�_?z �`�c�5^����rlV�L(�	�?�E��D��!C��gn��D����K��= E=�V�W�E���?.?+>�H��>I􉾑ȟ���%��>g�����-�伈==�[����=�8�=J��e��¦��6k?���>!��>E�7?�eI�6"F��ET��ER�O$��=;��><��>���>�F=F� �E��M�:ǥ��1�N�>�v_?XU?흂?S�;�=?�^���WB���(�\�оKą>� >���>�:������-��=��vq�(��}��E���i<wK7?Dz�>pȳ>�i�?6o?���WVt���E��0^���#�ɛC>�P4?= �>M��>��0=2���>��l?��>v�>����rY!�`�{��}ʽe&�>Wŭ>y��>�o>N�,��\��c������M9�%h�=��h?݂����`�t�>�R?O��:=UJ<E}�>�|v�w�!�����'�`�>�t?0��=];>�žM�&�{�$���?�H?4a�&�:��$b>z�?8�?Kw>���?�.�>,~о��=���>c�f?t0g?��?k�>��"�:ڨ�@�ʽ)��=[)�>Œn>��T<�ʵ=e��� ]��q�{�>:�>Ű�<�I�L�Y=}�����!�b=��>�ҿ�,;�1��)����&�ξ�^���ӻd�⽮E��yc��G����X������½{�����m���A�� X����?~� @���?���7����b��S޾"BI>�,��}�*>3�h��۽ �ƾЈо��|��*�vA=�V�i�4�i���'?����i�ǿ֛����ܾ�2 ?� ?��y?h5�@�"��X8��$ >^\�<�����������ο-���^�^?U��>t�Ѡ���>�M�>i�V>r`q>�W��jl��l(�<?^B-?���>�fq�)mɿgP���ȕ<m��?�@�B?���{> ����<F6�>�+?��>�L�$3��������>���?<�? m=Y%Z������d?�	_�bC�T��;���=կ=)u�<�2��#O>�U�>1� �)o�w5���;>�p>d_��C�b�M���'<)->�彟Z8�5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�����{���&V�}��=[��>c�>,������O��I��U��=���'�ϿX$���/�.<�=Ï��mF=�¼�P�@�����呾���� '�~��� <�>qs�>0�>±�>�%^?�ˀ?Ȍ>��<�Ҁ�y�@���¾��<zR�������^ѽ)�!���G��ݾcQ���ɾ�!�'��>�:�J�=�V�M���غ*�IQE��Y<�̼?j:�>BW����2�(����Ҿ�%;��;�P��z����k!�I�_���?�N?Z��5�C����3���w�i�1?�����־h�x����=��ҽ�>r=^`�>t�=P�ʾ�/-���H��8?�?�Ӿ�Ӏ��R=:�����=lN ?|�?6fڽy�B>�+?,�(��a�Z��>�d0>��7>4��>��;�,���*�T�>?N�?�8���Y����>�؝������]���=���;y|�P�>�d�<7'�)ϟ�*�=̧�=d/M?0��>a�N�S#��߾ۺ#>�7�1k?�n?S>t\m?:P?0�=+�� M������=��F?��J?�\?>K���2�#*^���<?Y�X?*gE>������T��
�?��j?��?��˽�U���Z���i���%?��v?�r^�'s�����V��=�>�\�>��>I�9��l�>S�>?�#��G�������Y4�Þ?��@R��?<<n%�(��=^;?[�>�O��>ƾV|������c�q=f"�>΋���dv����Q,�P�8?���?���>n���8���	>fi��bS�?!/�?��4�n����c1���Y�e�$�*��=ľ�=�Z�<Z�=�V��k��w����D�k���B+��}d>i�@�Z%�+��>��b�ݿ��ݿr����������n?��>���=lpP�����W�[I$���f����g>1��>�����x��w��������9�^f>9�>vR�>��=�/�5B�#�����>h�?��U>j�޼���">�?��;H�Ͽ��{���/�<K_?�>g?:_?a� ?*@��ۗ��Eק�Ҫ9f�T?@�G?*75?"��<b�"��C���gj?"���Hc�L�3��$G��a[>�t0?ł�>��.�vi]=>��>^L>�,�,3ÿ	���a�����?�"�?���Җ�>��?Z�)?=��,��}[����%�ӂq�ɒ@?n;>��¾��#���8������?"f)?$�?^��_?c�a���p���-���ƽUܡ>o�0�g\��(��ܣ�ZWe����By�T��?^�?j�?���n #�!6%?��>�����9Ǿ5
�<_�>
*�>�&N>xA_�߲u>n	���:�Qg	>���?�~�?|i?앏������U>a�}?�>��?�=I��>@&�=�����*��F#>�Y�=&l<��Z?mM?�1�>���=�G8��/�|F��9R�����C�O(�>�b?FnL?~8d>�з�ψ0��� �:�ʽ{s1��{�=�?���-���߽5>H>>�}>kE���Ҿ��?Hp�6�ؿ�i��#p'��54?3��>�?��|�t�����;_?Bz�>�6��+���%��}B�\��?�G�?9�?��׾�R̼�>>�>�I�>*�Խ����g�����7>5�B?I��D��q�o�s�>���?�@�ծ?\i��	?���O��!]~���d�6�H��=��7?�*���z>6��>��=�nv������s�3��>�B�?z�?���>��l?��o���B���1=FO�>�k?Cs?.q���¿B>�?ɮ�p���"M�Cf?��
@Gu@B�^?�ꢿ���������y^о�T>��>�#>�G��eMл�XC��g���a<�+���b>(�_=�W�<WM>��>jy�>}������^���L��/qP����as��m��Z���j���7���ǾO���v|�m�b�NX��d�m�e=�'�=LE?ɴB?uT~?ҝ?�?�9.>����푐=�ܧ=�.���A>D�?��G?�;-?��=��پL�_�-�e�����ugJ�FO�>+��<�t?�,�>S��>��=>��>�JW>�i�>xeE>�Bh��E��Ϧ=̿�>�n�>�� ?N9�>��A>��>�4��tʯ���j���c�T�ս���?-��]J��L���-��	���$��=$+?��=����*Ͽ竿�G?�Z����U�&�0�>]d*?�V?��+>�X���(I�Ի>�����y�1X
>���{Bf���,���S>��?��|>�#p>�oD���4�6�W�RY����]>^�9?m/����K��j��sE�*�߾gI>��>-GJ���7����ir�)R��+=R�@?13 ?a̯��5̾8�T���s����=�"\>jKu=}��=�=>�c��ꢽM�*���%�K�>� q>ز?a�+>b��=�Z�>��a�#L�7z�>�p>@�=d�=?��"?~������\y��\�.Z�>���>��r>���=Z4��K�=8�>C�9>�|��e�Ƚ�x��V�9�N>����e}����96l=�ǽ`m%>��=�&�ؿO�I�=�~?���(䈿��e���lD?S+?] �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�-)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�h�>_o�X]����z�u��X$=0��>q7H?	H��� P���=�;n
?j?']�J���4�ȿ'tv�K��>v�?���?��m��?��@�H��>F��? eY?�}i>I{۾FYZ�.~�>e�@?IR?��>S:��'�1�?ٶ?ԭ�?��I>MD�?R�t?FP�>:�R�u1�_���?o����\=�s�;�p�>��>S���߹@�ؼ��>u���j�hk�I�H>U�&=D�>{ ǻ��d�=>���,'���8s����>��q>�/>n$�>�?BB�>���>u-M=�I4�Q�������Y?�?�?�M�_�y��������O�Q���>x[.?X�	<���M�>��c?��_?&9S?�?��㚿�骿�ˤ�~i���Bh=�=?R!�>���8��>�ʪ�yJu�+<,> e>uq=��Ǿ���g>>}�[>���>��0?Sכ��P!?_�#?*bg>}�>k�D�Qi����E��ټ>���>�<?L�~?��?�ò�O�3������>����V�W�A>��r?��?�,�>������"���$�/}��Aˀ?f�i?m�
��?�?0D?J�@?�K>3�Ľ��˾}k뽅�y>+s*?��Ǽ��9�M5��� �Æ
?�>q��>�t���A�����)Ѿk,?4�??��-?�s�Bx�Գ�����<Ĝ:,�:���;�ة�X��=�h>>Ac�&�=V|V>1� =�z�0)��(�<f�C>E��>d��<3L��J
̼��+?��N��m��S�=��q�ѪC����>L;K>���l}^?-a?�Xn{�l��[����T����?~{�?9�?r2��	yh�s<?��?y'?6�>֢���r޾8a��u���z�ϵ��">���>�+�x�񺤿�쪿�'��>HʽR�j�p��>���>]�(?$�?|��=B��>D#3�sվ7��ap@��`���-�����H	�v/=�������Ƞ<f����k�D`>���X�>vL#?KE�>: >
��>d��=%�s=zG�=��3>��!>L�s;�y,>�.�>~M&��b��R?��>,�V�C4���cC?��`?Q)�>���\��U���f?�Տ?��?�=o>��h���)��?RJ�>��z���?l��=����R<x�����1H���`�i��>7���-9�e�O���W���	?��?«'���ľ;�ʽ]���o=�H�?w)?��)�'�Q�P�o��W�1%S�` ���g�_��a�$���p��ۏ�/]�������(�/�(=�*?D�?�������s��8k�82?���e>�3�>�>_׾>�J>�	���1�v�]��S'��Ճ�S.�>LY{?���>HLG?�$;?�<J?�^K? )�>���>Ᏻ����>,C<֕�>T��>ܭ6?�/?Z�4?�o? �(?�tb>`�������(־g??��?8?�;?k� ?�j��q1��n˼%��;u�i�J���=~<�T�Boy�	}=1�G>��?[����.�66���W�>�X2?qK�>��>"%���f���Q;�?*�>i��>髆>��t�w��,��~�>�"�?Mm�G]�<��>���=!N輒�%����=�I���=:2K������<�Z�=׶�=�[�<3!�9�}�oU�<���<�A�>��?�͋>�>ޟ��z~ ��v�h�=_�P>�ZU>�7>��۾\e��ʄ��jh���z>�d�?���?CWP=��=�K�=����N����������<(0?�"?)dT?��?W�>?��"?9� >�z�d����9������-?��.?D�K>ҟ)�胓����F'+�n2�>�	I?�ˉD��&��L#�Y��� ��>���]^����<��7�.���ˎ�<a�?��?a��<N�N��7����������T�a?��>�lY=3p�>�˶�u6��e����~���>z?,��>��o?g
�?̖K?��>1�p��zϿ��� �޽���� �>��?@�?���?�H?����<�j&�j�@�8q��=���S۽�N1�>�>R9z>�J>�F�>?U�>����cm�=�>G���Eͽ�	!>��?���=5��>�L>�ݵ=�Y>?��>4d������C�G�꽅XѽRCc?�?��?�w>P,)�_@���<0�>�p�?AI�?�_&?KZ���(>lّ��^׾��<��>0o�>g�a>c>�$Ӽ���=T��>1ڳ>���xo��H�rw��?v0?XX=+ǿl�s�,q�ZI��N�><ٞ��Ͼ_�$���L�W�o��=����T4��ƫ�ء_�6��t	���ܮ��Җ��\k�e�>���=��=g��=���<3�����<�*Z=�x<��.=��@�2��<g?4��K[9�P���i�@W?<�n1={�g�+Rľ��v?\�J?��(?��C?ؙ�>��*>�����o�>�w��e?ADV>t�C�V�ľcA�U�i1���'ξF�Ͼ�KZ�2��I>�$M�TA>f6>�6�= ��<a*�=�]�=�'�=,$����+=fȲ=eb�=d��=^�=��>Q>�0w?"���>���$7Q�5�罨�:?�6�>�U�=oƾ�!@?��>>2��f���e�0?l��?"Q�?��?-ri��k�>[������}�=��cC2>i��=��2����>��J>�{��I��u����3�?@�@ǝ??ߋ��Ͽ�_/>��Z>�T*>�S�Җ6��l�D+4���j�y7?��5�~Mξ�sr>�i�=�u;��.���$�E>.��=rb��WW�w�=�^�~�P=mf=��> K>�N�=fv��"&�==M��=V6/>�4$�r���������</WR=�}^>QA>��>�Z?�Z6?�~?���>�뉾Q���u�����=t��=��>�o����>�g�>��?�B)?pF=?!9�>|K����>a>��)�Y�Z���ؾy�F�1:q>��?/�h?���>4�m<����h�4�դK������?�zE?W�?�k�>|��>�W��L�#��P,<j�=��>k2�������M"u�j�`�Ʉ���>�=�o�>ؘ�>*�?R�>���>�W�>�c�=e��V�V=�S�=�8t=��#�UNk>&|o=|ݛ��r��
.߽���=i ���=��>���5%�ŵu�TE�=��>v�>FG�>A��=�|��sPI>g���^A�$��=5Ѵ���=��e���{�*�(���.�V�V>�c>c4x��܏�� �>�Jd>0z > ��?�Wh?YJ>c�Y�ƾU���䵁�&�V�.N�=t*:>+���D�J�j��L��ھAu�>c�>���>t`�>5��D���M=�̾.�@���?=�����ѽ��F�h8��󢚿"�~��\��Z+,?剿?>>y�?�X?w1�?U��>x8��49�!��>Is�9A��nVȾC�����?�S?ʳ�>j���|C6��˾G8���n�>��H�%�O�u��80���������б>;����;Ѿ$03�gg���֏��dB�XTq����>G�O?���?kxa��V��5O����E���{?�f?���>}�?fb?!"��Uy�������=J�n?���?4�?��>��>�D�n�>է�>O�|?AWf?���?������>p�Ⱥ���=��X=V(��a"A��=ܷ8�>�?��2?,�?
���	~���������(�ѽ>(��==��>�s->7eK>�e�>C+>i
>��>��>>�:b>+��>��>/�������8?�>u��>�;?K�>��>iɤ��>lv�;q�5���'�pͽ`?���M�= V��C>��>�=�>�\˿���?�K>��ؾ��?�E��oּ����=aꊾ��>�i>1r>��>���>߸�=��>bZ�>��Ҿaw>�S��P!��dC���Q���ѾK?{>�����h&�Bk�c����lI��D���b�Yj������==���<P0�?����Ek��)���u?�x�>�F6?����Ȝ���>=��>	�>�����d���������O��?K��?�?c>�>��W?Р?�x1�D3��mZ���u�*+A�We�ص`��⍿������
��3����_?|�x?uA?}��<�6z>i��?G�%��ԏ���>�/�� ;��#<=�&�>����`�ȥӾ��þ�H��DF>��o?�#�?�V?�JV��jм�F�=v@?X~?��l?z0?�@?�u����?�6A>Ę?��?]�?�J�>9P�>/y>�+>'1=��=*a���^�7彉��/8 �]��<�x�=Ӽ��~�=��������Pw��ݤ:���+����7�=�=
>v"�=��>:KY?��>��>�9?*`��`0��ڥ���'?�Ym=�}��D���������=��h?I��?��X?�f>�C�m�D�s�>5��>j\>��R>'�>ф��D�X�=��>��>Sy�="=��u�����q��	g�<�{>5�>:�>�`_���">�˛�t���}>:?T��b����[�g�E��'�9a}���>�T??7�O=x\ھ%Ȑ���`���!?��??J�Q?�=�?���=�Ҿ��9���J�(O ��r�>|f<�X	����������m;��N;��c>�����e����T>����M޾]Xr�"G:��H񾺞�=߽�9�=�j�?۾,`��}�=�I�=Y'��g��ᕿl���HF?��4=�֜�2?�����F�>)"�>V�>o�ʽ,/��^�8�=G���+n=���>�r<>FM��X���F��O��d��>x�6?��c?S�~?J�G��G���"A��-��ְ��GB���?��>�?�!>>������V�Ş2�e]�>;�?����W����7s����nƽŤ�>�]�>�(?�R?���>hB]?u�?�~�>\�R>^�E�w*ֽܧ2?�p�?��>�ga�ZbվZ�����+�a��>��?/�l����>��?��?c�'?��?#F ?@�>e����7ݐ>�_�>k}�r|��Q_w>�@l?g�J>�**?#�w? �>μN�҉پ��<΂l>���;��/?^U#?�n�>�R�>��>Fϵ�S�=�k�>T�o?׌�?*�? �=&�?..L>k�>I�>&7>'�?�?P1?jr?S�P?��?��[=ҘZ�+�m=�8;Z7�<�0ֽ�E�Z�=�P������1�;�>��2��ҽ��<1h;�kH=��c�Uԋ���>��w>>���V>�'ƾ1.��kI5>��μ�y��¡e�H!*�bh=�p>��>��>Ǹ!��݈=�8�>��>��� W,?�?�?Z�t�!c��Ծ�|_��|�>�XD?F��=�h����v���=Z/r?y�^?M%\����l�b?"�^?�ﾇf=�ipȾ�Y��辟9M?vF
?�$J��>7}?��p?Ȃ�>f]i�Fl������c��(e����=���>+���(g��Ǟ>sq9?�\�>ѕ^>s��=�پ��x�����5?�Ì?'ݭ?��?I?.>_�o���޿� �����]?@�>@���}"?���V�ξ`��E�Z⾛���d{��zE��2~����%�r$����ս� �=�Y?�Vr?ip?q/_?:���c�H�^�䈀��/V��)������D��0D��B��&o����5��"Y��ѓ>=�9_���F��p�?Ww,?6����>έ���þ[nǾ�Y>�_����
�>�ҽUo�=���6�l��"�!QZ���?}M�>�I�>�8?:gW�!�I�8E�gQA��;ξm�=sK�>�>ޙ�>	��;d-�Y+�=�þ����H�_�}>v�X?��o?計?m.�<(P�ɇ�������XT�e�:��>�>�=��>g8����=��P��zi�ayO���%� ���*	���j��41?�=�>�,h>�`�?�#?k�߾���`V�>�Q�%,�ұ>�5?���>q��=ȴ�=�����>�l?���>�$�>����T!���{�%�ʽ��>�ح>��>��o>��,��\�e��j����9����=֜h?ǅ����`���>R?鎐:j*E<;��>.�u���!�p��7D(��t>+k?M�=��;>B�ž�8�c�{���p6?�= ?��v�[�:�<�K?˅�>r>gdb?g�`>P��>�$��/?=�Q?� ?y�"?�A�>�5���p1=8���JZC�.�C��iE>~�>�ؚ=yd=iRɼ��^���W�򄷽4S�>����ͦ��>�O�='��;/�����=b׿�MF��X�Ih#��|ݾ�,ݾ~P��2�����ʽ]m� þG����I��~�K�0�,HP�ZC����SI��8�?b+ @�g�̢� }���sy��
����>aI����=O���N����1���ޏ�=�޾AD)�a�M���P���A��'?0���_�ǿ����9ܾx! ?A ?3�y?7��"���8�� >�\�<'��ĝ�*���4�ο����^?���>��+/�����>���>�X>hFq>��!잾��<��?ֆ-?d��>3�r�;�ɿh���	ä<���?�@��@?9$�����r�=���>\�?>Ò�]:������>b��?]S�?��<��Z��{D��Gd?ɴ��A�q�О�=�s�=O�=��h2>/��>�սgH��yv��B>�Q�>�3���A��K�L�<�W>[�ҽ&ʄ�.Մ?�z\��f�#�/�+U���R>�T?F-�>}5�=�,?�6H�S}Ͽ�\��*a?�0�?ܦ�? �(?1ۿ��ך>��ܾv�M?�D6?���>�d&���t�l��=	7��`����I&V���=���>�>}�,�Ջ�M�O�!A��c��=A��R�̿	S4�H/+��L�=.�$>�"`��������<�<�<_���=�i,Ľ~�U�{=�*�>�D�>���>?�o>��c?L��?�>�H="B�BH���;����j��r��<���Z��ǅ��`��J��m����������ؾP:���=!U�����@"�]��F���+?��:>����7�L��7����Ⱦ,���e��W���cždD,���l�G9�?��??Օ����P��{��f̼C�ǽ�wU?=�
�������rV�=б=�n�=$��>��=S8���2��wM��^9?�C$?����n��O�=%]���=<�?��>Xg;����>�:?��9�龜aP>�r�>���>Ř\>���=�\¾\�BY8?�Y�?qG@=�ȾZ��>�X�9�z�*Z�<��>�2���\�# �=����þ�	���k>��� �Q?V�>��D�����績�a=c
��"l?n{?��>!
J?�?��=�Ǿ!b_�Q���v�=ؖD?x�C?�9>�|�LD׾�A^�6�!?{�q?oz>�ܽG��L��]վ��?�/?��
?�v��[��E���K�ǂ=?)Sv?��]��T�������V�Vĥ>��>���>��8��>�z>?�#�s��屿�Q
4��ў?�@�b�?1�)<r����=r�?V�>�DO�X�ƾ�屽MP��.�q=.��>	��'v��$ ��w,�O�8?q��?l��>�i��I�O�><��@�?�݇?�Z�Oɼ�G����H�|Dվ���d���¦���@�=|p۾k�|��d�������EV;�#^>@�@�1�e`�> 
(�%��*�忠����U��Oľ5�>$�>����5%�|�l�@���=��\e��v�j��>)�p>�M��{�ҾWdj��+���6֏>�>�B?�V��"�M��c��H:�> �?��>%T=g���Ѝ?8���Ŀ�N��#	�DRJ?��b?���?ʴ�>*���鸾��f�ך�>Z`P?�A3?͐(?������
��j?_���V`�3�4�SIE�%U>h 3?F�>
�-���|=�>g��>_h>�#/�d�ĿAض�2���f��?>��?Fn����>;��?1s+?ei�E8���X����*��\0��;A?>2>y���]�!�K/=��ϒ�'�
?�{0?@y��-��A_?P~`���q�l.�TIͽ�;�>�P2���\��4ɼ���_�e�7���^{�Q��?1��?�&�?#���!"��_#?�Ű>
��NȾ	8�<ۥ>�Ӹ>�\I>G�Q���q>����W:��	>49�?�4�?�	?�����ަ�9�
>4�}?�'�>��?�e�=]{�> �=Vd���?E���">��=��>�q�?W�M?���>\�=ܥ7�HF/��@F��=R�L�H�C����>�a?��L?��b>\c��}x/�g� ��νL�2����6�?��,��ི�4>�<>��>0�D��Ҿ%?����Nؿ5}���(�4?���>�V?�2��So�-컓�]?�4�>����/���ȋ������?G��?^-	?$uվ��μ�>�Y�>���>-�ѽ�W��p[���|;>�B?x�������%p�X��>R�?��@�f�?��h��H�>�zվ<΅���������0�Tc�=��?�&���W�>C�?�$̼P���y���ǻl����>Nj�?�&�?��>|}h?��Q���?���=�d�>��I?�?AR�`�վь>M��>� �mh��܍�4Nz?
�
@�
@hqL?OϦ�
Z࿰��ЍҾ?�߾F&�=���=�d�>VW��3�={%5=ӂ=���==|=t�G>4�@>^�>���>�I�>�^�>M<��*U!��=��j��9�C�k
��bݾ��;�B��MT�t�ʾ�⸾�Й�� 9��Zg�q���g�r���VW�����=]�B?�;D?1�~?�<?G���1>�۝��=j��g�����i>�
0?B@D?c�?�F�=O`���O]���p��x��l@���F�>��p=!�
?�c?�G�>�͑=F4P>r�N>���>�m�>Oz�<��.�P��=l=�8�>��?Ɠ>؋?>�>�!��/����Ii��^p��ս�ע?7ߝ�J��ɕ������i��=��+?A>���=�Ͽ�x���G?���N%��N%��>$�/??V?q$>)�����m�е>�9���g����=�����Gl���)��M>O?嘲>�">�Z��~��{���\��k�=X	�?�}� {��WP�U�Q��Ͼ}�>�y]>�>>�*��0����w���a�ԥ�=!�b?�?8�5�"�'�I!���
�1>C�5>>�>�,B�M��;-�>	�>$�ʽ��y���c>:7�=ʄ ?��>��=� �>��������>3��=53�=\~-?W�4?�3>V��D����k�-�h>�T?�Ǣ>{h�=@�Z�� K=+H�>u�a>�'Ǽ�*��4Ͻe��� |>��V=~꨾`0�"~k=Ќ����I>v漙SH�e����=�~?���)䈿��/e���lD?O+?g �=z�F<��"�D ���H��F�?q�@m�?��	�ݢV�>�?�@�?	��3��=}�>׫>�ξ�L��?��ŽDǢ�͔	�$)#�iS�?��?��/�Zʋ�>l�|6>�^%?��Ӿ�k�>qw�/]��%����u�.$=���>q7H?�K��
�O��>� k
?-?�Q�䪤�V�ȿ�sv����>p��?��?��m�2?���@�Zy�>��?F^Y?��i>7�۾�Z���>��@?�
R?e�>�;�F�'���?�ն?q��?�*I>�g�?Sis?���>��n���/�=m���k��d�=-�:<��>>Vｾ�E��u���'����j��j���\>X$=�i�>k�߽�M��{��=fՌ��©�l�r�5��>��r>6pN>��>(} ?��>���>��=>���Ӏ�QV��z�M?���?*����p����;���=U*b�ޛ?k�0?��:kݾ��>
[?Cu?�?Y?Ċ�>ϼ	��J��_ƺ�j��:p9<��>>b�?.?�>g곽$j>ZξpjD�Y�p>�ě>8$�;jBӾ�W��$��;`0�>�?�B�>�]�=ޱ!?C}$?��>h��>�ZK�Sُ��x>�|,�>�F�>��?��??K���R0�/��n젿�>W�HU>>�!y?;?~��>�����g��4�d��"~��O��K8u?�l?�Wƽ�?�ۆ?�j:?�ZG?0�L>~Z佟�Ѿ8�꽅�>�^"?�����=��*��L�ǵ?G�?&��>�q�a�ڽ򥂽����J?�X?&$?����>c����ӵ�<V{��4���w�;(�9
>�#>�g�-\�=00>���=�qJ�>�/�����Va�=�٘>%m�=�7�������)?��2��vo�Yl�=�l��G?�g�>�!7>۾�O1\?�}6�s�]6������zZ���?|�?�u�?R����e�\h6?���?#?�L�>�÷�i�Ծ�̾�L���e�	��zk=6��>x�C<�ϾU���U���A���G�d�(m�0��>kP�>'>?Ґ?�#:>���>�Ͱ����ن��󾍜9�3�f'<���1�� #��0y���ӽC��.p¾�旾fق>EϽ֥>C� ?�s�>ų\>w��>��-=4�z>�	F>J,�=c�>E��=�wi>vb>L��=�E�� R? V���k'�G��d6���%B?Cd?\��>��k�5�����M?H�?>�?�v>�sh��*�%?5��>���+
?��:=;����<>�����j��Er����>ܸؽ[�9���L��f�'?
?W?S���; ׽�����<r=�T�?=�)?')��R�=�n��V��uS��*���d�򛢾��#���p�w��Z���̃���'���"=�u*?|��?/��W�|��s�i���<��[b>�C�>�7�>�Q�>�N>,�	���1��s]���&�Yŀ����>t�{?�b�>�1H?�k;?��P?��L?蠌>�ک>���ĳ�>�r2<�>h��>��8?f�-?�<.?3?\�(?e|^>p�+6��pVھ<�?E�?WM?��?y�?zA��%�ν��h�eۻ�gk���}�Jy=��<y����u�*��=V�T>��?�$9���@x�V��>�o,?;�?���>O"|��(~����B��>���>�'�>��ھ�ɂ�ܾ���>�?T�̻��<��I>$��=6�8��9�u4�=�����<zS��}"��H�<�K�=�ۥ<� ���e�6�G�1UȻ[�=�'�>	}?���>��>s�������ȇ�`"�=��V>c<R>�>�վA�����c�g��Py>ސ?G�?%\=���=�[�=o���SX��wp��m�����<>�?�##?s�T?��?�)<?��"?qm>��<O��J��ֹ����?��*?�>3��FWN��^���\����>P84?�l�!]���_��́�gR�>B��:H�J\���B����A4 �� &=��?�à?Y�|>�,��>S�X���:��;E?�qz>��>��?W.��T�s4��n>Rs�>I�L?I��>އf?Y2�?��4?ˮ*>�S_��F�������F��s >Bo?L�M?5f�?"*�?<ND?A���[y�����^���ؼ?���j����=Da=ԣh>�D�>�<�>��l��C �����;F��=h�=��>5	>�ҵ>�H�>*ٟ=��(?���>Cw�L!�対���1@<�!+>?$��?4`?�䂽u�0�"�o�7���>�F�?�!�?w)? �� XQ>/������_�O�qN�>�>�U>�=�=��$���=g8�>�ڿ>Ef����2"�@M�+A?�?y�d���ǿ�cu�|��'���%i</⊾_T����O�K�탟=�I�����uǪ�d�_���Z�����,���nZ�q ?�.�=���=E�=�Y�<�����<�%"=�f
<�.�<�0f��g�<1H�(�E<��p��5$�b}=�x=��� {ʾ�M|?�H?M�*?��D?�5{>	�>�dL�0�>���S]?X�W>��]��̼��@��H���*��U�־!C־��a�|I��R�>�jG�5k>jP8>��=�[<��=��{=���={Y����=��=���=��=���=��>7�>`�v?~`��Y����OQ�r7�3h:?3�>�ʫ=�ažڙ@?)>>C@������Gq��1??��?S�?��?�j��>��Oۑ�(��=U	���C2>Q>�=�1�!O�>��I>ͨ�&�����q'�?*j@u??7�b�ϿhL.>�Qz>d�=��p��*��ۧ��~�����82?�K�Ǌо�x8>��=�ࢾ��¾eX��} >p��=��n��S���=}O��9��=H}�=I~M>�d�=ς�=�DJ=,�꽉��<�(�=�o>�Y���;��l�D�d͞=Q�==�(�=�&>�I�>n�?b�4?E i?�̺>���W�Ⱦ�̦���c>��4=�m�>T��<1cK>S(�>mf2??5?�yA?��>�"=c��>⤠>%L,��l���Ɍ��q�=��?Zw�?���>m��;'G�lb�`A��hؽlw?(�9?� ?wL�>�����5�y"1�$rK<b�=��>�^������7��8ʶ<��'>+��=6�$>�>���>�j�> �?���> �>S��=�!*��|�=B
>c�=��uM�=��B<���=6��������==�q߽i�&>��x>�ʾ�ة��Խ���=�<�>@>���>6G�=���z\>�~��׷?���=��]�9��e��v��M(�f�p���X>�=p>�/T�%�����>p�p>�h'>���?��[?��6>Z�_�`������������!���=�6>>ѝҽ��8�8[y��?J�����#�>(~�>'˥>Lw>i�(���=���=V[ྡྷ�2�^��>�i���6������o�e���ß�V5f�[~;t�B?�v���L�=?}?�vF?�ɏ??
�>"݃��7ξ��F>�f��aZ�;��f�z�Ho�M?;�$?�0�>���L}=���׾�G�;-�>$T���-M� ����+����YmR�[�>�D��P���أ.�cPx��\��e9�2Yq�H��>qK? Ҭ?����s���<�ב�Q?ֽ-� ?��G?�K�>{q?�?����:�O��'�>ەs?���?���?���=6Q�=�A'�'��>=	�>��?9��?��|?���`�q>����:��c=Z�l����<����������>S?*�?$��s1�gN��r}Ӿ��f��>��>�K�>}�	>%p>���=��=k)c>n�%>pX�>1N�>��>7#�>cJ�>�*���
��@$?�>���>�1?z�>1>�-�b�=���Y�$���ͣ�Z׌�8O��Y�)��0�=�Z�M��>^�ƿTؐ?�2;>jQ��/[?�-󾫙�+�2>�kY>͕ʽsT�>J�d>��*>:��>m�r>w>�6�>��>��Ѿ]�>JN��� ���B�6Q���ѾK8|>9ě��=%�Wd��S���2F��೾S���@i�����n�<�m;�<�
�?v��.k���(�	����=	?M�>�G6?J�}���K>�	�>�D�>�|���B���ލ���ྐྵb�?���?l+c> �>��W?Α?�1�m3��oZ���u��A���d���`��፿����͛
�����T�_??�x?zA?�ۑ<QDz>��?��%�fϏ�3(�>�/��;��<=`'�>l��� a�S�Ӿ��þl>��iF>�o?A%�?lT?�yV��Db���>��9?Q'/?"�u?��0?{/>?2�}#?�/>i�?�?�22?b.?�
?g�>(��=���9	f=�U���܉�3�½�ý�Z�N=���=/�-�9;k =|�<�\ͼ�������A�����9<�Q=An�=h��=ׂ�>�X?�8�>���>~~5?�`�3�.�sO��W)?��=e���f���������M�=Z�h?F;�?�HY?�2O>B�C�c�A�n&>|݈>Fe">�T>�>���F8K� �=|�>�>�)�=o"*�l�y�H	�@���';=)�>L�>r�a>`8�(�G>z]/��C����>w�������{�/W�ƫ�r��s΅>GM/?
�?��q<+��ˇ��jmP���?��,?C�5?hɋ?O�C>�,����b��5A�K��Z��>�|U>�຾�蓿)D��{�.�t>��q>�b��h�h�sO�>0�n� ���j��(�ھ�n2=������c=����߾Ez�gް=᫑=^���������U���4??2��<����*
��!��w�	>�0�>���>X�a��ɽ�rR��䷾	�Z=鐛>� 5>��}��f�B-@�GV�h��>�V9?��a?!�?M�
����Q�)�$ξ������ݽ�n?܆�>��>e��<�n>4�Ǿ��E��r�<��>}m?�u9�Ei����
оiW$���λ�?A;�>�b�>�1�?�v(?&FQ?q>?N�?4�9>�h�T6?S�?��6=4�`������g=/�`�>�?A��!1�>�&?}�?�1 ?4 -?{�>R�#=��s��j��>C+�>�3v�\Ϳ�)>���?'�q>Z�?E�~?�M�>)<<�V	���v�>�m �h��>@�,?��>s�>���>{�����=�[�>�$p?;�b?u|?�t��?��N>X?7ʖ>�nt>���>*�>W�2?��}?o|L?24'?�h�;P3����6�("�;.��=��$�i��=ڡ
>>�=����9.���ݼ��; $=1R��8Ͱ�5�D<�>BU�<�n�>�4t>���p�0>�ľ�>��R�@>?����P���ʊ��d:�/�="V�>�?7��>�o#�Q�=�s�>��>����(?��?�?��+;�sb�Jyھ�TK����>��A?�y�=��l�$z����u�X�g=��m?�u^?�	W����Z�b?�F^?���f�=�k�ľ1Q^��1�:�N?˩
?XXD�Vݲ>�~?yFq?w��>:%h���m������Hb���h�;�=l�>ݯ�_�d���>p�7?�s�>�Ib>K��=�۾Cx�G4��|y?3^�?a�?j�?��)>'�m���6�Ծ�R��|fS?���>�ĸ��!?d�;��ҾU������&�ܾiա������-��x)���8O��؆�S��\��=��?~�_?g�?:Va?��C�d���W��t�=�J�\*�F��I�=���R�F�=�ʷl���Z��������=S�I���<����?.?�@����>��
��>p���+�>�S��z�C�Ŧ�=�s���2A>�~�=A|�y�&a��o(?�Δ>��>:�7?vqi�4^L��[D��3 �ѩ��۽=�,e>�>.�>0؛;$�F��F�|қ�������2�z}>��\?~JN?j��?y�N=�.?���~�2?
�ġ��q�Z��>�>��y>=�.�$�3=޸���C�N�g�/����� ����<J3?$�j>{�>w;�?٣'?1���F�����% R�<W;��TK>B�B?D5�>���>�������Y��>d�l?�U�>;�>ꌾ�!�̳{�A8ʽI��>�C�>:B�>�Mo>�a-��C\�X���u��~9�;��=��h?���
La�^��>R?}S�:�1><-p�>�ut�!�ͥ�
�(��4>��?��=?;>��ž`��W{�nꉾ+?y?W4����/�F�m>D%?`��>���>؂?Ϣ>��þOѻl?�W`?G�B?�y<?��>�$�<�D���T½�%��V�<]�>�oX>��y=�J�=e��X��m#����<�2�=����н�}�;W?��%�%<�R=��>7�̿]4<������W���X���r�j��
�{����q>;�������[ʖ��
	� �e=rZý̒V��9:��<����?�@�Il�����u����gv�y["�2��>��X�]�\���R���o��������֞�ƻѾ�9��Zm��v�R�'?�����ǿﰡ��:ܾ7! ?�A ?2�y?��3�"���8�� >2C�<�-����뾬����οE�����^?���>��h/��w��>ڥ�>��X>�Hq>����螾�0�<��?5�-?��>ǎr�.�ɿa���¤<���?/�@��A?��'���쾏H=�y�>��	?�?>�2���௾*��>�מ?��?iRP=t�W��'���d?7��;A�F�PۻzX�=p��=�>=�^���J>e��>�<��/A���޽ZQ1>��>w%�7D�D�]���<��\>�wԽ=���5Մ?,{\��f���/��T��U>��T? +�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?:ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=s6����{���&V�|��=[��>d�>Â,������O��I��T��=��g�Ͽh]�F!���=�wh=��]>��'=�$о�T>G㺾t�Q��Ƒ�f%�:[J@>Q��>�q�>`2?(��>�J?�g?:#>ȓ�=à󽵵�Ώ��3��Ny�=��������w��l����Ձ���V�ǽ־���<�	�
(����-��
>�_�Eu���T1�tgQ�\|B��a?��>�;}��+��k��(�پF���q���(=�������n���?v�S?0c���V�?�����_��ǫ[?ԯM��
��0f��Ϙ��L�=���(m>���=Μ����0�	Y��4?=p?��þ�̆����=t^���0= a!?���>&)�<�?�>]i?w�/�)�,H>Ry>F�>b��>��	>93�����,?�wZ?c �!賾�G�>:������鋼ɫ?>��I�ǽe�F>+ϐ<eu��W����k��4�=�pG?�P�>w�7��4�����o��=v�5���?�v?I�d>�8_?/|?}��=h��\��)��R�>)?��Z?�C>�zҽMM���yn�/5?LnN?��K>W/;�j��*��"��8�>?>E?{$?DŶ;�F]��7��7�+���R?��v?s^�xs�����L�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���xY4�%Þ?��@���?l�;<��[��=�;?j\�>�O��>ƾ�z������L�q=�"�>���}ev����R,�d�8?ݠ�?���>������?�>���׮?�	�?�����}�n'��	:�4�	�P�H���G;����8�=O���Z%�J������j� ��Ī�1�P>��@)�={��>ٝ�<A�ῤmпU�����ž"<ھZ ?�{	??g4=�����֗�{�i��-��Q5������ݣ>�L>K7��猒���{��(;�ir���Z�>~ �W��>�P�*ϴ�n���#�$<���>���>���>c���������?x�����Ϳ�ݞ����xGY?I��?P��?7k?��D<b�v�Z�|�ǒ��VG?U�q?�Y?���``��j2�y�j?nX��uP`�b�4�BIE�TU>� 3?E8�>��-�\�|=�>���>�N>	)/�^�Ŀ"ٶ�|������?���? q�V��>��?�t+?�e��6���Z����*�t!$�"-A?^2>ي��X�!�-=�qՒ���
?At0?3m�m'�[�_?$�a�N�p���-���ƽ�ۡ>�0��e\��M�����Xe����@y����?G^�?h�?ٵ�� #�j6%? �>d����8Ǿ-�<���>�(�>*N>#H_���u>����:��h	>���?�~�?Pj?��������U>�}?0�>z�?�B�=�\�>���=8鰾)}+�.T#>���=��>�:�?y�M?h5�>�0�=��8�l/�rXF�}DR�$���C���>l�a?��L?�lb>����1�!��Kͽlx1�2��W)@�.<-�"��)5>��=>�>%�D��Ҿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>B�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Ua~����7�m��=��7?�0�'�z>���>��=�nv�޻��V�s����>�B�?�{�?��>!�l?��o�Q�B�|�1=6M�>͜k?�s?Ro���b�B>��?!������L��f?�
@~u@`�^?(�&ۿ�@��n�žо������<ߔ�>.�<f��=4J�<�}�=��=��3�vx�>:׵>�%�>�g�>�>C'�>�:��2�"��.���슿�L���������̽2a���28���
�鐺�����������-
5��ߍ�gݽ5s&����=��N?��A?��o?g�
?�Q��g>��ɾ�t= 	ν���<��">�!?��D?�;?�>�=�c����R��s|�kY�����w�>�2>:� ?c�?���>A�7=^��>�ׁ>~bw>�Y6>E��<�
�<)^A=�)M>bA�>��>og�>��A>Z�>S ���r��c	h�q.q����O��?g����J�U��b���}���wc�=e)?>Sd��X�ϿƩ���F?�������7#�N�=��(?6�Y?i�>`R��v,i�5z>^F��Gr��>�> ��f�ʼ/�X�E>�?ۡ�>�!�>a�9�gr9���W�eb��u�F>��%?;]�B���㚿L�V�@�������=��ʽ"�ON���|���@��=��m6A?N
5?#�7��R�^Eo�;�l�8A�;�4>�EB>i�="ql=n����<*
o����C��=�D>*�?�=->4�=��>�ᚾ�/�+q�>"�$>��)>p;?gm ?���ղ�h)��W�0�,&D>Y"�>���>a6>|�O���=��>B�\>�������G����@<���7>�4��
BE��_1��	=�������=���=�.���<��N�=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ"i�>!u�BZ�������u���#=���>�7H?�U���O�&>��v
?�?�\򾺩��V�ȿ�{v����>%�?[��?��m��A��z@�s��>V��?gY?�li>g۾�]Z���>H�@?BR?��>%:���'���?~޶?���?�M>ͫ�?\=}?z��>۷.���8�l��[쌿��<�����>@�A>�ᒾ,oB��X��J�����^��+#��S>��
=���>�۽(�ƾ���=�Nr�乾}����>�j�>�n>f��>�?(Q�>~�>5�<w�I�l<�����L?ޏ?�Y�1�p�S0�<���=�&\�l� ?�_3?+�Ȼ�Ҿ9�>�9Z?�S�?��V?��>�������Cо�����s�t<�E>Co�>�a�>wA��e�R>r2Ͼ=CC���>�ƌ>�t��|Nھ���^�����>Ӛ?���>o�~=�w!?�#$?��i>��>c@F��A��ǁC��Ͻ>m$�>Y%?�U?M�?����2�
���3$����[�@tG>,�x?��?=�>���ĭ��P����Ѳ������}?igj??�ƽ*�?��?X??��C?��J>����_Ͼ"|ӽ�%�>�g,?��3=F�G�4^K�;d��ڱ?ag�>]�>��<?Ϧ��7�0�*�ž'?m�?�?a��i�B����E{=����9c�ʑ�=a�4��c�;�&�>t�>=�a�;��;��R��s���Vs��-�o0�=�y\>�>��+G������=,?ܞG�-ۃ��=��r��vD�%�>�EL>���6�^?�l=���{�S���x��N	U����?۟�?Bj�?��ŝh�#=?��?�	?�!�>zL��r}޾����Nw���x�{v���>��>��l��'���ޙ���E�� �Ž�z<ݍ�>�=�>Mt4?V��>�R�>(	�>�O��¾�@�K6&��n���I��Z?�L�#���n��:z�\-�������̾ �F��a�>�t�l?�	?��>\K>�?/=�>��>�N>��>�>λ_>��=J�>.й>���<�SR?Z�����'��龗̰�AB?vVd?��>�ch��p�����kh?�u�?�n�?��u>@lh�g+�<L?��>P��#\
?R9=1*��I�<�A��?H�4����-�j�>ݮؽ:��M��g�ba
?T?��\̾A	ٽ2p��S5o=wJ�?��(?�)���Q�n�o�W�W��S�uU��1h��c��k�$��p�揿_��s"��(���*=�}*?�?�t�؀�|���"k��?�:If>��>]��>�ƾ>WyI>��	���1�T�]�\S'��ȃ��T�>�Q{?�>�?H?�9?7P?��Q?�S�>\��>eM��>m��<�)�>zH�>��4?U/?p�+?�w?P�%?Q�]>QC��h���ؾ)J?j?j5 ?� ?��?x��!�����Ɩ���i�&䄽��=���<,>ӽ�Q�3bJ=U.d>9Y%?�n���7�(��g�>�UH?�(�>��>�>g�����,�;{Ҵ>� ?)�>�&��Cj�ni����>�'�?���=�p=�m8=u����	=�e�=X��"Ό=�����N���{h=��1=���K'�@IC�~�_=ԏ�����>�?�|�>�Z�>/�}�s���
���={�o>qG>hT>!ݾ����� ���f��M>��?%l�?�+�=<*�=8��=�����o��8��Ӿ��W�<�+�>�#?�1]?�[�?R�@?��%?*$>��������䂿@����w?R$?ht�>&N��폕��=����i���>:)?n2N���w�����6�q@:���>��5�KBI�V�Ŀ<�U�cO��e����P���?�I�?�E=�A1��kC�k��������z??���>�0�>�?�>n�&������;��]�>?��?Jt�>�[?r�?�??��>�4W��ǿ |�����-ߖ���O?�>�?y�?��?��?�p>�(�*��j�C�T�8nͽ�W��+�@>3Xs>y�.>�d�>|��>��T=�j��z>P�h�w!H�,�D>��E?w�>f�>�[�>�?�=�O1?U��>?���-�����C���[�t�`?�R�?m�?M��=э+��U�C��k�~>ʠ�?<G�?��?4<��_�A>�`� <����V����>���>�X�=��>"���g��rg�>��>#��<���W�>�L��t?�Y?x�L>�ſKOu���|��#��aw�<N揾�qV�ݟ�z�t����=�ә�2������`�A͗�@�������͒�U�}�4 ?���=���==8�=��<]⩼�=�<�M(=���<w�=�~�y<��7��A��g�"<A�<��M=A����¾$�x?�I?��2?��J?�\>3 &>L�J���>�]��?�}8>�H	��#�����z"���tӾӐӾG�Y�>��� >�/_�a�=�1->71�=��U<��=�{�=�M(=C7<��=1έ=
��=��=B��=��>��$>�5w?e���粝�@5Q�0_�ʶ:?�3�>���=�~ƾ�@?��>>�2������)b��+?	��?T�?:�?�mi�be�>W��2ގ�lw�=�����92>���=3�2�:��>��J>S���J��q���84�?�@�??�⋿ȢϿ�e/>
2<>�>4S��o2�P
`�YPX�_\��8!?9��
˾�r�>$��=��ݾ?kȾTa=��3>�~h=c���Y\��<�=Nꄽ��>=�R�=�<�>�%C>U�=����?�==A=]V�=��L>~���*cB��%��+=�C�=�[>�/(>?Y�>��??�2?�r?I�>#o���ľ�r��D8<>�%�<�5�>�z=3}>�k�>�C?�5?�9?�>��=+�>�i�>$�B�\�g��w����>rR�?\�s?��>��i�����,�^F��)����>�/?�y?v9�>Vk�xE��RE��m"�҃o�o�y�?mq>v�0=0�׾�vx>��D��;���=��>t��>���>�.?�K?'[>~O�>���=��-�r<�=B�=�e�=.�Ŏ� A�2�=1��)����=S���������=���;���=}/��R��=��>��>��>S��=H���|�/>�M��1(L��$�=�dhA��d��+�5/���;��>>�"U>��z��鑿U�?U�a>�B>���?#t?��>�_
�	�Ӿ	����h���U��e�=��>K�>�E�<�l4`�$L�Ҿ��>+��>!��>b�>�I3��&�PL�=Z^޾o�#�2�[>x���O���%ۖ��*���ힿb椿��j��I�#�9?m���z�=u=�?�G?�m�?��>/ ��7���X{>ݾ�Ž&��Y���S��!�?f��>���>��FA��G̾����ܷ>1BI�"�O�����ү0���ɷ�4��>������о�$3��g��m���-�B��Ir����>��O?+�?�4b��V��UO����+&���o?^|g?1�>�J?EA?�*���v�r���p�=��n?���?�<�?>�U#>``����?Ý�>�n?��w?�im?�g߾=Y?�>>aK�>�8�;S��������C�?��?V-?[1?4:(��z�4��!/��}�Qư�yJ�=U#�=�21<'��>'��>�=�>�x`>��6>��>l�!?i�>|�E=
܊>���������Z(?�T9>&��>!�6?1R�>���=�O�=6�>Y�ּ��8���"���=]��=[������bK�6��>�ſB��?�HH>�JB��t	?g!�m��4}�=�"t>7�ƽVd�>7�^> �8=���>�`�>E":>��=��>�/ӾM�>���i!��,C��tR�O�Ѿ�\z>Ԗ����%�����t��>=I�@_���g��j�p*��y>=����<D�?A���n�k�e�)�u�����?�U�>�6?PԌ�j鈽R�>j��>s��>�7��؏��ȍ�x\ᾼ�?���?�;c>�>��W?W�?͒1��3�qtZ���u��$A�e�̺`�s፿�����
��
��'�_?��x?*yA?U5�<�9z>���?p�%��ӏ�(�>�/�_';��=<=�,�>�%��D�`��Ӿ�þ�6�FF>��o?1%�?Y?�OV�����j:>�R5?)�1?�b�?�=.?}B?�Ve��'?��e>�D�>���>�$?iU<?�D�>
�%>��5=����"=D<���ß���ż��׽_o}�MY�=^�M<&�;� U=K��<�q=�A�<��������N=��=Á���k;�K�=a��>yc]?���>Pu�>��7?�{��8� ���]�.?�c4=#���H�����%���>jej?���?�Z?$d>BeA�u[C�]�>Y�>(,%><�[>��>���*%F����=�>��>b�=�|P��ׁ�B�	�yP��rO�<1) >��>��|>�׌���,>���?�w�HYe>�Q�4꺾)�Q�G��1��qw��2�>?J?�9?h0�=gX꾼6��]�e��^'?�O>?MM?�8?ƺ�=�پ�"9�g�H�X�%��D�>���<
������1���P:���0�-v>[]���%o�ɭ�>�#"�� �u�s��[�G����l><�߾P��=����
�<�����>��>��U	��㔿����[>?�f<MÙ����V셾���=���>��>�������L�M啾S׻��>)fe>��]"��^�T;辈G�>�6?�]?]6�?�ό�k���H���߾��ɾ@�P�F,?B#�>q�?7��=B��=����p��bJ�����>)?Y��\o�"A쾄_Ǿ�&;�����2��>M,�>���>�n?�U?�g?|.?�?G�>0���)�˾~a.?�?G1�=}V������.)��D��ܹ>Fm?5�{�.z�>��?C?�E1?ǣC?(�>�X>Ő����>�><ǐ>�h��rɿ���<��|?��>�?�`?��>F:5��Wپv �Y��>��O=��?��>*?	L�>b��>^o��[>���>G]?u$u?hӀ?dd�<�� ?�[�>��?ݔl>tF�>] �>M?~�h?3I{?��S?���>Rw˼o���Gm$�u��~��<D�;�O���=�CY���ｉ������=��<~6M��.�=�F���<M�e�X���>�O�>gj|>�����>�sȾqV~�r�D>ĥ�{����(��{[9����=-�z>�?�͔>P�4�1{�=G:�>��>�=��&?Z�?#?ٳ�;�g^�Z�Ͼ��;���>�??���=��j�� ���Ky�ڎ�=]�i?u`?�nV�Y:����b?2^?���i>��ž?O\�6����M?�P	?$�B���>�}}?_�p?Fo�>O�e���n������+a�$�g��>�=�'�>Q��d���>�7?�t�>xd>��=\n۾u�w�tD��Ss?<��?�z�?d�?��+>%2m��]��v���F���^?���>�4��p�"?	�����Ͼ'9�������������@���T��i�$�h�׽��= �?�s?NYq?W�_?�� �Kd�\2^� ���lV��/�2�N�E�yE���C��n�n[��>��E����G=D=���8�ê?��.?��3�=��>T��Cݙ�3���ZXL>l���+n<�4)>����'�b>��2>[:��$�j�6c��T!?Q��>���>�bI?��K��)R��E��l"�����u��%�>X=�>��?�/=�L�Q0B�_���������"2x>��a?�gN?��q?[ͽ�4�p!������������_>c> ��>��S�����\� ���?���l��*�Ǝ�����3t=@�3?��>@
�>΃�?�M
?�	�����3�[��j7�-�˼��>�a?��>�e>{Ჽ�r�3��>Z�l?��>⟡>�ċ�[!�t�{�NyȽ��>��>�F�>p�m>AJ-��	\�O\��9i����8�g��=Ԟh?����$`��Y�>��Q?V�Ź��7<a+�>�)v�"{!��[�a�(�[
>Tf?]��=�<>Ež�����{��鉾K�(?��?7Z��˿)���>�9"?ȷ�>��>U�?R�>X�þb����?Nl^?e�I?A?�7�>��=���9�Ƚ�g'�D	%=x��>��Z>U�n=ǿ=����Z�x� ���N=<w�=�Aüv2��?�&<$���m�<�a�<r5>ʩӿiz@���ξ�s���޾8�������-���ܶ^����-���"����x��#�M�E�pi�7�^�b��m�Q���?'D @�V��
��/1���&r������>F轆ݬ<�)���Խ,�+�sX���됾^��1<��oT�b~l�t�'?������ǿ�����;ܾs! ?iA ?=�y?��G�"�'�8�O� >�>�<U��Z�뾡�����οt���m�^?H��>5�|3��(��>��>��X>�Iq>q���螾,5�<V�?f�-?���>2�r���ɿY���I��<���?��@��F?�#��q����=`��>B�?Z��>ˡo��,�g��컿>9>�?�T?�IN�o�r��j�(]j?���_�-��@ͽn�<�j>5�:>v��<��.>��y>6��$���W�H�>���>�6���xq�����,��;�Zg>T$!�QBS=5Մ?,{\��f���/��T��U>��T? +�>U:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?#�(?:ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�م�=h6Ἢ���}���&V�~��=]��>b�>,������O��I��V��=�~����Ŀ��3�6�����<[@#;~N�rߍ�֟?<�G�+7Ͼ(�z�ڨ������<������=<!�>s�>3�>tU?M��?}�>��G=��佚Hg�/�ľ�z���M���۽��"�ζ���$����t�������5.���^¾�(�~F%>�`�'7��]1�q_J�?�?�	>?d	�>҉���8�=9F�eɾ��ʾ�(k��qJ=��f�Æ����i��I�?�tK?�Η���@���8���;E�-��?<?���=����g���f=�>�&f<Ɍ�>�\>!�T�D�,��S���1?(�?�����>���j#>�y�~�E=��)?���>_��;��>�#?� 0�����Y>.� >;Ũ>4�>���=������㽭�?��W?�4ݽ���y�>E����{���=�>/��T5���HM>O����Ă�nT#�������<�+H?�ɮ>�J���/�JT �Ӫ$>!�ʽyQX?I?s��>_W?���>��	=�+Ǿ3�D�����a>%s1?��J?�\2>�����xľJS��!C,?��k?O�>�FU��M����T�9��>�W5?�[7?���<^��+���g/�JB?s�v?�q^��r��#��M�V�>�>�\�>+��>{�9��k�>F�>?�	#�CG������^Y4��?Z�@"��?��;<x����=�:?=Z�>�O��=ƾWv������՟q=r#�>�����dv�����N,��8? ��?Γ�>����o���>�^�����?�e�?�zo��"��%P�X�."�%z�=	�0�H`>񻬾��IľE�4�<B���i<.}p>�#@�wٽu�>2ת�l�ܿ�:׿ۓ�!o�s6C���!?i��>��< �=� �x��m��?���:�ng˾Lg�>K�&>�Ὦ���j~���4���!��	�>�c=W(�>�O�q��%ɝ��M��ܝ�>���>��>�\7�����D�?2�羑�οV���b�v_X?�/�?L(�?�!?�4<s�y�㡅�K[�<��A?]�k?#�Q?��{��og�$n���j?\C���B`��p4��'E�+6U>�3?)�>��-���z=gL>L��>>l@/���ĿiԶ������?:��?>|�B��>'��?�o+?�R�r)���O����*��@X��;A?b2>���:�!��=�h咾��
?Ym0?��k���_?h�a�=�p�D�-��ƽ�١>��0��T\����'��iWe�����4y���?(]�?��?��#�E6%?��>����-Ǿ��<w�>;�>�N>6)_���u>S���:��j	>��?�z�?�g?��������KL>9�}?C%�>��?���=�a�>r�=7����V.��S#>\��=��>�}�?��M?�T�>5r�=�8��/��]F�xGR��%���C��>��a?r|L?OPb>6���#2�!�4xͽ�O1�`��%M@��,�g�߽.5>j�=>H%>��D��Ӿ��?-p�+�ؿ
j��wp'��54?*��>��?#��(�t�����;_?7z�>�6��+���%���B�V��?�G�?4�?��׾S̼�>8�>�I�>C�Խ���t�����7>�B?V��D����o��>���?�@�ծ?�i��	?'��P���`~�Ƃ�` 7����=��7?U/���z>���>&�=�nv�ʻ��r�s����>�B�?l{�?���>�l?��o�z�B���1=gK�>>�k?�s?J%o���8�B>7�?��C���UK� f?��
@Fu@e�^?*W�տ�ࢿ?���~������=��=)�>�핽�=`ɵ���y����=cL�=O�>���=��&>o�:>D҃>Lk�>Ȋ��7k$�8S�������cD��� �_���4��X�� (���Q,��އ�Nެ���8<|����S�_ڽ���*��ˁ�=�HB?@rN?[�g?���>3��' �>Z�ǾG;k A=�{�4e>��?A�F?�\'?�[<�,��3�Z��Dz�����
5�>B5>�	?7?��><p弫u�>��>�g>Fy&>���<�p�}�1=�'�>��>n+?�i�>�Bf>�7>bֺ�ԡ��!o�^7��lE��ҫ?�5��
M�V��w@ؾG�Ѿ��$>��?��>�P���_ֿ���9?*������$����=mX�>9Y\?{RQ>d˾���q=8�����9;>?j3���XM��5>T��>���>fL�>�7E�D�>�C�\�^]��$�>>�G?�6����~����g�[�7,���>Cۧ>8L7���(&����}��84���ؼ�<0?��0?���|������R	>���;�[?=�}P>�U>|E��,�l��&2�"Fռ��H=-e=��?�x->rE�='d�>� d<�#ׯ>o]<>�->��@?�*#?qN��
ə������T�xy>���>�h�>��>ωD��7�=<j�>�	^>Kh��$��A���0���R>~ꚽ��f��m���x=%���{�>	ք=���"@�?�M=�~?���$䈿��ke���lD?K+?���=X�F<��"�< ���H��=�?q�@
m�?��	�ݢV�:�?�@�?��R��=�|�>�֫>�ξ�L��?��Ž@Ǣ�Ɣ	�9)#�aS�?��?��/�Uʋ�>l�u6> _%?�Ӿ�
�>�;����z5��@�u�8�-=�ɿ>R'G?�Z���C��<�{
?
�?���_Y����ȿ{0v�h��>��?e��?mOm�(:����@�xQ�>���?xY?D�f>7�۾iY���>e�??Z<Q?sG�>�,� �)�r/?S�?j(�?[I>�m�?)�s?��>9r��n/���sp��D{=��=;�ؐ>��>�4��4!F�cʓ��B����j����N�a>�%=,l�>u�Y����=�1��-P��:�k���>s�q>0�I>�>�� ?f��>_��>�3=˝��J�������_L?0��?���nn�g��<�M�=�]���?��3?@VR���Ͼ�{�>�r\?���?��Z?�v�>ӳ�m��n˿�W���d�<�tK>�/�>u^�>�.���aL>�@Ծ}�D��>%�>⣡�}ھ ��:#��L��>؏!?J�>�O�=H� ?H=#?n>X�>��B�ፑ�_�D�C��>��>�f?�b?Z?��_3��r���!��3�Z��WO>9>y?�?睖>�-���g���/����R��җ�y)�?�e?x۽�D??̉?�5??�??Jk>�k��վ�p��1$�>�3-?�R�<��=�M@Q�-��!Q6?�� ?�x�>2�/���];x5�(�%�c��R��>ZeI?�$�>J�Ѿ��I�M
���o=�t�E8b�� �=�u=��>F��>_�=�U�=b�=�N
���V�X�[�t�$���	>��[>�n">t:]��R��;,?kG��惾͘=�r��qD�=�>EL><�����^?�e=���{�o��tx���U����?���?�i�?�&����h��=?��?j?��>�<���~޾��ྴew�	}x�Bq�'�>���>X�k���������H��!�Ž�1B�q��>`��>�H+?WK?zaL>���>㼋��J.������Ƈ�7H�� �ɡ:���R�X�#���W�3<½s�=.2����o�?��>���壒>??�;�>�?>���>S>	�^>�8>��
>�&�>��2>ٗ\>i�J>Rn>C�A�)ZS?
��E%�qg������+�F?�x_?���>򰫽��}�X� �g�?F}�?�E�?>l>6m�Z�)��?w��>y��v?�=��
��<� ���OԽ�E+��a��!�>e��CT6�MH�����a�	?�R?E�;?�������e���Bo=�N�?�)?��)�s�Q���o�֊W��S�4`��Qg�������$�/�p�fꏿ'X�����\|(�#e+=�*?��?"��=��
,���k���>�Zaf>��>�)�>E��>/|I>��	��1�v�]�;'�,���4�>6W{?V.�>�B?�e=?�&G?�!L?�В>2o�>H#��5F�>��=��>�\ ?��.?{t?(u,?��?~0?P�z>�N��@���u�׾+3?�K? �!?��?J$�>al��?���s{��|��ʆ�����L�=�.�<
�9��	��\,=�l�>��"?��Y���/�&��bJ�=��J?m�>���>BाZ�����<���>.��>��>�꾣���+��f��>��}?�DӼaI�<���=g�$=;����$=�c4>�����{=�4T�w)˽��ax�=�	�ђi:��y���<i�=�/��)�>�
?��e>�;}>?���6\��v^�?\�=��>̯K>��>M�ᾹL������Oe����>���?��?C=M�>���=ע������k�
�O���,<�?�?��M?�ɐ?�2?@�"?!z	>e�J���0�� �G?��&?J��>�0�?Z��z���g����>nq'?��`���`��g-�k�����D�ӂ>��"��*Y�ڰ���\����� �����L�?�W�?�>��"���\��{���v��+vp?�ʛ>���>�?#���/�%0��[�>�w�>L>?�Q�>�V?ʴ�?|�T?Q&?_W�ڹ��eB��ԓ����j=�?b?,Ё?�L�?�Xr?�3F?H?�>?���^m ���8�t+E�S��I9ֽ�">ȵN>�dZ>^i�>�*�>^�z=�g��í�=�u��[�MY�;�Z�>��>媭>wK�>��0>��@?���>��޾T��t�ƾ$Zv�b��eRi?�ƙ?��&?���<�`�M�;����Ĵ>�#�?��?��.?�~��r>�G�k�ľ�O`�p֚>D2�>��><Z�=�8D<4~>��>'"�>��ݽݝ
��,4��c��6�
?W;+?\��=�ƿI�q��q�����5f<�钾[�d�����V�Z��;�=����Ж��Щ�+�[�Nˠ��r��ִ���9���{�d��>��=�K�=_��=_�<�ɼ�D�<��K=��< �=>�o��?h<,�9�ӌܻሽ,���W[<#�I=ŋ��^�ʾL�|?�dI?��+?�	D?~�z>�9>'N*�?�>cdm��;?�S>��U�4㻾)�;�r���Q���;�׾�־]Ld�g8���>Y�I�j~>�4>Y�=,bu<(x�=�Aq=t��=h
��<=(��=� �=ޒ�=���=�>)C>�5w?b���x��� 5Q��l��:?�5�>c|�=O|ƾ�@?x�>>�2�������b�,?���?�T�?�? wi�Be�>r���㎽�r�=9����C2>���=0�2����> �J>'��?K��=���t4�?�@;�??�ዿ>�Ͽ�f/>ߜC>)f>�Q���4�Pne���C�5nG���?/�;��ž��w>���=��߾=�ɾ҆S=�>�ć=���&�[�)C�=	󈽡�=���=(�>�h>>�M�=	���6��=p�$=��=V[L>q���4�o�|�"��.=-��=��U>5>
;�>5�?��9?�s?��>p���6
ȾDB����F>ۅ�<l��>���:��9>s��>�:.?]�4?� 4?�>_�=ݯ�>�_�>��)�%�[�l4Ͼs���m �=Zc�?`�?$1�>�l�:s�����/��J4�8�N�C��>A~4?��?s��>]e	�fn�N �4��?7ʽ��P�$/>\�<?A�=��8@׾+b�=TG=���>>�(�>o1�>���>�R�>��>�V�=2�ͽ��P=t<�;�,=�[꽻�=~�$=n�=x85�!����G�V���n<������?<rnR���#��[�=��>`>��>��=�D��}D0>�ϖ�d�L�
�=����hA��"d��~��b/�X�6�SD>�V>+脽X!���_?}[>QMA>4{�?8�t?�	>��;־]*���b��FQ����=�T>�{?��.;���_��mM�\Ѿ��>o��>��>�ф>�`"�l<��n�=
@ھt�=��>�>񐾢 Y�4W�L/h�B'��S��ܭ\�y�=�2�5?���+��=�(�?q�B?��?��>����A��O>��Ag=#1�?r�����?�x?�$?����5/�!�Ͼe+��j�>{�W��lL�Y���T�.��
b�
��ޱ>����9�Ѿ,�4��_��zT����=�7�n��m�>G�J?��?�-p��^[N���g1�����>|�`?��>o?�q?��{R׾��n��<�=I�q??��?���?���=�+>�@��}Y�>��?ώ�?Ǹ~?_Ӄ?��.�� �>���<Қf>�$�6/��3�ʽ9���>{�?<B"?�?&�伬�վ>LԾ��M7���?�;��=Zׯ>�:�>�0�>ϫ�=;���_�>��&>c��>*�?̴�=X�>�6+>fЛ��S���!?�	>��>��*?L��>��=W��0y�=Lw\�pO�ݬ�QP��E�����=_�����<lb�� ��>�ÿzQ�?��f>�G�1��>����<>���=�]�+=�>Ĭu>z�=>˳>l��>O�`=
r\>P;>�rѾ5y>C����!��oC��9Q���Ѿl�v>�ќ�6�!����+��e~I��������j�X���=��Q�<���?�[���k�#�*��e ��^	?T#�>��4?�P�������> ��>�w�>L���+^��O֍�H⾉8�?�?>>c>��>��W?��?}1�o3�gqZ�ƨu�X&A�e�+�`�N፿c���ҙ
��$���_?z�x?�yA?��<�@z>}��?Y�%��ԏ��>t/��%;��'<=b-�>�#��~�`�^�Ӿ��þ�D�&XF>��o?\$�?JU?�PV�Lu����>�8?�-?6�y?�I1?��F?�!߽�d.?*y�>3��>λ�>�$?
i)?��
?�D~>T��=�Σ�3n<=�f��%M���'���彝����=��ａM�7�=~ ���W><�N���b<�b�<:�O=B��=7����g=��#>�]�>�\?���>x��>��7?+���6�Z�-?��5=/~��*���W��:7���$�=�Kj?a��? �Y?�c>RnC�	QD���>�p�>��)>�5]>5�>��l2E�CЀ=��	> l>�}�=�-H��0���!��U�����<3Q#>�4?|>A�ͽ��#>�t����F�B$�>�<�����Ï�CQK���!����K�>�09?�d?�H>B���T1�i�a��A?�T:?3�\?�m�?���<`-޾\�>�$M�![�*q�>��>c��<����8��[�!�F�<�HX>7�j��ժ�s��>ΨR�wl�����c���:��}�H$Ҿ��<���Z��!c=%<�>���>��ƾA�ؤ�8п	�q?�{��ey�������>/��=���>g'ܼ�|$���%��z�����>��>Q1Y=�bT�V��'ta�<��^p>5R2?�dV?sҍ?���XWm�w�^�������(�a�σH?v��>#s|>�ݪ>dCW=�[��"���y>�����`�>*�>W��K:��	���M�tI3�yc�>��1?��j>B�?�Y?_��>7pi?u�(?I�?���>qY��͝�'?&?�ǂ?�a�=\ν�]�t9��BE�F��>�J,?�W;�R��>��?U?��$?+.O?��?�B>Ľ��Z#>����>�W�>��V�(}���9^>�lG?�d�>�&Y?s�?�^L>��8���������:~�=�s>�2?�#?�?�>Bw�>H���tP�=0��>��b?���?�n?���=��?�5>�y�>Jޚ=K¡>J�>.�?{/P?��u? �F?#��>�"�<梪�/�%�|�������;tT<��^=��	�|y��t�o��<���:FU��	~��Z��a����޸�:O|�>��s>j���P0>�ľ����@>2���#���N�:�hF�=�a�>��?�y�>�k"�픒=��>�v�>����*(?��?�	?��;��b���ھ��K���>t�A?Rf�=��l�d�����u�c i=��m?�^?1W�5[��g�b?��]?h��=�J�þp�b�\��t�O?��
?x�G�u�>��~?6�q?·�>��e�9n����/Cb���j�%Ѷ=�q�>VX���d�M@�>Ĝ7?�M�>��b>��=u۾��w��q��|?J�?��?���?�)*>��n��3�q���[D��^`^?���>q��q�"?	��� Ҿ����H.��S��T���$���7��'��<�*�.��,=ǽ D�=F�?c�o?��t?=�_?w��N�a��`�nt����T��� �Q�YC�>�C�m�A�Y|n�(]��,��ļ����J=O'_�GK�2��?�$?�0�EE�>.����
�K�辣lW>$���M���J<h<�Խ�]#�G?-�&���I�սwo��ǌ#?H^�>�k?�4C?����6�o�B��	5�מ���r>e�?貀>��>��z<����g�������[���ۼ#�^>�&I?�S?�D|?����#�����I���:���)��>C�>��s���ؼL�N�����YG�I�c��t�������;��D?$my>��?b�?j�?��"��0�J�l� .��nWm���;��/?3>b-@>�5�X�����>Ml?å�>�D�>�����"��z�?̽��>�3�>�C�>a�k>�1��-\�m;���[��͢7����=܊g?*"��#�`��U�>��S?P^�;oL<Uܣ>@W��RT!�J��a.��^ >8�?�=B+:>{ȾQ����z�����o1?��?+����t<��~�>s	%?ng�>ii�>%8�?Vc�>��yJ�=�?�G?J�*?�Z?�=�>�t>�g�=�"��q*�K:)�a�>,�`>Ӯ�=B_�=��R���z���R<�i<� 9�1����f�<S��=d��<h�>[s�=M�b�1�=�Ҿp��Mz������#1M�}�s�����ያ��^��E	F��x��U�>1�潕䛽�-���;�?!@�v��h�ƾ�Y��`6d����O�>D���D<����;$�O�H�'#�����Y>��`��a��{�q�@?����-ҿ5���_�����h?���>Q�?D�"� �J���|f�^s7>��>@���c挿ɪڿw@־|9a?�$�>h����ͼ/�>���>3�Z=��>-'+��;ƾ�4C���>zf7?�ӈ>����߿�����ʹ�BY@<��?(�A?��(������R=f��>��	?\�?>�0������� ��>B5�?g�?��L=��W��w�ZXe?��<��F���ݻ��=eؤ=��=����}J>�>�>q���A�o(ܽ^o4>���>�%� 6��!^�:��<�]>o�Խ ���5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�󉤻{���&V�}��=[��>c�>,������O��I��U��=ܬ��Tſͤ��D ���U�c��<M��O�'���ӽ�s��H���Q���4߽6ĥ=��J>�ߋ>)�>��&>D�5>�a?��?q��>;��=/g��ᄾ�վP\��׶k��_̽����U�1������޾�!ܾ�E�uy�+��PQ־IvD���>%RW��֓�qF3�S�R��F��A?(�(>@���/D��t����Y-��X�=.y�������*6��}����?_�Q?����ISU����OM�;x��<?f�۽����.���n�=0(:=��=x[�>�z�;�����5�v	d���A?u�?�輾"پ�c�=^u�{e���*?��?�]T>̨��?㤱�&���e�=�� ?#r�>�?���>�դ���n�'9?Oo]?U�*�
����&9>�Q������i��"�r>7D���kB�u�==jk�qC�v�=t���kz#��^?cU�>�c��O�	���7潙�s=xH�?l}^?g�>��$?~4\?�?>�ܾuJ�_�϶=�^H?�"�?	C>�>����=E��O?�rs?��7>B7�����^ ��yW��L?2g?�?$�\�0�����U��wD_?��v?�'^�G7���)���V�ݸ�>B��>��>��9�Aҳ>�=?�"�����n���_4��՞?"L@���?�IH<M �.v�=�r?O�>�P��3Ǿ�������N�t=�\�>�����u�8���1�q�8?9Q�?���>炾]����=��-R�?H\�?6����&�<ڴ�&m����W2=���=��&��fB�h���`=��1ľ�2�x放����ǈ>{T@�-۽���>�Y� ]ῥE˿�|�m����d��$?˶�>�R½d����_k���k�`F�tBA�P^j�~ͣ>��> ��(���.|��v;����C'�>�Ӽ҇�>j?N��i��>h��s(<�
�>���>�ɇ>)���8L��ҡ�?Lk���Ϳ�Ğ��@���V?���?co�?�*!?M�<�}���s��#+���E?�Oq?	�Y?�/�7�X�c�)�4�p?.<�S�^���0�w1����=дw?�'?��w�<D��|>
��>��>����ʿ���k���~�?�T�?��;���>w��?K�*?$Y'��
��-�}��g>��ŷ=]~k?p<�=�¾���-m������E?2.?Ķ���)�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>eH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?7$�>��?]o�=�a�>oe�=B�-��k#>E!�=��>��?d�M?�K�>�U�=��8��/�O[F��GR�K$�@�C��>M�a?҂L?`Lb>����2��!��uͽ�c1�R�-X@���,��߽�'5>1�=>�>[�D��Ӿ,�*?u�:���տ9Ԓ��W�D�9?p}�>�#?���b�ž��<�oX?k>�>t㾛?��KǗ���E�$Ʈ?ɱ�?�d�>e�̾�N�=�_7>�`r>�v�=(D�=ni��Q׸���>��7?�ͼ�Ku��`��N>并?3	@䄯?�ye�	?n��P���a~���i�6����=��7?)/��z>��>��=�nv����� �s����>OB�?�{�?3��>��l?�o��B���1=PL�>2�k?�s?<�o���B>�?'������L��f?��
@Ju@n�^?I%��u4��jf������h?�=��=�tT>�L0�� %=fT�=�0���N����>A��>��>�>]�R>��>��=�B���!�n���d!��3KN�v�"�;��ãn� �߾o;�h�nа���j�c����$=��:��s�}�B����@l�=o�U?��Q?qo?�W ?�w�ު!>����= �n3s=OĆ>i�1?�J?0a+?��=�����2d�Gk���1���������>�;B>���>�:�>{��>Z�;q�I>.�?>���>��>#�<=d���e=�SQ>d�>���>x��>���>���<�������w�v��]�=�l�����?��|��N�Tj{�߸ξ��>�]>UW<?���=tŅ��;㿷貿�S?���� ̾��L��{�>��2?P"q?��?��Ծ�1���}>-��y3��	Ȳ<�x^�^f�S�C��P>�x?��f>�u>E�3� e8���P�@|��<j|>}36?�趾/C9���u�\�H�cݾ�FM>{ž>�D�]k�M������ui���{=6x:?x�?�7��Wⰾg�u�FC���PR>Y;\>�W=lg�=rXM>^c���ƽ�H�ki.=��=F�^>tW?�>�y�=���>������x�\(�>��B>�w>�C?Q?ڻ�Bp��M���I�tۃ>.��>��>�>C�c�YO>�x�>:ev>C�<Q`,���>��/B���c>�|�T���3�h�Z4�={��n>�I�<�H/���i�[PH=�~?���+䈿���d���lD?R+?� �=�F<��"�< ���H��C�?n�@m�?��	��V�I�?�@�?��)��=}�>׫>�ξA�L��?��ŽFǢ�ɔ	�$)#�hS�?��?��/�Yʋ�7l��6>	_%?��Ӿ�j�>e���Z��c����u���#=���>�:H?�X��l�O��>��v
?�?tZ�k���3�ȿ}v�K��>6�?���?Q�m��?��C@���>ˠ�?�iY?�oi>�i۾�bZ�ي�>M�@?R?�>b:���'���?�߶?���?_"H>���?is?�>侊���1��u���኿�5�=F�0�}%�>!�>ӟľ�@��Β��S��e�i����~d>>'=$J�>9������A�=L����1���b^��L�>�Ep>)(K>([�>��>�A�>5�>�*=i�|�oŀ�Ȥ����K?���?-���2n��N�<Z��=)�^��&?�I4? k[�}�Ͼ�ը>�\?k?�[?d�>=��P>��G迿7~��H��<��K>*4�>�H�>�$���FK>��Ծ�4D�cp�>�ϗ>�����?ھ�,��WS��GB�>�e!?���>�Ү=��?�G? �>�k�>�M��Ǒ��3C�o�>�b�>#?ꨅ?��?���j��瓿喿�t_�C�u>�|s??a<�>5㋿=���N9`�Iay��-A�
˄?�ڀ?���d!?#��?�b?�Z?X�>�������Gf0�z�>a"?	|���A�#�&�Gq���?��?���>|�����ѽ{��#�����?r[?a�&?pu��`�������< I$��遻b��;\\K���>�4>MS����=��>v�=�1n��9��|C<�=���>�]�=�d4�l�.?�����`�+��=��q�p�O����>$wS>��;U>_?4}!�Qm�����9�������?Q��?��?��e���D?��?Q�?�=�>|�������x��e���,�e8>��>����S��������=���9��Ո���5��c�>��>��@?�4?��I=�!�>C&��=�þ3Z\���!���e��&�X���s־L�<������ս������Ͼ6���q6�<�;8��">� ?)�X>�Y>��>��#����>�LG>\�U> ��>�n�>��%>l�~>!�&�}!ӽ�MR?����
�'���辞���T1B?�rd?�?�>�Vi���������?4��?p�?sv>yh��&+��t?N�>���)l
? �:=e���<lV������Z������>�;׽�:�3M��~f��g
?Y7?����x̾(f׽�����m�<��?5-?Zh0���E��f�|AX���T�>��;�>&�f雾q0�	d�tӒ���{��Մ�j����T=��$?=+�?�.��>�Ӿ_=���Ox�O�=�� �>I�>���>�(�>�ku>�����>RZ�4���W��U��>4~?�RK>�.O?�9?D? �P?H��>��>h����h�>G�n=�>��>��9?EN?��0?XD?̂<?��>>F~���m��Ͼ&K�> #?�Z$?�?{�?vW���'��^����?O�D�Y���=���<�2	��q9���=P@>G ?��vv8����]Hm>*�7?C��>���>�|��:#���W�<#��>7f
?���>������q�6����>���?��l��<�E)>[7�=*��k𗺌��=�}Ǽ�r�=젉���>�k�<�Ȼ=���=-�6��ɰ9��5;11�;^�<���>�?t��>K7�>x���� �A���ñ={PZ>�S>h�>�پCt������g���y>{q�?�[�?1�f=��=5�=l��畿�����0����<�?C�#?�{T?�M�?C�=?��#?' >�G��(���6������-�?�!,?ω�>F��v�ʾ��"�3�!�?e[?�<a�ȷ�8;)���¾��Խh�>"\/��.~�x��ED�&텻���E{��?��?翝?�A�I�6��y�ؿ��XZ��ΔC?� �>�X�>��>��)���g�6%��.;>v��>R?O��>�<H?L�z?oM^?9,I=F��p��E��+>��B>�y?-��?�}4?@�?�N�>USr>��X��M������$m7�r �;PB��m<K�>��>6 �>v��=���r����EFG���g�'�>��!?�4�>,�^>�=~�ν��H?��>������3������������r?�}�?�<0?=�� ���?�����Pi�>3Ƨ?.Ԣ?��+?i���>b����2���݋��C�>��>*�>��=���=9d>׶|>�>|Ҁ�Bh�&=3����9�?�@H?ҝ=��Ŀ+�p�~/m��S��GD�<����Q�a�{���H`�/ƒ=m%�����b����Y�ҟ�Θ���n���˛��{����>y�}=�9�=���=W��<��Ǽ`��<�|H=� �<^�=�ds��]w<B6�/���Y��U����F<cK=���	�;oa?8F7?:F(?iO?D.�>�L>rh�9q;>�Pҽާ	?��=�l��\7���"5�Y ߾~둾3ܹ�C�׾�O����H4�=������=��,>��>PK�<y��=��h��1
=@<@��=�6�=ו>��R=l�>,(>o1>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�F7>�E>$�R��b1�j�[�wb���Y��!?�';�m̾���>v��=�߾3�ƾ8�.=~@6>��b=���4\�a��=��z�vW;=&�k=t��>��C>��=u�6�=�H=��=;�O>�Z��l�6�*�gn3=$��=`�b>��%>���>h�? ?�.i?�|X>��W��� ��|�к�>��x��U�>| ļwG=�%��>(�(?q�*?p1?=��>��Y=��>�>���{T����	�=���!>л�?�?R(?rl���hƼ�*پ�BA�0`��"?F�[?��?�T�>�U����9Y&���.�"����u4��+=�mr��QU�I���Hm�2�㽲�=�p�>���>��>:Ty>�9>��N>��>��>�6�<yp�=<ጻ���<� �����="�����<�vż����u&�7�+�3�����;���;I�]<Q��;�+>�׳>�U�>�h�>��(>?����?>��w�x�-��r>��ؾ߼.�c2<��Q���f9��-��7�=�T>��켙$��&r�>�=[>���>���?A�d?�v>rƾ:���偿7��D־���=ʹ>����j���K��;��y����>A��>�l�>w.n>�l(���>�h�=��޾oX5���>0(��Lj+�A���>r�xͤ�AS���wi��&;f�B? 
�����=ܯz?O2I?��?>E�>�@���׾Ҵ.>���J��<����Mt�l��:?�K"?�6�>���E�_D̾����޷>�4I���O�j����0��?�3Ƿ�f��>	諭��о�%3�f��c���j�B��Ir�I�>��O?��?H3b��V���WO���� F��s?}g?�)�>�O?[=?��;r�Jt��<_�=�n?ҳ�?p<�?�>�ɽ���=���>��>���?���?&>q?�k���>˽M�<+�;�_=>�p�<u�>�W>��5?�L�>3�>�d�C���CϾI꾃� ���=;6<v��>���>�;l=�[�>T�O>jC >�H>1�>�j�>8^�>�>^H>=���:���?UM�=��>3_+?sv�>�=��%��W<L���,z@�hc8�$̿�d���n��2<�� >k,��Պ�>����L�?&�z>��&��i?�4!(���)>�V5>�����z�>��=\Y*>~3�>�Q�>`�`=�h>��>�?Ӿl�>���ph!��2C�xR���Ѿ�mz>ϕ��f&���������I�J^��[_�	j�,��iE=�x��<fI�?b����k���)�l�����?�[�>y%6?qٌ�U����>���>�Ѝ>L������Í�e��?���?c>'.�>F�W?q�?%$1�N3��/Z���u�� A��d���`�3ߍ�����F�
��G��K�_?K�x?�[A?ݚ�<��y>H��?j�%�f�����>s/��;��y==�!�>���`��AӾ>lþ�Z��F>��o?x�?p4?�DV���]�-ƚ>�:0?Y�?��l?U>?�o6?=d#�&!?ʨA>Gk�>_�?7>2?uS�>X3?���>�ݜ>Ę���z=�����YQ��zx�(}��|/�6�+=[�=�ܰ��==^�=9A
>ߐ��̖����>H��<W~�=�!>��1>iߤ<%+>תf?��?8Db>�G.?W�ٽz���S��Pc1?�a>�T��?W��GS�~��Gw>U?u?'
�?��7?�]W>��-�7��6�=�>��s>LC�>���>�pD�{)��H��B�="�=��>|��:¥�7F���M�:CȻ��">L��>1|>�ɍ�3�'>)u���Fz�v�d>o�Q��Ⱥ�G�S�"�G���1���v��C�>��K?��?2��=2Y�{��|Ef�`&)?�^<?�UM?�?�=Z�۾��9�D�J�!N�\��>}L�<<��(������8�:��g�:¤s>�6��������~>���7<�a�w�C�3�����h�d=6��2�<� 
��־��X��7>)O>�`��*X�({���2���B_?7�������v�����H9>�H�>mg�>@n��<����>�E�����=0��>�g\>�%%�k��hH�&_�_�>�(:?�BZ?��?DS��B ~���O���Bu���p����$?~��>��>PV>�j��Es��V���CX���+��3�>�x�>���{YO�d��O,���O�E>�>W��>�l�=��?y{Q?�c?��^?��4?(#?�2i>�Q�'L���;&?���?r�=�iԽ�U�b9�]*F����>�s)?$�B�'�>ϥ?c�?{�&?�oQ?:�?�M>�� �)&@�F��> Y�>P�W�#a����_>��J?2��>�=Y?�˃?�=>�u5�����`�����=mf>��2?�'#?�?b��>�'?Bc��fa�15�>"'E?b'�?��s?��b=!+?Ÿ�>��>3�=�U�>rY�>�?JRS?I:w??P��>f"�_l��č޽"Aƽ��G���9�L =	`=u ��Ƈ��N���XO=HE;���s>�<�q��L/���
?��of����>�m>������->�Mƾ3���?>��u��矾��s0��d�=*ŀ>�� ?��>N#�Ǚ�=���>���>���'?�?�?4��;F�a���ܾ��R����>X<B?�ѽ=�Vn��)��(�v�ȉl=��l?F�]?f#]�5@����b?��]?W�A=���þ<"c���龌�O?C�
?��G�^	�>�	?��q?^��>��e��5n�����3b�J�j� ��=�u�>HU���d��3�>Ɨ7?4?�> c>�=�۾��w��Q���"?,�?��?h�?:*>F�n�'࿣��\:��u3^?	}�>�P���#?5�����Ͼ�/���͎��U�<���ҫ����������(%��6���ֽ��=��?P�r?cq?�_?���c��C^�A��R�U����6��[�E���D��C���n�MI��u���՘��JJ=��I��,P��,�?�?@�}�8?��i����F��.J>Y�վ��c��9�=���&'�v��~���C�(�?�e� ?��>��>A�8?T����H�0J�jF&����2s�>n�>oθ>_E�>������Ҿҽ���BA�^�<s8G>��W?�@?l�?��#���E����$��S�9�ٱ���V?�w�>�[�=@�K�,���F���8�(�>�9J�&$������>�St?�J�>ˀ�>�u?A��>9�������s���x������ѧ=�.?>�>���>��n����Ţ�>l?�t�>f��>"v���!�ҝ|���Ƚ�R�>_�>�	?<o>:2���Z��ߎ�V���`X8��v�=�"h?t%���*a�*�>��Q?��9Koq<�j�>8ex�� ��N�Q�(��>��?�m�=Z,4>�ľZM
�'{����l8??��>ț���0���@>*y*?��?�y>��}?]?f���
y�<�)?z�I?B�C?�8D?�&�>�>03����׽�y!�y�:��d>_D>���<�,�=�g��Um�A'H�Sً<1�=���;�E��<Ò�Ƹt<��<�~�=c�뿏)X�
�о~��t� �4m� \��0,/���^ H��$��W���1��M�<B�=M��^7����j�����?YA	@�Jᾙ������RY����$s�>��w���E��G��y3�U��X�������ߐ$�eQb�K�i��ې���J?�����οV謹�O���h[?&V?o�?����өT�P�M��}�=�+?��=e۲� ��Պǿnh�?��>�D���-�=�l�>��b>3�;"��>y����̾�b���+?��D?�$�>�B��mjȿ�t��Lٽ"6�?�@��A?��(�x�쾠�U=���>��	?�?>�Z1��<�_հ��I�>+6�?���?ѲL=I�W��H	��e?ȓ<��F��޻�,�=3�=#=c��iJ>�1�>GP�<A���ܽN�4>�ޅ>�m"����@s^�^t�<�Y]>�Hֽ%���8Մ?{\��f���/��T��@U>��T?�*�>�:�=Ų,?<7H�=}Ͽ�\��*a?�0�?��?4�(?Xڿ��ؚ>x�ܾy�M?:D6?��>�d&��t�`��=�2Ἰ�������&V����=6��>L�>��,�ɋ���O��Q�����=rp�<Oǿ-L$��&��L�<m.��z`V��������c*^�p��p\n�_��K�v=g��=zS>T�>&�U>�Y>z�X?�n?�Y�>�>v@������Ͼ_R������a�p �����B椾Խ�F~�NL
�j�����V�˾�>�B'
>�_[�����=2��GJ��H���?��=Fi;[D�lF�3z��Rg�P=L}��Ͼi9������?kC?+~���wb�Л�q�@=ή���^?06��D��p~���|�=��k��=�z�>�=���#�7��y�0??̨?b���9�^��=����E麽}Z)?�?�~F=��}>��9?�������D��>N�e>�L�>���>�G�>��ƾ^�<g�X?�|F?94	;�B��'Ђ�� D�)Fc��U��:%>�-���4�;���>,��}(�����F{����=_3c?!�e>;�?�S%�^^����~����=��Y?Z[?E��>�pb?e� ?������/*H��ǡ�;}^>�f?0�Z?�H>��;����`���XD?�@�?oC>���k��P�����'?�ۃ?$H?Kr>P�s�l����V�8+?y�w?<M\�H���T�F-b��U�>k�>&G�>\�6�]�>@�;?'M&�v��_��� 
1�i�?��@X��?*�;��7�!=��>��>�O��,̾�۽xm��ʄ=�w�>q����r������K�(m5?Q�?���>�?������!>WǶ���?@��?r������6��/#R�T���V]>!L�=/=N�7;V�,!g���þ�����p؋=k�m>f	@K�E���>�B��5��N˿�X��n��)��H�D?��>4�a�Cc���Z���K�����P4�[
��L��>��>�����탾�}���>��ϼ�B�>!�<<���>�/�����h-���ߒ;��>���>s��>i�������?ol��N6Ͽ�˞�����L?�H�?-�?��?�|\=L3j�V�g��B�5�??��k?��_?��#<qQ�B�g�Cxy?�'�p�R��W;�Ve7��=�O?�� ?��c���`�A��>J)�>2^�>����Mɿ������nX�?�Y�?D�b'�>`�?8� ?�+�?N��+�*P�gӌ�]"w?�D\>�R��^��xO���ȾVH-?�Z?!3�T��`�_?.�a�W�p���-���ƽ�ۡ>��0��e\�GN�� ���Xe����@y����?I^�?a�?��� #�S6%? �>j����8Ǿ
�<ɀ�>�(�>)*N>�G_���u>����:�i	>���?�~�?Cj?��������V>�}?83�>@T�?��1>��>��=�о��W	��@>���=�]���v
?,~V?N��>k�=���#2�D�<���1�2־�F����>]bo?��G?��>��r�����*&��x5�5c�KE��8B���h ������>Ol�=�M>�<%�|��?O|�ٔؿi��Tl'�24?cȃ>�
?���s�t�WZ�'<_?S��>�-�a+���&���i����?�B�?��?��׾&Lʼ�$>�ϭ>0�>ĴԽ%3������[8>_�B?�*��F��n�o�%�>���?�@JӮ?��h��	?��M��`V~� ��� 7���=�7?��y�z>��>�=�qv�㸪��s�!ж>�C�?ku�?A��>��l?ۀo���B��u1=mA�>ߏk?|?:�l�����B>��?�������L��f?Z�
@�u@ǚ^?.좿�ۿ�����٣�⬫��k>ߡ=��\>�G-���3=/3<�C�S4Y<T<�={�>�>N6�>���>�Y/>�6�=�x��G�&��:���V��ӭ<�ɣ�����k�gh��օ�W��G���:�ž����y���Zh��O4�h������B�=ڲU?�R?�p?�� ?K�x��>����$!=��#�)��=�0�>HR2?ֈL?ݤ*?�c�=����g�d�HV��,C��f���>�VI>/k�>�-�>�>�h :EJ>^A?>V��>^%>H4'=b���S�=�CO>l^�>���>Ǆ�>�i�>8������b¿?Ah�Nѩ<̺S����?s9��u;�;����ܾ��G˨>��L?���=�ه��
Կ$ֿ��Z?)����
�Q5��~~�>�|-?�\?7��>��J��J��<%�Ε�`6>{�y;�[�������:>]+J?��f>u>V�3�d8���P��v��Qr|>26?����rH9�]�u�t�H�haݾ�@M>㴾>�QE��n�e������xi��}{=�u:?�?�4���԰��u�=B��m[R>�5\>^i=iw�=�]M>ac��ƽ�H���.=��= �^>g�?~^ >�W����>1!��JG(��Ӷ>HV>yvL>��G?'a?��2��8����A�ܽ�0�>���>q�>j��=��H�+�=>V�>VY�>(���������Q����Lj>bEV���T���ju=e��� �=�Y�=�<���&��=�~?���e����_�G<����D?#?n'�=�LF<N�"�3 ���Y��Q�?�@\d�?˂	�D�V���?L �?ĝ��"�=3d�>۫>��;!)L�D�?��Ľ.���D�	��#��J�?K�?'�0�Yˋ��
l�G�>b�%?"*ӾQh�>}x��Z�������u�|�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾;`Z����>һ@?�R?�>�9��'���?�޶?֯�?��;>F�?�Oi?+�>m]��M.��ɴ��Q��.-�=DUl���>��=N�㾫�:�B����7����X�Z�Ω{>V=m��>R(��c�¾��</hF������F#���>��B>�>E�>� ?�R�>��g>�='\�9rw��?��}�K?���?���2n�BM�<���=a�^��&?{I4?Xl[�T�Ͼ�ը>�\?m?�[?�c�>F��H>��<迿7~��a��<��K>94�>�H�>�$��zFK>��Ծ�4D�Up�>�ϗ>v����?ھ-��<P��5B�>�e!?���>jҮ=��?��?��> ��>��P�����)�R����>�>�??o��?�S/?�绾j���ڑ�I$��#�f��+'>�%h?�E?qD�>���H���)=pM�ԥ��ڧr?��7?�yx��{?�%�?�v6?i W?V��>W����;���d>��!?����A�N&����~?�P?���>97����ս�Qּ����~��g�?�(\?!A&?K���*a��¾9�<�"���U��7�;w{D�^�>��>����'��=�
>�հ=�Mm�?E6�e�f<�i�=\�>��=�.7��p���2?�6ý����K�<u�m�5�H�c��>O~P>��Ѿ��`?@�4��)}�������0∾8l�?�?s�?�����g�9=?�,�?=?�9�>�㩾���#�߾�<�A~���?3��=�=�h>ߢͽ�h��{᛿� ��k�������v��w�?N��>l	?$	&?[�>JM:>��r�Q�A�����*���l�>H,�49*��	��-�X�Ͼ����۠&��V��r7c��cA>O���6�=���>J��>��{>���>.Z�v�`>Ah�>1>ǔ�>Ō�>���>Y��>0$����MR?�����'����I����2B? qd?>;�>!Bi����Z��D�?��?0r�?1v>;�h��/+�p?�?�>����n
?v�:=#^�R�<A_�����5���^�Ӭ�>�׽M:�M��pf�]c
?�-?9���߀̾/%׽�㛾��-=L^�?)?�,���M�P�m���U�MPN�pSżŮk������� �&�n�����v������b�&��X=�(?D"�?9����9従����o���A��i>>��>a�>#�>ǪH>qg�%2���a��$�ٓ����>[x?�E�>�1J?Ë<?VQO?��J?/P�>���>����E�>#��<���>I1�>�7?=.+?s.?��?�n)?�wf>���m���о��?}�?�3?�A ?� ?	�_ܽ d�Fu��Sp�����w�=���<^[�?����K=��C>\?Xd�U�8�����ˑj>s[7?�Y�>���>+��47M�<%E�>I�
?�`�>^���Nkr��^���>A��?g��=e�)>���=Ɩ��BҺ�	�=�Y��˖�=� ���v;�^4 <y��=Wj�=�m�9���Q�:8��;1Ʈ<"��>��?@r�>�<�>G��դ ����Y�=d$Y>�0S>�>l6پQy���%����g��sy>�u�?){�?½f=��=Y��=�p���8������������<��?�H#?f@T?���?��=?�f#?��>�#�JG��J^��,��o�?� ,?Z��>P��}�ʾn�̉3�K�?}[?�;a���;9)���¾��Խ8�>[/��/~����D��A�����]|��D��?���?9%A���6��y�t���\��v�C?�$�>�W�>��>8�)���g��$��3;>o��>�
R?�۹>&nN?Qse?e";?uK[;1�j�0���fv��������=rX?�O�?���?��?�s�>��м��ľ����&?��g,��+m��2����<��>>C��>4�>��>��<�JD��@������=v�>���>��&>���>0�k>ࠩ���U?�	�>y
��
¾˶��eyξ��d=QX?Y�?�]R?N�u>5���_�0��x�>�p�?)q�?��%??m���E>�?�*����޾bC�>�I�>J�>Vv�<
q�l��>ʐj>O��>+4��M ������P���>�f?��=��ſ�q�f�p��X��U�e<*뒾7e�x����[�~��=�u�� �����ſ[�{ڠ�/����Ե��ǜ��~{����>L�=���=���=�<Ǽ/�<�TJ=��<��=
Rq���m<f 8��Żo����b<�iI=�m뻆�ξI~?�uI?�)?�lC?��z>X$>)B���>�8���m?Nz\>svc���ž��<��y��摾�\ھ*�Ӿ&�d������>X���>+94>� �='O��E�=�i=co�=����r�0=��=��=b��=Y��=֐>��>�6w?G�������4Q�[罗�:?�8�>�z�=;�ƾ�@?��>>�2�������b��-?z��?�T�?u�? ti��d�>��:㎽�p�=V���t>2>7��=p�2�5��>��J>����J�����o4�?��@|�??�ዿ��Ͽ2a/>M�7>
/>�R�3{1���\���b�1Z�'�!?J2;��	̾�4�>_U�=�߾Ýƾ+�.=�6><�b=B���=\���=`�z���;=im=꼉>��C>5޹=�௽��=GJG=ʠ�=0�O>�R����8���+�\3=ڧ�=0b>&>���>	�?�t-?��t?�m>?����5�(�x�g�>K�6���>�Nx����<�"R>�o?ɀN?�9E?��[>�=�=$��>�Cb>�"�
�|�����2׾�� >��?r��?H�
?�i�=10��pY���)���Y���U?��F?g��>QΊ>�U����,Y&���.�d���&	0��+=anr��PU�����<m���F�=�p�>���>��>�Ty>��9>?�N>x�>��>y5�<vp�=F猻Bµ<������=d�����<tżn����a&���+�
�����;���;>�]<٠�;9��=���>�"q>��>_j6>�����/�=�h�A�Q���!>j�|\���b��Tk�� 7�:���OU6=�C">!��Y8��m�?h�]>^8U>�;�?��b?�c�=���l�澉��-�
�����%A�sY�=6'��V�x/x��Q��!ྦྷ��>�'�>EB�>��l>^�+��:?�Poq=K���Z5����>ư���|�����p�H
��$�;i�g.��LtD?�6�����=S�}?{�I?��?V��>T.����ؾ��/>
&��2�=�Z�br�����h�?��&?Z��>���v�D���Ǿ>����ܸ>	�2��NP�����2�<U������٩>����~Ӿq�3������b?�hYh�vn�>}!O?��?�wd�d����Q�uB����4�?[�g?�p�>�
?D?0͙������E/�=�Tt?A�?��?b>3v��*�����>`�>!�?�2�?��t?N׾���>��'���=�*���>\�=���=/ۗ=�?F�>2�?�Gr�=*��'
��=�2-�Yq=�0l���=�ɓ>]ʐ>���=�ܼL'c>�P?���>��R>���>ѻ�>\�>�����$���$?��=�k�>�r<?p	�>�)�<_,�����eUV�P``�#�:�8}:������kļt��8=�A��>����伐?��>�d���?<?���=���>
lc>}�߽�	?�h>yP�>x_�>B�>6*>o.�>�8�><CӾ}y>H��f!�!,C�ƀR���Ѿ�z>j����
&����}��X8I��k��f�j�.��==�D��<�G�?T���9�k��)������?�]�>k6?)،�5��J�>��>oʍ>6K��Y����Ǎ��g���?K��?/�a>��>4�W?7�?�90��?3�!.Z��!u���@��Ke�*~`�	�������&�
��<����_?��x?��@?���<�^y>�m�?�y%�]��yO�>�/���:�ڂG=��>�t��_f^�:ZҾ2Nþv��ZF>�3p?E"�?�?��T�6h߾]�>��?�(
?���?Z�F?��]?��G���?�76>q�>�;�>feL?�q?�O4?,6J=T �>eB����>�ýLᐾʼ�=W=H>��>\�=�?�=�>K���oY=8H�Y�½=�=���=g�'>߈�=�=\=��U��������?JY?BAl>�bQ?�Ͻ,���|!�q?y?���~XN��y)�>��d�<��O�>,�?,��?���>]Y{>Cm:���C�/�i=����5P=��>�"?M���'[���=���=J;,>ι>-�ؽ^&���u�%gP� ��<��#>���>��|>&Q���(>l,����y��~c>�Q��s��7�R�9�G�U�1�_Hv�"�>O�K?Ԝ?z��=����9���Yf��/)?�<?>M?��?"��=N�۾�:�0�J������>��<�%	��������:���S:�ps>1����	����>��5�o`��:|���#�Ax�����$�b�<�!�A��zȐ>:Z>�Y���h-�t��ӎ��ruu?̕�������W���Ⱦj��>G�u=`?	��=:#�g:E�P2��-�@>�Q�>㾆>,�=w�PW�L��Qw�>��D?�)_?�?�F���r�"ZC�U���.`��H
Լ��?���>��?�=>熬=�7��˦��(d���E����>��>�����G��m�����q$�)[�>=�?�>�D?�Q?sv?�?`?�)?�,?��>�a���f���?&??���=�Խ�T�@�8�F����>ց)?˸B����> �?
�?��&?��Q?��?�>ǫ ��>@����>�Y�>�W��b��� `>ɨJ?b��>C9Y?Ӄ?$�=>ԃ5��ᢾ�驽�l�=�>��2?7#?��?���>��>�]����<Ԩ>�W?%~�?Wl?�P=ض?-r�>�n�>�Ύ=._�>^��>A?��[?À?Q\?qV�>Ӏ]<9��2�彏9.�3�r�*�b���;И�=�F�mA���n�C�5=��;q�Ƽ�e<S'��X�̽)�밋<��>©>L���[_>�A��T[���]'>=ɶ�[Ǜ�)�t�v)�SP=\=u>�h�>��>M���=1�>�2�>�R��m"?�O?}s!?���<�3^��ξQ/���;�>� 5?n�N=��o�˕���{����<
�e?�la?��\�� ���b?I�]?*	�.�<���þ��c�m��o�O?��
?��G��F�>v0?��q?;
�>1Of��:n����h"b�F6j�̶=uj�>(?���d����>��7?N��>�b>�F�=��۾�w�����`W?mʌ?���?�ۊ?�z)>�n�@��+��\��Y�a?�?�>Bɳ�\&&?`ج���̾�����b���}��@���m��t:��˵���9��"���ýb>Ҵ?�ph?�{?%^d?����xd��^�{�|�ON�8��6��<�>��B���C��n��X�A���帛��=�{n���D�ʴ?��?%�o���>���|��~�ؾ�W>T���
JĽ^��=�Ε�^�e�;�b��j���u���$?�̦>���>��G?
=��f�B�-�6��54�� ��m>�C�>	�>���>�P�t<b��X�wjؾ�����E<��>H�T?ٺF?"7{?~J&�Cz0�A���xξLT�A"��ì�>�sj>�[�>���O�Y<�eQ�ښB�2S���P��9"��8�'���c?�-g>���>��?���>��ؾH���(����ES���������r]?�[�>�$�>ֆ����	��&�>>c?���>$�>^���m'����y̻>��>JR�>n�?��>X�
��I�3���*���A����=w�d?�np�P�`��Bu>c�R?ŹD=p��=�Ն>Dؽ��������Z�U��<�?�Xz���S>bӳ��,�6�g�с��+?�
??���+��By>]7'?g��>���>��?�ư><0��%��:w?X`U?x9G?E)G?�s�>���=C�ŽA7ƽAj"��2�<E�>�3[>��Z=,��=����^���&���8=^��=j�Ƽ�g��=$d<���|�;���<�J+>N�ῡ�9��̾Wz �_��� �r��x�����tN'� Z��.Bv�*�O�<�<(������s��+����%�?6M@f��&Tؾ�Ŝ�~Vo�����[?>����6�K�q}Ծ	�|��þȸ��m��{O��T�L�[��y�K�4?n��.�Ͽ�a��S�<�4?��'?¿�?�6�w�|�Q�P��+p>r�>c��<T��z��� ǿ+Ǘ��;?�n�>�xd>YE�>Hu�=�:<>�9?�DZ�ޥ��xȈ=BV?�a?�W?�^���_ܿ蝿��>ݳ�?~�@O�A? �(����d�U=Y��>8�	?��?>�g1��1��Ȱ�mN�>/6�?[��?ɗL=��W�P��ƅe?�	<2�F�8*޻$3�=g�=ן=%��|bJ>YG�>�J�rA���ܽ��4>��>ݭ"�_���\^��|�<]>ֽ����5Մ?+{\��f���/��T��U>��T?�*�>a:�=��,?X7H�`}Ͽ�\��*a?�0�?���?&�(?2ۿ��ؚ>��ܾ��M?^D6?���>�d&��t�݅�=F6�z���~���&V����=Y��>b�>��,�����O�J��d��=H��ǿi�!�|D�v��<d��v�>�Cw������������SU�@ׅ�Mh�=���=&>�={>�X0>f�M>��\?5
|?���>4��=ͳ
��ߍ�H�̾fP�H%v���2(����-�Kf��+N�3޾õ�q4�{���Ǿ4\B���)>��V�tS��vg(���Z�vX?��J?J��=3���T#N�����̩�s�i����<9�㽅tܾ��@��t���1�?	$K?A�����T�9u����<�#�++P?����������%t�=��<��I==�>c� >ޝ�T;�}�d�h_??�?
$׾ρF��+B>��J����,?��?+N9>s@�>�}B?�)/���9���~>�>ۃ�>�}�>k��>5�ľN����J?�a?�C��o��Y��<@s�IU̾J7<#>�����s9=0y�>^(⽘0��U#�,1��>�W�2�\?��>]�'�B�����N��)�=�P?�J?�{�>�=d?��R?[[��ae޾m�&�5�ƾk��=�8j?�X??�=�s<�5���w���4?��2?��@=����!R�rT�J�Ծ�?�@X?�o?$i=���o§����#`E?��y?��V��!����i�S�?��>���>�
�>� ���>��6?_` ��s���i��.�*���?I�@�B�?�m��+��5�=���>ٲ�>��0�����q��^ ��R�Z=���>�@��Sg��4�Щ%�x#5?��w?���>�gq�������=�1��?Ŭ?���?���I<�?��j�
����<�@�=O6��5�'`��w9�vEǾ w��c���sg�a��>��@/��)��>\9��>�fOϿ����)�ɾ�j�Ii?Uީ>*vؽ�塾��i���s��F��bH�y�����>Y6>�c���u���`{�D�;�����`�>�߼��>�M��<������ޚ;���>���>�h�>N~��xû�M^�?,y��Aο��������V?c��?��?��?�<�5m�d�{�-�L�E?%�p?٬[?���*K[�~�K�xSg?~���C���J���D�*�=�Y?\%?�ȁ�Nʴ���}>���>b��>W.9��̿m皿Y��Q��?:V�?��þ��>���?��?����(���R
�GC"�U�]��T�?�|�>l5;�|�H��f.�B��ww ?v@?vq����(�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>eH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?��>�	�?|��=�>�}�=F8��0y��~�(>���=݇���d?�7H?���>�Y�=��1��1��7C�z�M��'�H_C����>g�b?c�Q?	�i>�9̽Yl*��U%��2��0��I�a�_�^L�;����,>�>'>�'>C�a�ܾm�?�u���ؿ�i���'�054?&σ>�?�����t�����B_?��>6�U+���$���V�G��?WF�?4�?D�׾�/˼��>v��>I3�>^ ս�������e8>$�B?@3�E��4�o���>���?L�@AԮ?ti�)	?u�� 9��`�}����.8����=@�7?�B��dz>�"�>M?�=�v�+���m�s��O�>+4�?&)�?|��>�l?�Go��*C��9)=2��>(�j?V�?�'D����(sD>�'	?�������Rm�(re?��
@�y@lW^?�뢿�쿓f���⌾u���£�=��=�E>~�C���=���E�N�<��g>��?�0�>˅�>s�,>V�Y�d�=K���%����,��sG��c�(sﾗTE�|!��L���c �?Ē�E"���ǥ�#]<�^���H/�z��H���,��=��U?�Q?�
o?/�?!l��(>����G��<Q�%��4�=j��>ft0?�uL?��*?�q�=�a���c�v����`���W���b�>~L>p�>7��>�Ӯ>�V�;ڑJ>��A>�q�>���=6z/=�Ȫ;�=]�H>�8�>Ԅ�>���>ڼ�>(S=l�ɿ�V���r��MM=ߗξ�͙?84��t�?勵��о�X+=nX>+IU?\�=c�����俪�ɿoR?�����-�E��>� ?��;?��?��|���C��=о�yu?�Bw��$�{� ʥ�1�(�.�>B�-?�f>u>[�3�Me8���P��{��j|>�36?�鶾�D9���u���H��bݾ6GM>�þ>�D�
l�6������ui���{=x:?�?�:���᰾;�u��C��9QR>b8\>�R=�k�=�WM>�\c�N�ƽ�H�[m.=��=;�^>b ?,�&>,ɭ=���>�n���L���>��V>��/>�08?޿&?��]��	���\��۵$��4M>���>rm�>�>��>�~݇=���>�p>�aļ50��3��Q�S�x;{>�������J��;��{c�~&�=w�=�ō�g�T�?�]=�~?���X䈿��p��ymD?M-?�=�`F<х"������B��s�?��@l�?Ӄ	�B�V��?�@�?�
����=ڀ�>�֫>�ξB�L�m�?/ƽ�ʢ���	�� #�S�?�
�?�/��ˋ��l�:>�`%?�Ӿ�i�>+���Z��g���u���#=e��>g:H?mW����O��
>� y
??0]�:�����ȿa|v�Z��>�?���?�m�j?���@�l��>���?$hY?hi>�k۾"XZ���>��@?uR?m�>R=���'���?߶?�?��I>� �?ggs?�#�>�C~��G/�1/������mv�=�);Vܑ>�>����rdF��:��;L��wWj��5���c>pZ&=�n�>�}�W���7�=򳊽�b��dBv��:�>�l>��D>�,�>�
�>�`�>R��> !=�Y��P��⫕�|�K?���?���2n�>Q�<*��=\�^��&?oI4?�a[�2�Ͼ[ը>Ѻ\?g?�[?�c�>$��8>��9迿W~��֪�< �K>�4�>�H�>�%���FK><�Ծl5D�Ap�>�ϗ>8���?ھ	-���Z���A�>�e!?���>�Ю=�^?�]?
�> �>
o�w���-�c��
	?gV#?f�?4��?��@?�#��ﾓ���A��]�[��E�=��}?|�?|{�>�����&���f>������ɽ�&u?%=?�_�W�=?��?�I,?��e?U��>|�8�+驾f.��o�=v�!?`��A��M&�b��~?�P?���>�7��Q�ս�Jּ��������?�(\?�A&?����+a���¾�7�<<�"��U�c��;��D���>W�>񊈽*��=�>>װ=Om��F6���f<tk�=��>��=l.7�Et��69-?��v�~�d���=.n�\I�vˆ>Ywd>*�޾�;a?�^��Y��F裿ۘ�������?zλ?{�?9]����f��;?���?k�?Qg�>�������Y澑�`��n�"�LM�=��>2��<�鼾M¤�2/��d
�����"���>�Z�>5e?��(?��=Y�[>R���:�2����� !�v(t����"�A�	�6��("�U���U��=I���ž�
��dq=_�{�t��>Q/+?y�>�p+>��>	{3��$>��>~��<rz�>�\�>#��>>dO>"�R�#��4LR?9�����'����Ž���4B?_zd?GA�>��i�A������|�?G��?�n�?�"v>��h�W/+�Yp?�K�>����n
?x ;=����l�<D_�����9b�������>��ֽ�:��M�^�f��R
?�3?�Y��@u̾d׽�m�=����ٔ?3v.?`�Y��&8�+�c���=���<��[
�����9Z���%�k�h�)w����x�����B�8D�>)�!?_�?,&���搾��ξs����[��+�>�!?���>y�?�+>dr+�f��λV�B��m��r�>��\?�r>�}N?�V6?�F?Y?'��>˒�>�x���j�>��j:#�>���>nx'?�'?��3?�f?h�+?�i>�B۽�b���NҾjO?Js	?�&?Z" ?!��>4������*�$�.l;�=t�[����Ħ=���<�q
�aq�� �E=n#;>KX?R��	�8������k>V�7?{�>���>���;-��#��<��>��
?`E�>} ��}r�%c�V�>-��?��z=��)>���=@���8�Ѻ�Z�=H�����=�K���|;�0�<�=V��=�t�b/����:θ�;Z|�<���>��?ğ�>��>���O ��I��=i�Z>?jU>[>��ؾ�L��� ��qg���z>���?^��?`�d=���=OC�=���2ƾ����==��Q�<E�?7�"?9�S?|�?9�=?0#?R�>F���X��3����|����?'#,?�E�>|��[�ʾN��3�x�?Oj?�Pa�����)�x�¾D�Խ:q>�s/�0(~�/���-�C�˾�����6�����?㹝?�A���6�:}�3���_N��ϜC?���>��>���>��)�S�g��#�+(;>n�>��Q?=�>h�N?�Fz?��Y?|�D>Ze<�#����9��|�����>)D?���?�P�?Ԅv?yo�>Α�=��G�E<۾�&�}'����?p��V�=�+`>n8�>���>�t�>�Ƃ==	߽(ǽ��`����=;�">m��> �>+9�>FAu>o]<ݝa?tu>���6
׾��]�e�]�>��?{x�?3�i?��>U"��qh�� G�<v�=���?�`�?��F?�4���>>jے�z��O
��T�>��?l,�>��Z� �=:�?�w>/]�>� �>6c��q릾���=��"? ?xj����ſ�Jq���o�U֗�Nb<U�����c��#����[�1h�={�����&y��~1\�8M��ȯ��V=���n����{����>��=���=l�=q��<A��a�<�F=�M�<ej
=�p�d߃<��9�h�������	���t<�GN=xDʻ�k׾{�{?��E?Q`!?��M?>l�>d>�uƽ��>]����k?)K>-M���Ѫ����Cx����b���žs�Ͼ�a�����$�(>0]	���=�>���=N��<Q��=�(�=�Y�=_r�0�=`�>�)�=�I=��>�	�=8�=c<w?Ϗ��R����/Q��I�X�:?O�>��=�)ƾ�<@?��>>�$�������p�E ?<��?LW�?��?�i��R�>L䢾+T����=k����1> ��=�d2��h�>�AJ>g��5�������!�?�@�g??���Ͽ=�/>;z7>*7>J�R��1��1\��ab��_Z�֌!?sG;��G̾��>&��=5%߾F�ƾ�.=w6>�$b=0Y��K\��ə=e\{��(<=c4l=v��>FD>���=�=����=]�H=���=��O>Ȗ���6�9�+�°3=�$�=�b>�&>�]�>�(? �#?�bz?ؕ�>0������͘��q�>$k�<�N�>��,<d�;,�]>`�?x�0?6�:?Q��>^>=V�>i=�>�B�����q�P����=T�u?��~?WT�>�/P=�$$��L8�
�+�Y�<��;?2GU?I�>n�>�[�X��M��)�$U���߯����=f�j'��j#V���mH��5\'>���>�$�>lh�>�\u>e�>��>a��>^$�=�,�<x��<vu�8K�0<�I���H=1���a�=,;�����<���<m*G�a�������=�	�=A��z�>�>҄>n�>\f>J. ���>L�A�]�u���>�Ӿ_&h��u=��]i�C�H��S���e�=�\�>M%~��Ǐ�͜?�c->
�>���?�j?B=ĒV��Ҝ��f��~����h��=��e==ʸ��-��Vr��^R��������>)I�>���>�Ul>�[(�rA���n=��ھ�[8����>����6�}�"@��vn�L¤�6���sf�ץ�;&�??�҇��/�=�v|?�K?�ԏ?���>�+�� ;޾ݥ.>+ׂ���;�[��v��P����?�"?k��>5��)�C������ƹ�h��>�����K�#���X7���$<�g��$��>�Z��/ξ��?��텿�+��n�4��U���>Q?萪?TX�r�����`�9n�<۽�{?+�b?z�>� 	?$?����jD��ꄾR�	=�>?�?�?
P�?Y:�=չ�=Q��[��>��?��?�?FVp?1zG��>�?_;�>6������=0�>�2�=��=
H?U�	?7�?C{�����©꾪��3�X��=��=Zr�>6I�>�1o>���=Mɂ=g��=E�b>9��>�q�>��b>�У>��>��������X?6c=���>�d@?չ�>�ý=�N��ӣ�>�z�@f ��E�ǋĽ�~��\i��Yͽ+A}=�f�����>A���Ÿ�?<�>n!K���?���B5�7�R>i��=�ɽ���>��>q��>�ء>g��>�g!>���>�կ>�EӾ;}>D��'e!��,C�s�R�վѾbz>z����&�o��<x��r@I��m��g�mj�`.��x<=�t��<�G�?���F�k�L�)�������?D\�>�6?�ڌ�#��{�>��>�Ǎ>�J��F���_ȍ��gᾺ�?F��?��X>E�>'#H?�y(?`н��F��Q���i��,���R�B)P��މ�~q���	�̒���R?�n?1?��<��`>0u?��r˾'ϛ>_���1�N�o=�R�>��[bc�?Ú�����*s���~>��?*�?j6?�ҽE4׾���>��+?$�>{?E�2?�D]?k����}�>ǒV�@k�>̐�>��>}oE?�#?F]�>���>��-�U��=sp<�L�j��4���v��C	��� =��A>�r=UPR>�<!�<��&=���=vB�=�m)�+��<�_A�j辽��{=�Z>kIm?2N�>ؑs>'�i?����+�'�Q侅�?/Ǘ=�����m��'���þ�ؚ>J{?r֟?�+K?w�p>�'p��H���>��=��)>ݾ�>�Mz>L��~,P�_��>�7>n�d>��;ʵ�v�k�����O<:t�= ��>�p�>7q�g�n>�R��Z��1�=>iW��,��^��z9�=�9�;gn�g��>b�B?���>�i�=�pԾ��
��e��� ?G9?2Ec?��z?T�;=Ԯľ+�M�.I��C�sR>i�q���aa������2�RJ�=�#R>5󺾴lǾv5�>*1�Z�#��'o�gH)����!*��n����=2#	�;�73;�>��p>������&������h��.#x?#ѽ�d뾟|5�mt���ym>�
>|l?$\�U���C�V ���L>#ʔ>��g>�	I�c�� S����f�>��D?�2_?#o�?�Ã���r��C�!S���W����ż�?�Q�>� ?,wA>%��=�����Krd��&F�
��>��>�(�$GG�BJ�����$��]�>6�?��>т?�NR?a�
?�]`?;*??��>㴽���B&?ۇ�?���=��Խ��T�d9��F���>�)?�B�V��>�?��?��&?Y�Q?�?��>\� �??@����>�X�>��W�Ha��� `>?�J?̘�>�;Y?k҃?��=>��5�vꢾOé�jS�=�>x�2?t3#?�?	��>���>hЧ�{�>=�R�>8Fb?��?'�n?�<�=��?I>n��>��=���>���>�h?��U?:Ly?�N?�)�>�]e<TO��~O��4W��Sj[�:���±�;��f=�8�,��������<ݿ;尹��n?�X)�j���!Qa�Z�f<��>�x>~�/�'�u>�̾#Ǿw$>Q>�B�L̈��mP���_>�Z�>[�>*tl>2MY��r\=FD�>r��>�R���?��?�?�ӽD��6����e�X��>�2?�v�= C\�x[������`#=~�p?Jrl?�=�����'�b?a�]?]�=��þ��b�`��_�O?a�
?��G�|��>��~?��q?���>+�e��:n�/���:b��j��Ŷ=�o�>�U�W�d��C�>��7?H�>\�b>a�=�s۾�w��r��s??�?f��?���?�(*>?�n�m.࿪����w���^?�g�>���:�#?��9�dѾX�������(쨾�����┾󥨾iu)�J���ѽڌ�=��?�yq?�s?�a?ܗ�N;d�� ]��~��rS�)%�5��Q
D��VD�)�D���m�A��,>��YK����u=3I��j�L���?2?�ye��?�Ȟ�p���s��>k\����@�=��������Y���~U�����:�����)?��>7�?,�J?�E��WDE���)��C,�1˾A�y>H�>9��>�ɾ>�'���G��$v�<þ$ 3��}�<ŀ>�U?�yM?�q?��7�pm(�s����Z�(�����k>#R�=F˅>�m�����+�5%:�O�f�D���튾��
��^;��,? j�>��>�ш?B��>1��!������D�=���9���>�b?��>�kc>�}N��@�i��>��K?G3?���>����6���x� >�/?��>��?�n�>r�����T�)9|��Ʉ�����==�w?-�h�h,���=�tG?����*>���=�yA�����þ��`���`�>(��<�i�>��þ�]���M��m���8?���>����/�b��>*�1?���>GZW>1Ʌ?�^�>Ʋ��2g=`�
?b_0?��B?y�_?.�?V�&>��D� �ѽ��έ�<7J>=�J>�=2h=h��� �� �>�n�0=�P=U���۰�7��<֧��hF����/=�UC>S����=��ȾS#-��.��7�wj���&"��_���흾�2������=M=�n����:�ľ�M��/��?;�@��ƾ����,����b���#�M�>�ӹ��[B=P�{�u�A���%����������ceD�h/m�D���*W4?���N�ѿ;��������8?EA?0��?3�:~��{��>N�=�>w���K
��kƿcf��-4.?���>L�����E>Z��>zLM>.�=�� ?gu*�K�ھ�$B=��%?�6?\3?�[����ݿk,���PC>P��?�h@�A?&�(�w���K=��>,�	?�'A>�2�Kp�^����}�>��?̄�?ۃ8=��V�.ܼ[Kf?�h<��F�t����=W!�=�U=�<�#�H>��>����C�T�޽��4>9��>��%����\���<5�Y>�׽�^��=Մ?{\��f���/��T���U>��T?Q*�>�:�=��,?a7H�!}Ͽ�\�j*a?�0�?��?Z�(??ڿ��ؚ>��ܾ�M?RD6?���>�d&�&�t����=j.ἄ���H��0&V����=���>��>Y�,�����O�BQ��.��=��R�ƿ��$�}��]=s�ݺ�[���罽�����T�M#��fo�U���h=��=r�Q>�k�>:$W>�3Z>�gW?i�k?PN�>�~>:佪���ξj���H�����˥����F�wR�˩߾}�	�������ɾ�|N�N�s>-�]�� ��x�'��P�� K����>���=�ױ���>�=~����c��]����=j7ܽ�ܾ�I�[��㤰?kn<?Cɑ��#U��V��%R=��O���b?;Wս����l	��uA�<Y8�=*�=���>]��=�z��N=��ZZ���6??1L��-8I�
7>���F�^=t�"?�d?�ʴ=���>��%?�[����D>��T>T �>r��>�FA><ỾU���"?}W?�Qѽ�T��?`>5瑾]t]���C=�T>�K�4Be<�f�>E��<�%��Ve;�N��=e�P?Z�}>E7 �{`��Z��������=.��?�#?�a�>��}?Q�x?�V7>�n����K��j!�_"���Z?9�R?�m>�-�⃥��ž $.?�KZ?�a>.������ �ȃ����>���?�h?H�b;�f�n����Z����+?t��?ɮ`�����]z��z��M�?܀?���=Y¹�*V?�?b>;<a�������{��ڀ�?g�@{��?^y���R{���=tV�>ҏ>*"ѽRJ��/g*��񉾖L�G��>^���kl9�%��C}�|!?$�,?.l>�^L��������=��h�?��?����g<���:�k��z��E��<GΫ=1G�X�"�2��!8��ƾ)�
��o���n��Ɇ>TK@���8��>ƒ8��5⿃@Ͽ+օ�0�Ͼ�p���?*M�>1�ɽ�s��U�j���t��G�жH�1�����>�>�&��*����:{��M:�!���8�>�����>��F��|��x"��yi�#��>��>&�>���&2��W͘?J���̿	��$����S?}�?�<�?t?,�<�mm��M{��U��wF?��n?��]?��u��\��2n���d?2[���\�s_C�&HP�&��=liU?t3?{o�u.��'�>?��>�o>y.(�3̿�욿��MD�?`��?���3�>���?��C?����Ya����,�B�<�����?��5>uB�Η+���M��G�u�C?�
Q?O�.�2_�]�_?+�a�N�p���-���ƽ�ۡ> �0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>]H_���u>����:�
i	>���?�~�?Qj?���� ����U>
�}?��>z�~?�c9>}��>6��=K����:�>t�:>�\�#?+c?��?N�5>�K�+Y7��MB�f`3�MIҾ?���|>vpb?��=?@�,>�鎽�wQ�Q6������z6�?��u�8�������a>[\H>�c>�1�����?�p�%�ؿ�i���p'�~54?ù�>O�?[��صt�|���;_?�z�>�6��+���%��)C�S��?�G�?�?R�׾kK̼F>�>�H�> սh���������7>0�B?* ��D����o��>���?�@�ծ?$i���?Jy��	��P_�����>����=��6?�Ծ��i>(S??��=�u�S�����]���>;��?=�?f��>�+d?�Zf�	�5��z��/��>]U@?�o,?�A�;�Ͼ� �>�q?���O��M����@?l�@�@p�J?	����hֿ����SN��L���9��=���=چ2>�ٽ@_�=��7=��8��=�����=w�> �d>!q>6(O>{a;>��)>���M�!�r��Y���R�C�������Z�@��Xv�Uz��3�������?���3ýy���Q�2&�&?`���=I�V?-@Q?��m?��?�r�%O>�*���) =\��>�M=$�y>�?,?d�G?[�)?�f�=|���<b�@�~�����E��h��>:>�>[��>~Y�>-����Q>�uB>��>��>#�B=���<�;e=�W>��>��>���>�:d>F	�[�ο�s����r�A긼pė���?6t̾D�d�╿zھ��׼uOg>ڥM?Wͼ�^��Y����Ds?	 �$Q����	4�=�&?v�v?��>o�z�a��ȟ�=�S<���a��=H��]����I)��ƭ>bF&?�f>�u>��3��b8�d�P��t��n|>[06?S�~O9���u�z�H��_ݾ�PM>V��>G�D��k����E��ti��8{=/y:?�?�L���ذ���u�E��UOR>�.\>�E=o~�=XM>83c�}�ƽH��p.=E��=3�^>�?;3>�p>��>�C��[U�����>�c�>�]�>I38?4sB?�4!>?�<9�Ľ�/߽�&>�Ĵ>e�>�K�>�)��=��=��>l�N>2�=�*H��?���߽'�>~O��?N��J��[�=o3�l��=z��;5���=�����=Ȗ~?À��刿�0{��umD?�/?0�=��E<Y�"������B����?��@Ck�?q�	�£V���?�?�?;��Z��=K��>�٫>-ξ��L�ճ?��Ž�͢�k�	��#�AR�?C�?'0�h͋��l�PC> d%?��Ӿch�>�x�AZ��8����u���#=��>�8H?tV����O�3>�|v
?�?�^򾪩����ȿ|v����>C�?q��??�m��A��l@�܂�>��?+gY?~ni>�g۾�`Z�<��>V�@?�R?��>y9���'�d�?�޶?���?V�I>ۏ?�	s?���>�.��H�/�e���������=48T<Gv�>'I>+Ⱦs�C�&#��Ѓ��?�j��V���|>@�'=���>�l��ٷ��,�=ʱ������1���>��~>iO>��>���>6[�>Oأ>���<?Z�������K?���?-���2n��N�<W��=)�^��&?�I4?k[�|�Ͼ�ը>�\?k?�[?d�>=��P>��G迿7~��H��<��K>*4�>�H�>�$���FK>��Ծ�4D�cp�>�ϗ>�����?ھ�,��]S��GB�>�e!?���>�Ү=��?��?���>m��>M�N�����Ub�	?��*?��?5��?�8?zʾx� ��͓�	|��%�G�m�J>z?�+?p�g>`˅�iV�c��=MF��C4<g�x?j.n?yӎ�K!
?��?�U6?0~9?v"�>��Y�B��S��Cv���!?�1�w�A�J3&�/���?�1?���>�"��.ֽB�ռ���,j����?!\?�6&?���Ga���¾eb�<n�#�¸l�-�;��B���>�>/���ǡ�=k�>Ұ=�$m��T6�3�b<ׯ�=���>v��=:7�`����<?�j��.���O�=g�O��# ��>`;�=S*��;�l?LC,�,�W�Aס�[됿��!�u;�?#��?���?!Z��4c�O�;?��?��Y?�>Qnݾʾ(]�l������f��@�=�JY>h��>kw��U���b���Z��7�>/7���?�=�>X?�?F?�?>��=t¾�:�gZԾ1~2�}b�Fr�.5��e��������ZP��,�(�`;	���D��m=v%��߈>���>\u*=Ҭ>s��>�J��bE>�">��d>죧>�t�>Տj>Ñ�=���`�=9FR?ܳ��u�'��^辺���k�A?�Hd?���>�Kg��u��܇�L�?���?lo�?C�u>��h�[1+�R?�`�>8#��`
?5�;=�����<i8��`��F�������>
׽�:�o�L��mf��O
?�'?;�� �̾�Pֽ�Ђ��)�8�?T�=?�M�� 6�V:\��?���I�,���?-�������=eY��L���xd��@��K�����>D�%?��?��a��f���:���1jG�qJ�>^1?:/�>��>�N>�����1�l��sѾ��x�;F�>�E�?�Y�>�GI?�:?~EO?UL?`$�>�K�>T �����>��4<�#�>K�>�07?�-?�h0?�?9R*?�\^>����W��q�־5W??R�?:?��?D䄾��ɽ1���4×��Py��Z��l�=���<K��bᆽ�T8=��P>��?�I��Z3����%b>�h-?��>|�>�҇��7y�г:=ʦ�>n�?'��>�E��:7s��7����>[�?�����=�U1>���=6y��+�9���=̻j��j�=�����:��,�;��=lh�=rQ>:פ�:��B;��:��=N ?�q?Ҋ�>�؈>@ޅ��. ����#�=��X>��T>�>*�ؾ܂������-g��D{>a��?z�?	f=��=�|�=�P���c���l꾾�<�?/	#?�T?=�?`b=?ҿ"?'S>6��|G��UZ���O��CJ?e(,?{�>V���ʾ�먿[3���?C�?�Fa�����)��4¾��ӽ�/>�Q/��>~�S�����C���t����Fp��j��? ��?6\A���6��G�ɳ��?���<�C?(H�>�A�>�.�>`�)��:h�;��0�;>��>�R?ɣ�>�L?~My?s�\?�D>q�8�M}������L�>�>�&A?� �?�
�?eTu?(�>6>��0� ؾ}�뾇��Ė��n���o!R=�7a>|��>8��>�Ʀ>�W�=�ڽ����B����=� ^>�|�>>�>a2�>1v{>�<��^?s��=jvþ㬾�����@@��w�>�?ok�?��u?�1�=���(6��w�"�Ӽk>���?���?SE?���� v?>�޽���Ҿ߬�>�r
?��>{��U�5>�t�>�6���~�>*�s;^��4���#*>�??H�W?e&�8�ſ*.q�Zp�:5��C�n<D5���Le�y��\��ġ=ӱ��Y��b��Q�Z�R��1������͜��Oz�>�>ؙ�=�p�=4��=���<򳽼Eq�<�G=(��<��=�nq��pn<q7������Ɔ��~���d<�hM=F�)W���?��-?�b�>w-n?��>[�����/�ų�>z�����>��G>#��M�Ѿ�< �4���ս'̂�ї�7g{�&���7O>��_NJ<�� >�9�=��;;w�=z��1+�=$c,<+u<>XE>�C�=���<�+I=g��=���=a�w?G$���H���pP�p���:?�O�>҄�=9þ-A?�C5>���������K'~?y{�?�a�?��	?�2l�b��>�������ز�=<(��\�)>˞�=Z1(��ѷ>�7I>�����j������?O�@�2<?"����	Ͽ�b8>�f7>1,>�R�L>1�h	\���a��:[��q!?�%;�_̾%!�>�:�=��޾��ƾ�A/=!E6>%�a=P��"\�x�=��{�p�8=�@k=>��C>�Ӻ=�ï����=ڳH=���=O�O>m��b�7�jh*��7=���=��b>@w%>�k�>��>�~?�i?��>�DB����Rr����>��=�$�>c<�;V.>= k>�I3?@x:?D�;?X��>��>�W�>I�>��/���h�v�־%�¾+�>�l�?M��?��>�Gv=�t罖�,�	+;�4����=?Z�T?���>X�H>�U����9Y&���.�!����m4��+=�mr��QU�R���Hm�2�㽲�=�p�>���>��>8Ty>�9>��N>��>��>�6�<yp�=%ጻ���<� �����=(�����<�vż̗���u&�;�+�+�����;\��;E�]<Z��;n�=��>%;>7��>�tX>����*�[>�1\�QVg���=����&:-�,�@�e�J�F�+�z����L�=� >h��7��ja?� >� >z��? �i?+6��͜�'�뾲1��:����x�P��<�E���츾��X���h�gwS������>�>�
�>Q�q>��,�z�?�f=�۾�"3�ǃ�>����&	�F�
��9p�(���Ѓ���g�wJ��ujE?����8��=$�{?�"I?u�?�G�>���ܢھ[w,>޺��A:=qE�Ju�㢽-�?9�&?�=�>E�LeC�Y�ƾ��ƽ1�>�U8��qO�_t��53���v��{����>L���QӾ��0�Y`��V����_@�r�7��>8ZP?�)�?.�a�@����LN�rh�m4��5�?ye?��>k�?�?rӔ��0𾗐��id�=�Bs?i��?��?E��=��/=&e#�H6�>\�?��?���?e�d?VL��w�>Wk���>��w���=��>���=��=eG?@�?.?M������cm�5$꾘Yq�C�q<���=�(�>'H�>k�}>���=��<A6�=Ǧ�>\�>6K�>��`> ��>��>��ɾWV��?#U>N�>�;?�h\>��@<����8#	�o�K�(0j��R�{� =)n���!��c�ؽ��8�Ѯh����>:�¿3V�?��>��B��/?/	�;/�WX>��0>�얽��?n�5>�>�r�>m&�>�4�=�n�>��9>GCӾ�>���Sc!��-C�T�R��Ѿ��z>8���L&����	���~6I��k���d�Vj��-��4==��Ͻ<�G�?������k�j�)�k���ؕ?�V�>�6?�܌� ��,�>y��>dč>,H������ƍ�2iᾎ�?U��?�j>#�>�fP?�f?R�>���c�a��j�1�;�S�d���U����-zy��M��6��bU?C�m?$m>?}�W=�v>�v?�.��>�����>j�)��1�\�=���>J걾��[�V�ƾJþ��4��-W>x�y?U�?5A?8�f��_��6�>H>9?���>�+s?�T,?<@?X��uc?����G$�>���>��?�R?ܻe?�A>+<����&��i>Bm��v�C�� ����8������<�x�>�۽3֒��}���mh��,��ν��=jRB>�Tż�Oɽ�� ����=҃�>��^?���>ñ�>e�<?+�	��8� ���,?.{U=K���^l��T���1����>^3i?�J�?"@U?��Z>��J�1jB��x>'�s>�)>�<k>��>
y�_�Q�iQ7=͂!>Gh9>�t�=�:H�!�z��s�������=�%>��>���>�S�1IY>Y�^��]k�Arb>�E�w0���,��y,"�zu�ށ���>�+F?��?۹�=$��0Q�e�n�!�#?�5?�%1?ӆ�?��>Ԟ;i8;���i�[∾�>��G�����Ԟ����y�B�6�m�w�I>L�澿Ю�'�>q�.����3��X��·�+Ұ�����PE=�����ξ��<���>���>�����"��}���¾���p?޸O�R�þ*�˾����D��>�2^=Q`?UM��Ͻ]�-��-��q[W>[D�>w>w�w� ���*R�������>i�D?�t_? �?9���Er�C������'���e��]?���>�?�xA>��=���d�̕c��TE����>9��>����G�松�
#�m��>E�?� >�Y?�R?ɋ
?��_?�{)?d5?F-�>�P��C���!B&?,H�?��=�gҽ�.U��8��-F����>~)?֙A��,�>c"?�f??�&?+.Q?��?>�* ��Y?�ť�>���>�@X���l�_>�J?�ش>�Y?A|�?I?>p�4�<���V���U��=% >G�3?]�#?E�?�Ϸ>S��>s����i<R��>�lN?<�{?{Jv?���=]�?wy�>w��>&�'=Ra�>;L�>hk?4gM?(�?��\?�>	�	<���}��Rs�u}����_<�,��mX=.��zu:���q��]<=N�	���m�d��;G�@�էǼ����AD<��>c�`>�G;���3>O'ž�HӾĆ=�n=���d@�%�6<�e1>ь�>��?C�>ք��'`�d�>z�>���:�?��?_?бT�}P�r�����8����>��]?Vb�=v"p�cC���ރ�Q�R;M�Z?yMh?�y!�=E���/`?s�W?���z.�lLže������P�E?-)?@�q��>Ma�?xkz?�?�9���6q�����nxd��C�r�=�3�>����s�)��>�J?kz>p;>c��<����u�}ۮ�(U?�P�?���?�5x?O�=zYt�0ȿ�������U^?p��>�餾"?~ ��VоfC������!���a:���虾���}��Nh���G�	Q�=��?�+h?uu?MA`?�	
�`y_�@6_�9l���RT� V ������@���>���@��Pq�O������p���g=h9e�l�I�ղ?��,?gq�
K�>�ٕ�����Y��D>m"��Ag������J�G�k�=Ƽ��)LW��#��a�*?�$�>T�>��:?��D1��3���:�����Vd>��>R�>f��>WLj��떾*Yڽo�ϾB�s����xEz>�<`?<iN?�sk?��	��M2�>������P��z��fXR>��>�J�>��M����#+���=�2%o��[
�S펾�}���=A�1?g(z>���>�&�?�+?K��������2���;ͫ�>�)c?��>�=�>�������~�>�/h?��>�m�> S��G�!��8}�'H��&
�>;Ӱ>�@?d>��-�oV�V���?��M7����=��g?�р�=�[�s�}>�P?��g�И*=N֠>�P��"�����u�2�D�=4?#�U=a
2>W�Ⱦ�� �~As�����#�*?�
?-u��&���r>r� ?�w�>ƹ�>�z�?1�>�J��w���E�?O\?��I?X�@?���>1��=6>��^�ʽ�&��M>=���>F�U>YBl=�c�=h��^%[��b��</=E��=�#	�l~Ƚ�V_<�4Ӽ��<�;�<N&3>%�濨8?�X6���@�v8�|���\|�ܙ^�3Fq�%�����������Q�=}W��=�3(��2��Q#¾�0�����?M.@�־��ľW����_{��-�X1 >�~J��� ��ό����Py���'�$�R���D�C�+�V�/bu���%?���j�ڿY+���׾ �?���>�#T?�)���%.�	d�W�>��>����	�5%��xƿ���@�f?���>�? ���;�ԃ#?5�=��>�?��W��y���E��T�>e�j?���>^��H�ӿ*@���>�9��?�"@�|A??�(�N���*V=5��>W�	?��?>=1��>���`�>7�?���?m�M=�W��o
�ue?(r<[�F���ܻ1�=�=c`=����wJ>yf�>�i�LA��ܽy�4>�υ>o�"�J���^�v��<K�]>H�ս�\��5Մ?'{\��f���/��T���T>��T?�*�>�:�=��,?H7H�Z}Ͽ�\��*a?�0�?��?5�(?ۿ��ؚ>��ܾ��M?cD6?���>�d&��t����=G5�ˉ��}���&V����=K��>7�>��,�֋���O��J��b��=��ƼƿX�$��z�{=��ں�t[��罢�����T�`!��}ao��}�I�h=��=߆Q>d�>aW>�&Z>uhW?��k?@I�> q>�N�ц���ξ�-�4A�����������壾LE��߾��	�������ɾ%BJ��3>�S�\Ǐ�q�/�R�W�:$E���>{�>�����t=��}i�����GP�G��=z�e�dw�W�:�mς����?�qQ?���[@T�)!�Sx�=���O%E?7��'�ݞ�����=��=̶=h˴>i)=�����#���V���0?��?.��fَ�"�%>x��}�<��+?��>P�;`�>2�&?S$��w����[>#>I�>KO�>/I>�����zڽ?ӁS?���A���g�>����C�s�d��=rz	>�A6����^M>���<������V�E�z����<��R?���>.�r��K�W����}*�Dc?b�?���>0�x?ģa?]��=q��!e\�-���(���<?��[?�5>��<���1�̾'�=?Łw?p�~=���
�.�F���N~�>���?�;??��ѼYu�q����!��1?ty?k����Q�����u���P>dC?�7?Z�b�E��>��1?�4��y��0c��_�X��Q�?��?��?'�N�dې�d�=��%?W6?�'���(�)ʾ7M>>�%@?�&��Z���E9���M���?V�?�i!?��AC�_��=B���3\�?8�?SȪ�$�g<\��xl�xs��m��<p�=A��"�@��P8�j�ƾ��
�����Y���ҳ�>�Q@��+��>�Q8�20�PEϿ�W�Ͼ��p���?듪>�CȽ�o����j�Cu�ŪG���H�<�����><�>*N���n��E�z���:��`���<�>\�����>�&J��s��M��ׁO<�2�>3�>�)�>�好Ӹ��sӘ?����#ο�!�����b�T?�&�?��?�>?d<�<~^k�4 {�.�B�XF?do?�:^?<̼^)\���U�k�j?�]���O`�l�4��DE���T>�3?�G�>�-�oL|=�B>+��>�l>2/�j�Ŀiض��������?���?Pn꾊��>Y��?qp+?�g�87��QV���*�!�,EA?�2>����y�!��2=��ƒ�T�
?�|0?D\�U.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>gH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?˙�>RW{?���=/�>L �=�lӾ	���k�>>���=�슽x�?j�T?	3�>�G>����U8��mR�I���ᾲb?�x��>�Tn?��B?�=>Է�����p��"��C������]��PW��E���D>$H1>�(>Rv��Zо[8,?�>�V�޿����5C���0?�M�>78?t�Q���z߽��?z�>(�C�}d���i���]�ZV�?��?~Y�>����%>���=�H�>��(>�#��,\=/:���~U>p�{?}鲾�ԡ�^�[��]�>��?%�@���?چ��?�[�ž����������y9+�8>��<?��
���(>�t�>2��=�o��,���Mz�
v�>z+�?�/�?���>��`?O�l�l!,���'=�9�>�EK?�+?e	��1��e)�>0�?��5�/���E񾅽M?ib
@�}@>pi?�����ֿJ����M��XU��j��=P>�f`>��6�G=c���0��$&��3�>���>�{�>�z�>\�6>f~>�Z>�6���%�֗��Z��� <���+���S�v��<����	��c��h�ξ����Ľ�����T��e5��
��\��=-{U?�R?6�o?�� ?(�q�"�>�V��%�=q $�d��=]Æ>M2?��L?��*?k�=���/td���������5�����>�CJ>��>!�>�4�>a,���:H>��=>3�>�� >��*=v�8�3=s�M>|�>��>w~�>.�<>��K>�|����ͿQ�K���=m`�'!�?�����5�����]�{�%�<�Y>6?G��=�/��3'ܿ��ÿw)B?\d�����f®��>lw�>�?�ut>�{��w�k�ī��Müyu��������k����"�M�>�g'?<�f>�u>d�3�`h8��P�2t���S|>�36?>EG9��u���H�[ݾ�LM>%ž>%7D��l�������Cni�nx{==v:?�?�&���䰾b�u��?��\TR>�9\>�I= q�=�KM>r�c���ƽsH��U.=g��=��^>��?���=���=i`�>4ָ�@&r�泥>�g>�f�>/�c?.*1?��"�@�Y�� n��|>#@	?�_�>��=�&H��0�=F��>o8�>`~ܼ����G ��Z��QG>�9ͽ��T�ZIM���H���]����=��=�A����<�r�B=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�#�>J�޲��wt���Ou��70=���>MG?�u�;~���K�;[?��?����S��YCɿ�7w���>$1�?�Q�?��m�펙��5;��b�>'T�?�.[?��o>=7۾ԏa��N�>�B?LsO?o�>�3�����?��?���?a@J>�+�?��s?e�>QC��//�#��_ɋ�̵�=��;,Z�>��>�����_E��s������6aj�[z��c>(�%=|h�>�a��I��>��=s���������\�;۶>2n>PZG>8�>"G ?v��>�F�>�=������	����K?���?��;n�zD�<3˜=R�^��(?�@4?��[��Ͼ�Ѩ>�\?���?�[?3`�>���r@���鿿�v��GP�<�K>�'�>�O�>�D��F?K>T�Ծ*D��o�>MǗ>����@?ھ�6������8�>�_!?A��>��=��?L�>���>���>��]�v�����:�V?8k ?]�?�{?]�0?��߾�	������7����G�O�`>I|X?�?K��>�����s��[=<��X��r�?Ȝb?N���3>?9I�?��(?W�`?�R�>�������BJ���=b�!?>���A�xJ&�c	��v?�C?���>�C��sֽUHռD���m���?A!\?�3&?P��+a���¾�:�<�J#��T�;]�;�[D���>^�>�}��Rv�=Y>���=Im�1T6�Ef<K��=�|�>��=:7��n��і3?�kg��bb��y>��j�%�^���>��>�
u����?�6�K&i��ꏿ�퍿�����?W��?xϕ?1L��h{g�%�a?,��?��?�6 ?Cc(�N��U���[;��UྀE#��Ņ>���>{���sQe��X��$ɼ��ǔ��B�=ç{�5?�>��?��h?\�>}Y�>Ri�11H�������G�Z����'���2��|�#hϾf�f��@���������½#��>�\��1Y'>0��>���=f�j>���>8o��.�d>��5>���=�kl>H��>V��=�Q>ao�=�,W�8JR?)���B'�2��r����@?J�b?^��>=Io������ ?�E�?pŜ?~�u>��h���+�i�?�5�>N����	?�IH=���j��<�B��t�����t��0�>�VӽB�9���L���h���
?ܿ?� ���ʾ�@׽��p���F,�?X�/?��F���7��]���U���M�p�.<��|��ϙ����lzj�Zȗ��h����p��+F>��'?��?{�پ@.������s�,6�}u�>�6?�G�>]�?Yh~>�Oݾ�5���]�l �����Х�>�Na?86�>�H?�;?#N?��N?a��>�v�>Ԋ���E�>K�麉��>jV�>i�8?˞.?t�2?�?��)?d�_> ���t����ܾp?�n?�(?&� ?WZ?���k��#o�7'ü5v��Y���=ѕ�<\R�UU}���7=�Z>�e%?CTJ�VU���.��=��>�tA<�^�>�����x�Mn�>!?�,+?�=;??���5��r�8��9�=Iց?0߼ +���|R> q>�+�;�����1=��*=H~�m !�">���<�f���|=/��>���X�ý<��=��3=%u�>��?���>�D�>YC��\� �ȵ�@g�=Y>� S>�>Dپ�}��#$����g�%]y>�v�?3z�?(�f=��=;��=�|��sU�����a���<��<��?�J#?}WT?���?��=?qi#?6�>>*��L��&^�������?5:,?�>�'���ɾ�a��gJ4�F�?	�?��`����/�&�����>н�>84.���~�)��ݏC�/.9)���ژ�З�?�<�?�{F���6��l羫Z��������D?�J�>���>���>��*�Nf��x���;>�&�>��P?ɰ�>��E?��?�gQ?Ș#>5�;��ά�^����=&�C> ,E?_ks?ª�?u;p?Fy�>��=��B�^�Ծ��Ծh�)�z��kMi�S��=@_A>Hs�>�3�>�g�>���=�%߽S����:k��=�]�=e>�>:�>C��>��}>Ō}<I�T?.>�Ǿ��ʽ?jɾ������>R��?���?"}?v	?���K�:��Ƀ�NeV>���?9j�?9�:?4u��rj>kný���G�ؽ[�a>�>lD�>�0o�Z?[>�)�>��M>�Hi>Y���s�m���;P�<�
?gEX?�ny�H�ſq�Ln��[��Ld�<����c��喽Uu[�A�=>�h�vũ��[�vџ����������%��Z�z��d�>�σ=�=S(�=%��<�ƼV�<�PK=�<��=��k���y<��4���лv�����%�`<rI=lO컦���D�?�sW?|�>�bO?Z��>g��=��
�>�PL�3�>:\=@8���ʾ	��=�o(ཊHs�Ǯ���4��Eٞ��H;>�!��K63=��=��D=�p�c�N>�J>><�==m�;�9L=4��>
s>��(:�=��>.�>l6w?򝁿尝�2Q����y�:?�A�>[��=��ƾ�@?��>>E5��䔹�
f�� ?���?�T�?H�?�ui�Y�>���������ΐ=���$82>���=��2�*��>��J>ʆ��G��38��d2�?��@@�??������Ͽ�k/>c�7>�2>�R�х1�
w\��ub�O�Z���!?XG;�AV̾_1�>��=F�޾6Uƾ��.=d/6>q�`=8��+?\�)�=qB{��<=��k=�̉>X�C>p=�=Z诽	�=X�I=O��=��O>}��Zw8�#�+���3=(��=��b>�&>���>�"?�*?�V?�m�>%Uv�t�ξ-V��S�>�!>g��>:F-=�6>���>b�)?��"?WF?�Ҹ>/� >�>�>�b�>ʙ@���T��پ-�ƾ��Q>P�?a"v?9�>�s�=gB�}v�o�%��q4�g�F?��K?W��>�I>���R4��<*��.�Xg2<��~=�><l��E����̼H��O}��]9,>���>���>��>�1>�q=k�2>uH�>߄�=u�<�[�<SEN��2Q�t�eǡ=CQ�=�4=G!��"�<S�i=�G&�m����S;A�;��<�?�=�>dK�>f�>© ? �t>��$��h/>����!����<i�ľ�9&��E�2~�md�v=���>;Cg>���s`���}$?�B>:�>J��?���?:�=+�Ǿ�ZJ�V\���,��ՠ�j�����=Fݤ��vR��Q���FS�f8ɾ�.�>�p�>< �>6l>h�+�~(@�4U^=8ྙ�3�0�>ʐ��&���p�n�B?�� ���Ii������D?G凿:?�=I�~?��H?��?;`�>vZ����־�4>��~�h&�<y+�;hs��r��Me?�[%?��>7��n+D��!ȾƼ�q�>�C��sO�����X1�p98�쳾4��>�Ѧ���Ͼ�1�1K��`Վ��D���o�Qܺ>��O?�ޭ?X�_��с�`N�M������?�Mg?�۞>�<?��?����H뾷}�Vj�=8^p?k]�?+%�?��>G�Y=���d�>9z ?��?��?�h?�c�[t�>���Ǹ >�I���O�=��=�;�=Q��=G�	?��?q$?矽�l��뾙�|�o�K�<�̴=
'�>N��>��`>���=��=�Ҩ=%�O>�͛>�!�>�a>��>Gl�>c$��Z���=?5{>�"�>�(?�&�>�b=�&�
n��)39�\�c� c���L �����:=	 ���<���;U$�>������?^x�>�J1�,#?˴�g��l�Y>�^>c.׼8�>�*�=�*>S�`>�C�>�[�=��>��#>c7ȾM�>�C���/��=��G����%L�>v2���]'��f�L�޽���<���^���j�b���E���.�J�?H����o�b �H
��?�>^��>h +?�~s�|��}��=��?'ȏ>��������������?G�?Jp^>�B�>�cW??�%�`�(� �X���u�%PA�1�e���`�ܵ��\���{]�O���^?Q�w?��@?)�j<��t>e0�?�i$��Ô�Q�>L�-��Q:��q<=�<�>q�����^�9�о��ľ���ѿG>(Jo?J�?�c?��T�о׳n>i)A?)?(�{?��J?�g*?��3�?5��V�>г�>�R?�?	aG?��3>Q�N>lU-���=
h;�`\��G!�}��=���<�F�=�[>wP�Щ���1<�&<7}=��=q� >�Hu=�=O�M<��ؽ��=li�>�c?���>��n>r-<?�1�$�2��\��L�)?��z<�퍾�����}���t�#>�sc?��?�DV?��P>QJ���S��%>B/�>6_>��=>�׫>z��=��U�=�>��>c�=g)�M�x��o�l ��j)�<a;>e�>�7�>a���0>J��� qh��Q^>�Q�b&��}�]�ZH�=1���~�F��>	�K?�D? і=�㾨N����e��(?ri;?G�K?DR�?�p�=ݐԾ�\>���K�Q� �4��>��%;}�괠�+���A�8���<;��k>�q��>5��6��>PuS�{���|��p��oeݾ�0�1��2��>���]���4	>��=�eȾB�&�D��á��0e?U��=MѾk��	�ľ�>r�>Pc�>bj���y����"�{%�=�j�>*�E>�������A�$<�D7�>��F?Z`?<փ?�O���Rp��p@�����b��F
���?܇�>V�
?g�@>��=�����s�A(e�^G��W�>��>ĳ�e�F�&N��lb�Ï"����>Y�?�>҂
?MhS?�t?�\^?Q,?r�?숐>�e���3���A&?3��?�=>�Խ��T�t 9�BF�t��>i�)?	�B�޹�>H�?�?��&?�Q?̵?P�>�� ��C@����>zY�>��W��b��2�_>��J?皳>k=Y?�ԃ?��=>R�5��颾�֩��U�=�>x�2?�5#?T�?	��>���>�桾xw�=�w�>3�b?�?|�o?�e�=��?'�2>TE�>�/�=��>��>��? �O?��s?�K?���>�R�<ᬽo���op��L�0�W;vH3< u=f����-r�Ǌ"����<���;H	��Fy��/���4J�������;��>�Br>�\��lc0>e�þ�����2A>�?��o���T��K	<�a�=��>��?�'�>\Z"����=s��>V��>i�8�'?&H?B?��㷋sb��Eܾ�\M����>�A?��=�%m�b���q!u�KWs=�[n?��^?�YV��!���b?�^? ��H�<�b�þ2}b�=U���O?�
?��G�F�>�~?=r?���>%3f�
Kn�R���Fb��6k�A�=v��>fg���d��o�>�y7?B�>��b>x��=a�۾ǭw�%����?�ތ?��?�?�&*>!�n��4�]��1H��c^?�t�>v#���"?���v�Ͼ�\�����D+⾵��k���N���~��7�$�x׃��׽�!�=�?�s? Gq?��_?�� �p�c��:^�N	���WV��%�O'���E��#E�˂C�?�n��Q�����$���G=Ho���A����?
�#?������>�l��� ��;)G>f+���$	�F�=]Q��X!==�z=(d��(��t��C� ?���>ѡ�>3>?~_� �<�7+8�cp:�Mj߾P/>��>:ӂ>��>��<4���N���Ѵ�W�y�5r�1_s>�e?UL?��m?��_;/�ۀ�n��GDW�$��CH>A�>G��>)mS�^T�b�'��|@�OCs�a��\����P��>T=��1?�>`C�>*Ֆ?��?^z����`�w�	�,���N<�?�>(j?��>1E�>FؽDh#����>$�d?�
?�`�>Q �����\c�>���߫>���>�?��.>!ĺ,�/��͓�ۈ���IR��:|=�p?R���Ͻ㌬>�aR?x�ýx��=�w>�����5�/u��r���>�?�k���sH>�Ꞿ8��]a|�j���O)?�J?�撾O�*��6~>I$"?)��>�.�>�0�?3*�>oþ��F�ư?P�^?�AJ?{SA?\J�>Z�=� ���<Ƚ��&���,=���>��Z>m'm=��=����r\�_y�,�D=Xw�=��μ�S����<n��v�J<��<��3>�}ֿͪ#������+��� ��1�<���0Q��,�yrw���ܾ;��O��,�/�Ώ��E����C�>\�Q�^a�?�� @ �����m��;��r��'�h>�B7�#;�>N^��Ei��C�����xQ���O�ndx�x�W�)�'?�����ǿ-����>ܾ ?m? ?Φy?>���"��8�	� >x\�<^b��9�����ο������^?}��>�������>���>��X>�Mq>A
���䞾���<�?r�-?��>ȏr���ɿҊ��-��<���?��@��A?�(�F�UU=���>&�?��<>��.��J�/���Qa�>/��?�g�?�B=��W�LK�݋e?��;�tF��Kӻ���=4�=��=�����J>�>W��s�A�˺޽��6>�̆>�? ������^��3�<�]>˘ؽ�����ӄ?�r\���e���/��O���j>��T?yO�>E�=��,?�H��~Ͽ��\� a?�-�?��?��(?"����՚>��ܾQ{M?b)6?K�>[W&�j�t�e��=E�߼/p����㾡V�׼�==��>�N>�v,�ъ�}O�\җ�S��=���Ϳ�����*�D�O�--m:"`=��[N���ҽ���pOǾ��?�����2[>)�V>��m>��{>�Te>���>�5D?��x?���>��>=H�s=�ٮ�g�þ>�n=��I� c���:���"��}���ɾ�yξ�
�R�$N��Ĳ�E4<�>�d��ܓ�a�(���|���9�П?:>VW����P�'#Z��A��sp��R�꼂�����Ӿh�9��=i���?�S?|��Q�F� ������Dͽ�E?���ȾR���j
>�=btR=xm�>�6[<��G�?��]�78?-�?��������r�>�5s�,��<�D?���>��<�	�>�?@�+p[� �w��c�;�ލ>���>h�>a���5 �+�?k=?v���:���ϱ>���r����>>��ɾ/*>��>5s.��!��d�;�U7^=#�=N�W?b��>^'�����r����B����<��y?�?��>��k?CBB?< <ۤ����T�!���=}kP?�Kg?�!>7�j���̾~���3?��b?��U>ۺd�!��w*����@�?�m?�O?�[̼��{��S������5?�iy?�`��������r��YC�>��"?��?��=��>|zf?>�$��?���������<P�?���?��?�؞=����>�1?��.?�h��������Lt��d�=W�?�o���ؓ����� �;B?��?Y?��8�Vcþà�=�ٕ��Z�?{�?s����Dg<J���l��n��ǀ�<�Ϋ=���D"������7���ƾ��
�
����߿����>?Z@�U�*�>D8�O6�TϿ"���[о�Sq���?R��>F�Ƚ����'�j��Pu�S�G�1�H�ܥ��ը�>-�>s���*��$�x�7�k �ʢ�>��߼���>�]S��"��짾M��<���>���>���>�>�������?���Ϳ�`��4��3V?��?�Ɇ?�?X�<YM�-f���;O�EH?�w?�OZ?32�u
G��VB��j?�B��$`���4��)E���T>�$3?9
�>�S-����=�	>6+�>Z�>F�.�ŃĿ�϶�t���mצ?8u�?qi���>���?�g+?/C�,���n��<�*�.�,EA?��1>[����r!��=�����:�
?x'0?����]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?Ե�� #�g6%?�>d����8Ǿ��<���>�(�>*N>bH_���u>����:�i	>���?�~�?Qj?���� ����U>
�}?��>ή�?�%�>�K?;|�<�˅��<��>>�[�f/���?��i?�'?md>U�l���I�:8n�>I`�,1%��M>�+�>�?�)8?=�>}��{ ��fؾ�0��	٦���t���=ə���z�t �>݁>�8>&`��*�$���-?�A�<M׿���㤾�9d?��?���>ܳ��Z��t5��-�?�C>6H
�:��o닿�48�,Ԥ?Ι�?���>��Ǿ��=��q=U��>m�>�>��f;�2�׾J$�="<V?$�/������gj��6�>��?3@}ܣ?s����?��|���������ؾ���K>
�3?EJ���!>�?��#>��y��謹�Eq�]�>CO�?J{�?.f�>�@`? MU�b_��u>UB�>qF?Ck�>��=�Z�b>4`?��#������
��Ip?u�@v�@m]W?	1����ܿ{)��K���b�[h������݊�z4� R�>-Y>�縼uRҼhJ�=�n�>1��>��>rb5>6>�=�J>�T����#�����Ҏ���1��W���y(��2Ӿq��Ol�s0������̾������Ǽг:=A#M�� Խp�Ἲ���M1f?4J?髑?H?Ԟ̽��=�ǾA�R�<%^��C>g��>C?�aE?�	?���_���Io�����+1��;��6:�>u	>^��>6�>Y5>�Ľtqw>hI�>� >S8�Z
���8����#H�=�}�>a��>��>uC<>��>]ϴ��1��|�h�w��̽�?c����J��1���9��t����h�=7b.?�{>���?пl����2H?j���W)�2�+�T�>��0?�cW?Z�>���3�T��:>w����j�p_>�+ ��l���)��%Q>�l?�f>�u><�3��Q8�o�P�w��r|>,6?�U���I9���u�=�H��JݾG�L>�{�>�cE��i�������i��g|=G^:?͂?�β�X����gu��/����Q>M:\>�=;�=>UM>��d�Ȇƽu�G��.=��=:�^>?�5>��=5ގ>���/w��`�>@�8>�^2>u�\?/�2?�����i��������K�=��>ol>��>�7s����=Q?d�k>(�t���߼4*&�첔�DÄ>��=�Ǌ���˽�RO>�)=����=�o<�o������Hj{=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ\��>�h�z����ሿ&G��֤<�>t3?���뭻����5�0? �?�J�-u���*ȿA[��Mr�>l�?9��?��}v�/�k�e��>�i�?�D�?�W->)/þ�Ͼ<O>%�C?�\?ڲ�>�I�("ݽ'�?���?B<r?L	I>���?u�s?�y�><y��B/���������1}=ET;U��>��>�f���NF�mѓ��k��<�j�e����a>OA#=\-�>k�体+��{��=�ዽ+$����e���>"�p>r�I>���>�� ?�C�>,�>I�=O>���逾���5�K?���?���i2n�xO�<=��^��&?I4?xy[���Ͼ�֨> �\?L?�[?8c�>���O>��Q迿e~��<%�K>4�>�H�>@%���FK>��Ծi4D�p�>�ϗ>�񣼧?ھm,��k)���B�>�e!?��>VϮ=T� ?Ր#?߉j>m�>�ZE��6����E���>���>+5?��~?e�?�߹�#Y3����1⡿/y[���M>}�x?uM?Oƕ>	���M}���*F�&+I�m���a��?�ag?^D��?(-�?�??��A?��e>d��<ؾ�׭����>�!?o�˫A��B&���fj?�:?���>�ݓ��cֽ�ԼV��������?\?n)&?���,a���¾b��<4� �OsX���;�;B���>��>�b���P�=�>>��=7m�#�5�n�i<�R�=�u�>�z�=X	7��$���G:?t�����d���=�q5�u��x�>�؟>��1��HD? ��˜|���8~��[	�#��?�[�?�}�?�D��-U���.?�;i?�u?��?eϕ�Ƚ��t'��ʪ�{ؠ���n�M>^>��?�_|����������ǯ����h�V����>��>z?n}�>��:>��>�@{��Z���#���B���r�R���2�Qx
���05�h�����?9X����>C�Q�?�>�i?�P�>$q>��>r�;�<�>��{>Ii�>�x�> Nj>$�]>���=�V<*Q���KR?������'�v�辖���>3B?�qd?[1�>i�������u�?���?As�?L<v>h��,+�an?�>�>2��Fq
?�T:=�4��8�<�U�����_4����n��>5E׽� :�wM�jmf�qj
?�/?���`�̾�;׽������n=�M�?��(?P�)�$�Q�I�o�>�W�S�[���5h��i����$���p��쏿�^���$����(��l*=&�*?�?����!���%k��?�pef>�>'$�>��>)uI>v�	�u�1�"^�M'������Q�>p[{?KD�>��I?-�;?�yP?�L?��>�q�>���`�>�?�;I��>���>D�9?��-?l#0?fY?7[+?�Oc>���������Mؾ� ?��?�A?�?��?�煾"�ý����0an��py�Y��B!�=��<U9ֽ�/t�N�T=��S>��#?o��B�'����D�:>�~?�Z�>�r?�n���M^�=��?�x�>�X2>�s� �k��Rݾ��>ߤx?�"��z�=,>��=S��<c�u��I>r<<)=��=ci��f��Kw9>�T>���P�;#	�����<��\=I�?Ĩ�>~*>���>��J�Q@߾�-\�ɼ��Y�b>��}��V(������l���؛�C�C�^��>X �?���?��=�^Y>�6����7�ų$�{�3�����k�;��J?�~�>xU7?d��?�`6?Nc?;�K>���
얿ίH��K=�a2?0,?���>�\��Aʾ���%v3�]{?�?��`�T�
�=(�6'þ� ѽR�>۾/�Bu~�n᯿F�C���4�� ��=��?�z�?Y�C��+6��W�뱘�5]����C?d��>��>���>�c)�xg���.�6>#W�>*�Q?)�>_�O?�<{?�[?AT>܋8�������8�c�!>�@?ು?��?�y?aP�>�P>�1*��5ྙn��?�����K���LW=;Z>߂�>��>��>M��=1lȽ�u���>���=�~b>ϴ�>棥>t��>�Pw>D'�<IM?�_~>������ھI���EpսN�k>��?z1n?�T�>���>%Pi�eq��d��`?�Y�?=�?��r?�M��r�=���<渰�{&��y�>:�9>�\z>�X.>�D1>��K> s�>Ln�>�}��>��CB�bB��?j�???o <D)ƿ�1r�?�p�!E���.<<y��+g�����RZ�b��=׃��U��L���KEZ����S����N���\����z�H��>��=S�=j��=���<�¼iS�<ƝF=V�<��=�t��2o<.|6��}������s.	��c<�L=����پ�{?"5E?��.?�;M?�7�>��&>�n�W��>x�:'H�>.�0>�Y =i���=%B��۾�#��h����b��ީM�����d�=����'�>p'�>��^>O)>~�b>f�l�k���M1�������xB=��>	�.>�&X>2�s>d�>�@w?���vd����P���轞�:?���>��=��ƾ��??|B>�6��}����}���~?���?S[�?BT?lsg�E�>f����?��s�=���v0>-�=L�3�w��>��L>����f���*����?I@�x??e����/Ͽ�/>��>���=�++�E@��G�ڻl�!	����,?2[����>�	T>;�W���}
����==�>� ��
9/�+hH=��%��-�<��<Μ�>@�w>IF>� l�G��;Mu�<v�:>�ڨ>�ش= [�<���{�=r��;ސ1>�a>�|�>�`?r�*?��\?K�>u':��aԾ ����q�>4S=��>_g|�O�=|��>�P??V]?�:P?��>|ȶ<o��>�ǣ>c�0�og��������J��=�8�?�Ft?T�>�H>\Ӆ�:@G��n �{�[=��? )?�?|��>����w�N	���>��Ӭ��J��׽��<�S�@�o&e�u�Ҿ�����>��?��?�>�Հ>��;>ru�>�u�>mAE>�:̎m=�M/>�r$;=�=���=������?���ѻ�"U=p�=Vi�=���<&$b��C'���@=y�<�7,>r?�>i�>~��>L��="����!>�?x��b�1jE=�ܾ��4��$K�Rm��ԙ5�g)��>}|>�_�%����'?�^[>��Q>n&�?d�X?B�	>#���-)�����b�9�!�����>���aք�ÁG�a�q�U]z���ԣ�>͜�>�`�>�fk>Jf(�U�<�I7g=��~�0����>v���3N�ʵ��f�����d?����l�K����G?�����G�=}�~?G�I?lƉ?yw�>����/WӾ�>�݊���<	�;�R��Ͻ��?�g$?y-�>��hBD��%̾Ix����>H@I�;�O�<���o�0�����з�7��>����о 3�c������0yB�<r��>ŸO?p�?.b��W���6O�B���U���E?�Xg?�^�>�@?�*?�袽���)D��h�=/�n??��?�5�?��
>a��=B��ڜ�>�F	?��?#z�?T�r?y�;��[�>�
�;�>�&���'�=d�
>Cț=��=�N?! 
?�
?�ޛ��/	�8�{~ﾙ�]���<H�=��>�X�>T�m>���=��]=W��=��^>#��>}ƒ>��i>�Q�>��>�D�a��g/E?��G=$�>�p0?�>�>5ʾ*��<w����ؼ(�C�]3m��B�pЊ=��v�U����f=}j�>C���M�?�K >��)E?��|>����?^�_><���_o�>��6>%,�>���>�\�>��w>}��>�c�>SR��N6�>�+e�M��Pk�C���ץ ��;�p��F8>�m���m���]]��ʾ6M���r��n����V�u�5�T�?l����v���II��2?�e>==U?��T�7.��Z>�?��=� ��T��P�����(�?�@{�>G�W>�J?f(+?�%�oQ��Q�Z�����;�#aZ��:��{�����p������G<-Lt?��z?^�D?[5����>
ia?�L�n �>h��%��sW��F�����>\/Ǿ�)�����s#��a�<��>��w?�u?��?�!��_,ξB]�>k�B?\�?�c�?ylG?n�7?�S�,"4?ɂ=��>�~�>�N?iT?��?x��:LPz�IN3�)�l=;��x|d��A��2��h�:���<��=_�� �=j��=�.�=��J�Q��%�=�N=l�>�2�<���;�58=F��>ۤH?���>
�> +R?U�< *0�_��M�?�ڵ�12ξt���G̾�����
>�vw?��?�U?��=��Z����I%�=��>���=��>^K>�L�������t��lrS�_��=�r=p��fQ���m�`����<�8Y=:�>�Dz>�ዽ�t'>=���N�y�?dc>MpP����g`T��QH���1�Ǧv�[�>�;J?��?���=���̚��(jf��y)?j�;?�#M?ǒ?=^�=A�۾;:�'�L�����>�Y�<X��ա���2;�����j>���GH����{>�������f�m��h�����h�����nȵ=g�#�8����FS��&�=j��=�Ǿ�W3��)��������\?)�>�;$�g�������;�8>���>k�=>�g�0�8��셾U��=>�>�E>㭉�+x���8F�g���9�>*RE?�U_?�j�?e���r���B�0����~����Ǽ��?��>�v?�8B>�í=����j��d��G����>���>^����G��"���(����$�l}�>�/?_C>��?��R?��
?��`?� *?�D?#@�>�䷽ ���A&?Ԉ�?�=U�Խ_�T�A 9�iF����>��)?ܻB�Z��>��?��?&�&?��Q?̵?-�>�� �D@�^��>�X�>��W�mb��R�_>�J?���>=Y?�ԃ?(�=>R�5�u颾�ԩ��O�=�>��2?l5#?9�?`��>��>e����q�=���>�c?'�?��o?��=3�?�2>;��>B��=�t�>"��>?�\O?�s?q�J?�v�>�~�<h7���-���r�L
P����;2jF<�[y=��qu�����E�<0@�;�Ϸ�&8���x�ReD�b�����;���>��r>����&1>x�ľoQ���(A>���0?���\��!�;�(v�=ݍ�>�?�і>I �(2�=�,�>��>�,�'?)H?{\?J�9�eb�(�پ�qH���>� B?Q��=4m�����H�u��Ri=on?mK^?%�W������b?��]?�b�@=���þ�b���龍�O?��
?"�G� �>��~?��q?��>f�;n����nCb���j���=�t�>�W���d�h@�>\�7?gK�>��b>�=6y۾��w��l���?��?Q�?��?�,*>��n�4��0�����V?,��>oj���?�Q�K��2nZ���~������*1������%����,��k��wf���y�=�]?�t�?u�c?�d?����Y�o���\��g��}\�� ��j ���I�P�A��hB�O�k�����b�������;�Q2�\?�T�?z ?:RV����>Dk��*��q���M>fO��"r��r�=S=��=���=��O���%�{nS��?���>�sV> II?��Z�� 7��]:��I�IzѾ��	>��g>J�>I�>ST>�V�;޻�x����>�����^�u>m�c?�K?3�n?���1�	����}!�� 1�R`���C>y'>��> �W����wK&�Pe>���r�8�������	���}=��2?�c�>���>�<�?�?�e	�=���wx�l1�ρ<8�>�i?�?�>��>�IϽ�� ��D�>hi?�K�>#F�>��Y�����W��鮼�\�>]�?�?5?ᗯ>�I�=7F�땿�W��A�L���=ϊ�?Z*���Dн'd�>�N?Č:�P��=��>�Q��	�4�I���C����o<>$�:?�%�=�z>*��&�M��Ly��)꽘X)?/�?0`���q*�I }>$�!?�w�>�>�ă?/Ĝ>�vþ�⏻��?��^?ӢJ?�A?���>�x=غ���zȽ�'&��/=��>�3[>�k=MK�=� ��A[������G=t �=�YܼUt��r<W��|�T<��<�3>��ڿ��A���ྜྷ�}�O�g��]���ڑ�q����6)�#��=���H��O)�BwB�ф����Z�¾�R��h��?X@��t#*�����l����� ��>Մ�Bi�w�����!���T��A;Ŗ���!�\l_�*�x���u�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >YC�<-����뾭����οB�����^?���>��/��p��>ޥ�>�X>�Hq>����螾{1�<��?7�-?��>Ďr�1�ɿc����¤<���?0�@|A?��(�*���V=ζ�>̈́	?��?>(=1��B��!��%t�>3�?K�?��K=��W��]	�ȁe?e�<��F�dݻ&X�=5�=_�=����}J>�'�>y���DA��rܽR�4>��>��!���H�^�W��<K�]>�ս������{?�S�h2�e�5�rHx���>��[?�.!?��L���n?L�/�ڿ`Y�خ]?���?���?E?w�ƾk�>�_���,?�_H?�i�>�?��m�b�3�*>aA�=���=ؙ��M
��
�>3��>U>6�νTM�N-����:��M<���8̿�^ ����ۃ':׆�<��h�v�4��9�<�>��N�����5�"}��lz�=́�=KQ>4�c>�/>a\>J U?�3i?Eö>�u>UZ�앾��N㽭�C���׽m|��8��|P����G߾���L#�L��x·�t1�Hh�=7I�-���1���]�M�G���-?�A�=1�վ5Q�r�<�Ⱦ����WҼ!����D߾)�5�3p�gƕ?#�G?�Ą�oT��[�!������_?�����U�����M�=7 ��u%�p>:��<��徍�4��[��i0?�?�&�� T���)>��n�	=J�+?_� ?E�S<8�>6#?2�2���罌2Z>��5>w�>�"�>l>����i5н�"?^dT?��ｽ����~�>Խ���|��>[=��	>��0���ż
hb>@�n<�T���ϊ�N����c�<WnR?V�>���
��{����qo���j?�u?�-�>��|?�LA?R
;��R�f�����5�=C�T?�:V?B[�=��9 ���q���J/?�]?q�/>�N��2�}_�"澙��>��?iP*?�+��̊�����_(��q9?gQu?7�a��H��P���ꈾ���>�R�>T�>��-�Y�8>�;?�����U!��څ3���?j� @i��?�A<����­=[Q�>Z��>�������'�ﵱ�_�,=zh�>�8��� }��z��@ٽ��@?ѵ�?��?��t������=�ٕ��Z�?o�?7����Eg<[���l��n���|�<�ͫ=��E"�����7�c�ƾ��
����D߿����>8Z@W�_*�>D8�I6�TϿ���[о�Sq�e�?'��>1�Ƚ����+�j��Pu�M�G�#�H�⥌����>��=��q��I��Ʋy�IR8�⪧���>�ֻ�h�>��^�
���^���5�5<z~�>���>��>S�p�����{�?����ο����� �g�M?2�?Za�?�*&?���=0��]���~�:�2(?�f?a�T?t)����2=!�j?�_��lU`��4�sHE��U>�"3?�B�>I�-���|=%>~��>�f>�#/�r�Ŀ�ٶ�'���`��?܉�?�o� ��>i��?vs+?�i�	8���[����*��,��<A?�2>���=�!�;0=�lҒ���
?O~0?�z�h.���_?�ia��to���,�����x%�>�3�yma��.�Ƅ��<e� ț��.w�E�?��?��?K��"�"���%?��>7��%`ɾ��<f3�>�b�>SM>��b���v>C��g�:�&�>xZ�?�j�?YN? 쎿�[��S>�8}?��>��?� P>ph?U�>,�s�����a�.>�μ?"�<��?��m?�3,?���=Iy��]WL���e�}D��
Ҿv K�Du�>��%?Ŵ+?�G�>�)���	��@� ���Ǿhv��q�*�������<P��>�u>ˉ�>����bv��e)?��,��-ܿz{��E��/� ?�->Y��>Ot羡ٸ���R��)b?ɜO>��/�3�������� ��6�?���?P?�'���t�c�K����>���>O�`=u!�.tɾ��C=x9R?o}A��T����[�#�>�9�?<v	@���?<�x���?,���Z��Ԫ���:��ܽ���=9�?uN�8�=~��>��=�[x�ٸ��x�P�>6u�?[��?���>�:^?gi� ;�'T�<��>36w?_�?��G���p�@>ͭ?OD$��?��}�辣�t?�W@�@�n^?�r��w̿,p���T���}��9�>�%.>��>���}�|>�ݔ=]���vV�=X`V>�-�>�QT>q4>��>Q>ITi>6��EZ&�]���s���V��v��e�H���}��3ʂ�ɔ%�c����!��27��5���-��D�?���Խ�{�^��=ҊX?c�P?i�p?[?�[c���>S���F1�<�H,�4��=�!�>�{4?��J?~&?jg=E|���a�R ���䪾������>�J>�
�>���>�M�>�v*:�N> C->kr>���=��<hݹ:��=��P>�װ>���>ֻ�>�I<>��>p����)���Yh��w���̽�?{֝��J�Q&��P$������˞=�3.?>���o8п����H?������R+�B>'�0?�bW?�'>C��'�R�-�>
���j�o�>@ ��El�e\)���P>�K?�i>lJ�>F�*�4@�e�3�/а��?%>]�D?S�ھ�k[�@q�Z�6���پV>���>;�+���'�>̗�C����i��p=��9?{��>d�1ᓾ��/�35��Z�,>w�u>��=��= 2>�����ٽ��C��Qp=2[�=� >??�">��=��>���1_����>�'P>�>��;?!�"?s{����cds�D��>���>�>��=/FL�P��=��>�}>�f���O��dJ�7�H>\\���FR��'��*k=>TS����=ԡ�=�V��D@����<�~?����㈿��$f���lD?�+?5�=ÑF<�"�0 ��I���?b�@ m�?�	���V���?�@�?Q��g��=�|�>�֫>Bξr�L�'�?�ƽ4Ȣ�X�	�D*#��S�?��?��/�rʋ�Pl��3>�^%?ɰӾem�>��:�/J���%��)B���R�[�>��2?3O����S�`����E?;C?�R�v�����ʿ���崣>փ�?dx�?9y��%��Q7u�7��>5@�?ho?��i>>q�-����
�>q�-?U�?®7>�_!�����%?QH�?�<�?hI>K��?ɜs?�g�>B&x�`Y/��5��5����V=�[;_c�>H\>�����fF�kד�6h����j����
�a>�}$=��>�K��2��F>�=��6H���f�2��>�+q>S�I>V�>
� ?�`�>飙>�^=�q���〾������K?Ω�?���Q9n�:��<���=	_�M?R�3?�	a���Ͼݴ�>U�\?��?��Z?3%�>���@��^���\k��	��<DL>k&�>xN�>Gm���K>>�ԾYRD�ۍ�>��>o��ھ�ҁ�&Ȣ��%�>�Y!?�M�>V�=� ?�#?>�j>�%�>7[E�7���E�k��>��>lG?�~?,�?-ι�4Y3�,
���硿v�[��AN>��x?�P?�̕>T�����k�D��H��쒽̘�?jmg?���z?Z.�?-�??1�A?=#f>t��;ؾ%���>��%?�B��1�����J<����>آ?|��>h4&��?����Ž��?�����Z!?4�k?��D?�'վ�U�e��R��<"+���i����6ʪ���>�3>էG=�%,>��P>��=�?����������d�=�?�>��>o�3�_�i��I,?��\������=f�q��jD�T�>�O>�����]?��;���{��*��U���+P���?�Y�?c?�?L����g��=?�#�?�{?��>b���_l߾`ྍ�x�՗z��4��C>�`�>�?���Yѣ�	���ʃ�:�ʽ����)�>��>1�?g� ?�N>���>���3Q'�������W^��I��>8�/�.��z�a?��"�$�4��6¾>r{��M�>Y����>�u
?Uh>��{>���>�m��w�>�Q>(�~>�1�>��V>�(4>�>�;<8/ҽ�KR?�����'�������}2B?�pd??.�>�*i�����5���~?J��?�s�?�Av>�|h��++��m?U>�>����p
?�?:=4k��<�V�����%��0�t��>�E׽�!:��M��nf�sj
?�/?�	����̾�@׽᡾csp=)��?��)?S*���R�p�#>Y��Q�4'�Obm����!0$�4(p�3����5���U���J)��!=$�+?���?/�����w�l���?�^h>
v�>Wŕ>f��>��J>����1���]�Y8'��Y����>��y?��>=�F?�
>?�KP?]fL?�c�>g��>1�����>4�3;���>A��>�z2?�
0?_2?9�?�5,?	�\>���F����:վ��?�X?��?)?u�>�퉾�����@�%�����k�f�x��=w�<}Q�-Z[�	XI=�K>�X?F���8����k>m7?y}�>���>��/���K�<~�>��
?A�>L ��|r��`��Z�>+��?��`�=��)>o��=x��uҺ�S�=����l�=p���u;�N�<됿={��=^>u�v���Б�:�ņ;ii�<q�?_w?y��=n�|>���]%��k�徥��=�{�>�7��o��>�\J�7���`����mx�C�_>�C�?M��?�^�0��=�Z>7�g��Ĕ�1벾�Ƙ�zȽl�>w*?ØA?��X?��3?��??�F\>Z!��،�ا^���=��>� ,?��>�����ʾ�憎ˈ3��?�\?|=a����';)�̏¾� ս �>�Z/�%.~�G���D��K��`��B������?H��?��@�1�6��r辪���A]��;�C?�$�>�W�>��>ؾ)�P�g�E#��4;>���>)R?M��>�L?��{?h�[?��[>�5�	*������Yм�d >hx<?=�?�@�?{?G��>75">��%�k[޾j����t�[J��t"w=��I>��>��>�¦>���='ͽ����&P�?�=p�o>�]�>?�>GK�>Nv>��<��@?�m>ٰ�\
���
��f���)�>��q?� �?=�?�u>,�E�h���/����>i��?h*�?s�i?�<N��=�z�<����]r.��>�>�DZ>�U=��p�����u�<?)��>&z���:��L�9S�<��?E2v?��+=S�ƿ(s���p�薾�A<������d�������R� ��=�<�����S�X[Y�u1������\v��L���tz���>t��=��=���=²<�|ڼ V�<�r(=h�<�?=g||��m<Q�D�E�
x��%�K��eb<�FI=�һ�|���?!6?v�?��v?y��>�)�>�=F=J._�R�?���>%�>�@������q�ȾA?!���b��$Ͼ�Ǎ�b��hW>/����>{�	>��y>�=g[f>� >�0��!e��D]���v=`��=��8>�O>��n=��&>A�w?A	��^/����~��Ss��!Z?+"5>���<;�Ծf]?�%�=�������
�#8u?���?~�?�?�K�d��>O�4��`�=��=>+Fl��ɣ=�>���=ke>
~�>VN�zͨ��L��g��?j	@��B?�>t�{ԿKP>��@>�60>��I��f9�l2�4�r�Z��,E2?�=>�z�ھC�A>7"�==�޾�PҾ��<��>]#��	�S�b�s��A=��c��8=jz�=;��>�z>><��=pr���$�=�)�=0�2>�.>�N:�`v��s�j�m=|<���=�W$>B��=��?�N�>�+.?��Z?��>c�Ω�ә���)�<�ڽ�Wy=�D1��$�=^�*?�T?_H?+�I?�Ȉ>�Jq�X�>�/>��Z��3p��dL����ϣ>�1�?�u�?d��>	���4Eƾ��_@���Ѽ��>x-�>���>�%�>S��NO�x���}*���l7�=U\�<;W�#��=wk��S�*��eN>���>���>ч>�>�=?c=^,)>5�>�%O==xu>!$��l�<)��
1"�zL
>�U>s��{Q=x���F����j;�19=��<L��3N����=��>7V>��>�F�=� ��Dr.>�4����L��ؽ=~�����A�G!d��~�I�.�M�5���A>�CW>����%��0?�MY>�>>�^�?��t?��>����Zվ7��7�d��R�.۷=��>�/>���;��C`�n�M��Ӿ'��>-^�>�k�>��m>��+���>���v=����M5�;��>N����6�����q��5��E ��[di��R���D?�A���T�=��}?�I?gǏ?�%�>�♽HLؾ�-.>d ���o	=Κ��xp��鑽_?�'?�q�>77�s�D��,̾�J��OǷ>&XI�zP�D���,�0�߆�᪷���>��o�о"3��e�������B�-Cr����>��O?��?"Xb��V��^O����؅�O�?�}g?��>�L?�Z?
T��d��Z���60�=��n?[��?U?�?F>ä�=pp����>�4	?���?�9�?R�s?��=�R�>�9�;b� >+����o�={G>�	�=,d�=�N?�H
?�?z1��T�	�>]�S��-c^�7�<�l�=ӓ�>@~�>�Yp>�=��m=���=��\>|~�>��>��b>y��>�u�>� b��m��I�J?�n�;�#�>�?)?u��>��=����y=�Ꮍo��8�.�\� ��$�+®<����j׽u�+��~�>��Ŀ�$�?k5�>�I��3�?��վ������==y>A��[��>B��>���>���>=�>G��>E��><��>���}�X>�cD����FZ��L��OlA��/0=1DF=�`Z���:����<�P@�c$�����/�}��>���q_���%��"�?�?��;�M�_�/t��G�
?��{>��^?�nh�C	潼P�>D?٠�>�����J@���A��J��?K��?��m>z��>��[?�<?tz���+�}|[��w�|/C���d�u�^�H�����~�����h��4`?�}w?�$;?x��<9�y>iy?�~+��g���o>��+�I:�O��<M�>X����{���Ӿ����/��!7O>v�e?-��?��?@3U�7���nv�>��3?�?�P�?�7-?.^?pŶ:�2)?�>1�?7.?��F?c�?㳮>vx[=�"B=�D�<5��=��o�����'�ɽ����5�<��=�M̻�sP���l=9m^����=��>_�=<�=�_	=�oC<�_� 4b=X�H=��>r/K?T5
?�ɢ>��7?��8���0�o���?�Eռ9�r�����i̾�_��fQ>.�n?x	�?��G?u�>CH>�o%9�.�>S�>�X>Ƶm>^,�>t�&��~�@��{Fh=�"Z>�a�=�?������"�Hw�?=���=I�?�l�=� �=��=��3��O����R>�{��;t�� ,�`�8�Op4�<n�����>��`?a�-?��=��ܾ��½G�O�45?I)?��1?�G�?i�N��!��)���H�Y���a />!�>;�󤏿���3�@�I�L����=3LϾ�ϳ�Z� >mѾ��澛Ѓ��t$��:�����\�,�=�;��rվ:��� �=�n�=Pľ�-���������CD?��?>��r��M��W��?>�Px>V^�>(�὚����*9�����i�6=�+�>J\�=�	����V������M�>�DE?�N_?�g�?���s�r�B����J`����Ǽ?�?�_�>@]?OB>�$�=D���7��d�nG�S	�>���>3��[�G�e0��N����$�8��>�-?�>x�?g�R?��
?�`?q*?U<?l�>s9����8B&?���?2�=��Խ2�T�A9��F����>��)?R�B�%��>��?�?�&?��Q?��?��>�� �zB@���>�X�>�W�b����_>J�J?���>�=Y?ԃ?Y�=>��5��뢾�٩��T�=�>a�2?�4#?��?���>y��>H�����=��>3
c?r.�?��o?�y�=A�?Z22>���><�=���>���>?�YO?��s?T�J?y��>>��<�@��6T��#Ks��:P�	��;2xH<��y=����
t�r����<���;�N��R��:�pD�:V�����;�J�>[ri>�꓾B+'>�ž�7���H>-�{��-���ބ���F��O�=��>��?a��>���E��=��>��>R���o)?�o?�t?F�;~La���۾]JP�zu�>j�B?͈�=P�h�s����w�ĉR=�l?��]?4gR�͜����b?I�\?�j���<��-þ�Hn�S���P?��	?�hH�b&�>�o|?,�p?�"�>Ld��{m��<����a��g�*E�=+�>Ԅ�?�d�Z�>�$7?\�>��d>��=��ݾ�w��]��x�?|�?
Z�?�	�?�%>�n��Y߿���EX���4Y?�u�>F�Ծu�3?��Ľ���uj'� �_�ܛľ���#y��s{�����Y�����ד�U=�CB?(�q?��g?��K?��!�q�D���i��~�d?��@ݾ����fB�	D���;�'g��
��K����������{�OMA�H�?�&?��0����>����n�Vʾ�@>����&���=ɷ��;UN=��e=3l�m�.�J��� ?�'�>���>��<?{4Z�hF;�mM1��f7����� 3>�>j0�>��>n�;�!$�p�ؽ_ľ���/�ͽ�dc>�pj?�GI?� g?����0���}�k��� ��ג���J>>)>?��>Y�Z�-�K.+���=�p�(s�ꯜ�P��2#=ۡ0?��>#��>#L�?!��>���ۧ��B���0�W&?;!�>'j?h�>��>2��Bq����>�te?���>�#�>��x�1d*�*�^�^�Ǽiԧ>�[�>)�>*��>T=���U�d돿	���,05�g��=��`?����>&;���>o�0?��:�� ��f�>v�3��!�oV���!���; s?�>1�T>1Xݾ�C'��&��n])?6 ?C�����*��N}>��!?�a�>49�>�(�?�ǜ>�aþ�E(��(?{�^?FmJ?|�A?��>�=gJ���Ƚ¡&�Ć/=�>�Z>�m=���=OH��w\�s����F=�G�=gfҼ�N��ui	<�\��'X<R��<b�3>�&ݿ��k�%֐���˾+���t�i~پ9Y��D�x���s�� ����_�Pti�����{�R���:� �c���������� @�n�?�/��΢�֓��9�Y�.&)�o	7>�?�O�<h2Ͼ����;f�徠ž��PS���e��m�V�'?����ǿ���:ܾE! ?�A ?E�y?��-�"�ɒ8�ҭ >�D�<�'��[�뾢����οJ��� �^?���>��v/��}��>���>�X>~Hq>|���螾�/�<��?)�-?=��>r�r�"�ɿh������<���?'�@��A?��(���0	Z=e��>�{	?�?>X�/����L��a��>�<�?l��?3uD=6�W�e��e?w�A<�F��	�]��=���=8�=�%�
FL>z5�>?K��4@�LD޽��4>�r�>�C��� _���<x�[>|G׽����΀?/�L���Y��#��[q��3<��@?f��>,`_>92Y?/,��>տ��z��\I?��?��?A�A?	 ��Б�>�wݾna0?q^,?�q�>{���QQ��*U>��;��}��G���u�ڄ�=Y�T>��(>2R��:��m|��Ǜ����=d��^Xǿ�� �X ����<�+<L�\���ｧ����\��2���f�&�ݽ7w}=��=��N>{R�>�Q>'uW>�kZ?X�f?�!�>�)>R����y�|�оu���:y�����������w)�0�ݾ ���h�����˾��7��=J�P�����*����f�?�E��V.?�j">�+ƾ�
N���;ʜȾ�ѧ�=b���@����Ѿ�40�!�i�Z��?�@?w���KU�K��0F��y��WoZ?�b�H>�J���B�=�֥���=��>K�=GL羧4�w[R�1�0?�	?���<����(>LP��w=��+?�=�>6�p<�1�>�j%?�F%�y���zN>ϼ">d�>���>��>OE����Խ3?��P?,~ �቟�l�>�;��c�~�^�t=��>o?�?���J�`>��<R���"��T3����|<��X?}d�>s� �~ʾ�7���=���=
�}?��>�$=97z?dހ?Kic�F)�Ybz������>:G?VbO?VM!<˄	=�LѾ����3v�>��?�xX>	�j�	u��{�`9���?M�?.�?����)\������Y�I�q3? �u?$dT��������P��Y�>��>m(?G�7�Kl�>�3C?���-����¿R�5���?D�@g��?���9$(�S�x=j�>H4�>�S�D���M��ر�z%O=���>7����R^�A�� O$�NC?�Az?q�?(z\������=�Օ��T�?��?h��s�c<��#l��Y��݌�<�c�=?3�3	"����(�7�#�ƾ��
�����D��ǔ�>�W@S���$�>#8��0⿖SϿ�	���fо�|q�y�?�^�>[<ɽ������j��Tu���G�p�H�?����p�>E�>\����֍��{�B�<�T�˼K��>1��v�>��Q�ͫ�������m�;�˔>-��>&��>Ǚ�sɹ��H�?)� �wnͿ\���i�"�V? 3�?U��?{�?��;p���&ʃ��J�8*J?��w?}Y\?b#��g��J��wj?�����_���3��C��OP>1�2?�)�>6�-��Z�=Ѝ>3�>e$>"Z/�J�Ŀjc���v��~��?���? �����>���?;�)?hf����汩�ݔ*�E��O�B?��0>;�þ=F�Q�:�rُ���?9�,?��6��xU_?�h}�ѯ���"T�K>S����>��=L���v�>Z��<��R>��N�~��?���?�t�?��1�4���G?y׮>g@�\���!�=?�?��}>�{u>���>���SdR�x՝>F��?N��?�#?LՃ�qP��}����?���>r��?���>�a�>��6>x��Tn�<��]>t��4w��+�&?llm?�-?�b
�۱㾑Ko���d�Y�M���U�y�ߎ�>�:?E�?o��>16c�Ȋ����ٖ0���ɾj���kZ���5��b�>
;�>X�>��?��-����?Mp�9�ؿ j��"p'��54?.��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>A�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji����>�!Ҿ0'��5�g�?1��:��Ѥ�;GO'?��־Z�>`��>ÅY����g���4|j�珠>ܤ�?��?(V�>�ރ?Ӹr��!d�v;j>Z��>d)?�`*?�ua=9q��r>�(�>,M��䄿*�Ⱦ1��?�@[�@��D?���chֿ����=N��&������=���=K�2>�ٽr_�=��7=1�8�?�����=m�>��d>q>�'O>Va;>�)>���6�!�	r��I���L�C�����A�Z�>��;Xv�0z�4��
����?��t4ý�y��	Q�W2&��?`�^��=�Y?[CP?��k?��?�苽0t>����G]��N�;���=�؎>�f5?B`E?��#?�7=����b�a�C��*~��a���+�>�dS>�[�>�O�>ڼ�>gI���=>.�9>��R>h��=Ѹ<Hs��d�c=�1W>�<�>A��>>��>�I<>�>:δ�$0���h��w�V̽�?`���]�J�m1��2;��΢��p�=�`.?[u>X���=п2���E/H?3����&���+�x�>�0?�bW?>�>�����T��1>k��@�j��c>" �g{l���)��Q>�h?�ˋ>D^>��,��1�;;���,}f>��<?©�Oy��?x��A��ʬ���i>���>�T<�qP4�lW���Tj���c���f��J?�X�>`�s�Y�g��Xu������OE>�I><� �4�=͢t>Dx���.<��X�z=�5>�>�'?��+>�B�=u��>㌔��-y�
ߛ>C>�)>�B=?|k?m=�'������x�)�p�j>;��>*U|>�>�S�6��=@�>��X>Ʋ���ę��3�X���zA>󘰽�M�0)���Q=y؏�[W�=K�M=���M�K��<�<Mn{?"����?��)$���q���-?˄.?R��>.֑=�J���r&��`��?c@뭦?�.Ѿ:W�(��>���?�!����>��A?�o->_q����X=?��&�r}
�Zq~�h����?�?|7��Od��b��!K>��>�þNh�>xx��Z�������u���#=L��>�8H?�V����O�h>��v
?�?�^�੤���ȿ6|v����>W�?���?f�m��A���@����>9��?�gY?woi>�g۾9`Z����>л@?�R?�>�9��'���?�޶?֯�?I>%��?�s?:k�>-x��[/�b6��T���6q=�\;?b�>�T>����kfF�Hד�h����j������a>l�$=��>}P��3��T8�=.����G��
�f����>�&q>��I>CT�>6� ?�`�>J��>:c=�x���‾����L�K?V��?���=.n�^k�<.�=̨^��*?�?4?_^�f�Ͼa��>v�\?S��?��Z?U�>n���:���࿿�w���Ĕ<�L>�"�>Q�>�È�L$K>�վ�#D�{e�>l��>Y*���)ھ�&������_P�>{c!?���>M��=�� ?Ƃ#?fj>��>-E��T����E����>Wq�>�8?k`~?T�?Y���W(3��撿ʡ�^�[�T�M>]�x?E?�ҕ>x���Kf��ΛH�%'K�W��v��?g?�l罇�?���?aS??�~A?.�e>�E�Baؾ5l��Ȓ�>�w"? ����A��t%�j!�&�?Q�?'K�>�䁽C��͚�:���B��L?.�\?]�'?W��"Ea�rh����<s�U��3��gܗ;"]��Ϫ>�L&>c�k��Ѹ=P>�k�=�bl�s�<�%�<�c�=n܏>e��=�W:�ѻ�� �,?taE�bփ�h�=�[q�H�D���~>��P>�0��C]?��6�Ucz�VH���ݜ�Y�Y�Ԣ�?��?�m�?@ ��Rqg�<h<?<k�?:?$�>5&���Y��+��s��~�B��ϸ>��>eq,�m�羀飿\h���\����ɽ������>$��>��
?�� ?�;>���>;ᓾ�'�_������Z�j���26���,���>��T%�:���þ�7��0��>�ѐ�L��>�#	?�k>H�|>��>�X����>�IM>��{>���>op\>�X5>�� >��;N�ν�LR?JM���'�E��ɰ�7�A?��d?\j�>3=k�~l����.?[��?���?\w>�6h��-+�n0?���>�'��^�
?~�@=Vm�v�<ղ���6�7G���R�^E�>�ֽ��9�l�L�K�g�3
?
G?\�����̾bٽ�.���0=Z�?�u?��7�A[;���|��`���F�������i��C���%���k�)l���T��>����$2�[����t(?�B�?v�󾗶����qI]��:��h>m��>&��>���>2�+>����73�^q`�C-��������>v�z?R��>QZI?�<?�gP?YcL?�Q�>�>59����>�P�;G~�>���>D�9?��-?�40?�m?)7+?��b>�J��z���Ֆؾ��?��?/,??�?5م���½��pb�4�y�5������=��<X�Խ|�n��0T=,&T>��?�����8��e����e>b=/?���>�m�>H��~������<��>k�	?���>j���
q��K��>�n�?�����<w?'>���=W�|�}��;��=����q�=��ＹnV��Y%<���=���=�kg;k�w_i���Ǻ�|M<�L?2?`>�l�>�&0��˾�F����X>�R>���=�~�>'+Z��ȋ�������v��^�>���?�z�?<�i<Ǟ=��4>.y�������ܾ|,��j,=�$�>� ?�/?�?�<s?S�8?;�4>����Ռ�2|���b���?�!,?=��>U����ʾQ騿�3���?[?�5a�I���;)���¾ǬԽ�>cV/��-~�p���D�$�����B������?޸�?��@�7�6��{������S����C?��>�T�>)�>]�)���g�}��(;>��>�Q?�h�>�3?��|?�]?>^m>S�5�%���Ȕ����O�=�6?�pi?��?sl?�b�>ck>��!�m�Ҿ�x޾1M�T���ju��>�B>v�>9K�>-�>���=��⛻rr]�y�=�z{>��?���>�%?Y�;>�w0=CN?
�>Լ��C4۾।����@>��s?ɡe?{C?2T>�!	�M_l��Q)�1m�>��?U��?>�a?�3'�II�==Zݽ:�ƾ�c��.{�>��J>��V>�C>��`<b��R�>~��>w���-�ĦY�)�I� �$?��J?�7�=,�ȿ'�u���d����l�<쬉�S�a�*����K����=�P���K�����9P�����萾VR��	қ�]v�a?��a=I>�� >�_:�;��8<ok=*3�<�w=�#.��<��*��8t�؋��}����<�wA=���= ���`?�r?j�?�|o?"�N>M�>�}D=Q��g��	?TX�>�2�>��������4��ҧ���Ng��9���N����=���i�5�'r>��r=��;�V>~�>�v�=<��zr`����=�x=��>.Ё=�L�=��>R�m?�/h�G����7�ҘJ��?g>��=�m��P�??ah> N��4��(���q?M��?F��?�?�g9��b�>���Q1����Bo�\[�>4�d>��|����>�d>��V�����fT=�8�?��@ȴF?�g����ȿI>�?>�|>lcR��./��[���{��rU��#?G9�	̾�}>	-�=k�ھ�¾�d+=�->�:=�x��fX��W�=�)����==��B=t�>bI>���=�᤽ut�=5=n�=�lO>w�<h���V�P�1=E��=��Y>�G>Pj?]��>fB?f?���>=���h޾(������=�U>�Ɵ>�a���u��z�>��P?�i?/�P?5Rs>aA��8�>C�]>E�;�f�R#%��¾c��>�w�?I��?\�?{�%>�od���ЩH�V� ���>��?�O?e�>���w��Z�h�/��LԽ:=�0�<�v�u3�<�̺�ez�wwt���=^)�>V��>C��>�6>�>��T>7�>5��=ur�=I">>�p���>>�%h<F�'=�G��K�����=t`q=�B=5I�<��N���U�|S^=����X�;[��=!��>�>�>JV�=3繾o %>$'����J���=����n�A�M�b��{�EV-�4�5�a9>=�U>Ⱦ|�����q?��K>��<>"��?Avq?.�>����p{׾� ��~]��kY��K�=Rd>p�A�^<���`�p�M��ҾM4�>@��>ɲ�>��_>�&���>��E�=��Ծ��5����>?M~�{qm�n�⽹`o�󺥿�ʢ�ْh��}�݇A?ǧ�����=܀?/�A?؎�?�]�>4���Tپ�4>��]���==����H�qi�(?S�#?�\�>T���G��;�x�;�c�>�i�����mqR�T�n���R��)�>Tਾ����dZ=�k�}��q���l�чҾ���>9�Y?�?ce�L���ݪݾ2�žU2߾K�?A�l?W�t>G�?��>t�<���fm;�1�5>�3{?�U�?%�?{� >J�=S���[��>�y	?<��?�e�?%�r?Aq?�ev�>�S;T>�1���&�=�>��=t��=LB?M
?د
?=����	���𾸤�e^���<��=v��>Q׉>{�s>��=X=�X�=�a\>%��>B��>h�f>�>�ވ>h_�����[)?�Bu=�3�>?��:>x�=��������r)��6H��ǽl�X��`*�O=~8��=�w�>i�>d���e�?�>��Ծz?����F�+��V>+e>�㽽Dr�>F0>�`>*��>%�>��>��>J�G>C&�����=Gvg���b���w�g���*v7��9��[���ҽe0����>��Њ��Ѿ ��;�|��/��O$g�����.�?�o�=�V[��gA��w��{�>{~�>A 1?� ��fp���8�=Ч>��^>�w��ᐿ�͐�.z��?��?�d>�5�>:W?�&?�.��x1��[�'7w��B�drd���_�Xō�ƻ��x�	�����X`?b�x?1�??<��x>�\�?�s%�����\�>�X-�J�:�L�9=��>�>��H�\�+�оH�¾;���E>��n?���?�/?ЭV�&nC��~i>�C?O�(?�r?*�*?p+0?�뽟�(?i�=�<?J	?a1+?mY?7��>v�=���='SD9�!�<Ioֽ�Ћ��[4�s
����S���5=���<|�>��9=�Vb=��<����z�4��<F ��Hu<�â<B~�=Ϊ�=��>��S?v�>&��>UP6?�0��`�A���從�?���<��X�⋚��N¾���6�#>`�q?��?�QG?V�=u�;�D��[n
>5x�>=�/>V}>|��>2���sU"�^�=@'>8b[>���=Ev�������lď���=�>ʍ?�L=��Y=���>1���A��!}>�\���/�� �1>��7�@/4�/�e�(L�>�N?=�>?{�^>��پ�R�|�J�,GP??��v?��?�/�=�^�x�f H���ʾ��?�C>�7��ē������"�7὘�k>��+�>o�2_�> ����Ӿ�y� �R������v۾�<�ɞ��Ͼn�c�ڸ�=@Ѵ=����a2����tw����T?��<>�ߐ��`�����^��=��O>ߎ�>�H�<uwƽ'�)��:ξ�)��d�>
�>
���y�>��H �9G�>YCE?�7_?_�?�����s���B�����Q��ͨǼ�?h�>�_?OB> �=���_(��d�	G���>5R�>����G��������$��U�>)?U�>��?ٺR?��
?��`?�#*?�E?�*�>g����A&?ˇ�?�=�Խ��T���8��F���>.�)?\�B�ӹ�>	�?߹?��&?ԅQ?;�?��>�� �GC@����>
X�>Q�W��b��'�_>�J?l��>�@Y?�Ճ?�>>τ5�k碾۩�k4�=�>��2?5#?T�?C��>�$?a�w�!�=���>]�W?j��?ηr?��X>��>�,>�?؟3>�<3>"�}>���>%K?�J�?˭{?*�>�p�`B���T���W��,L������<�S���f�5���9=i�=e�6=�⽰��K6���$���ż�g�>`�M>�����=>0Ѿ ���[>0A�5 ���Vr��!g��x�='��>D�?�ע>(���u=倴>���>D���,?:�?�?��;��a�߇��h�ȼ>�??�>B�\�򚗿<�{�7�<Mh?ՍZ?l�5��D�b?�]?�r�"�<�r�þ��c��q���O?��
?P�G�v��>-�~?V�q?+��>��e��6n�i%���>b�
cj�D��=���>���d�
c�>��7?��>܈b>ŋ�=�a۾�w�����?�?2��?��?�)>��n���k����ӑ���[?-��>橨��v?�F1��kѾb��e������ا��˨�����Yg����!�1����Dҽ�5�=t<?Wju?%�r?{�_?њ �r�d��]�o:}�"S����!��UPF��)D��A�*�m�ɻ������ў�^�*=��x�R�?�ȳ?��,?���O�>*f��X� �Лپ��7>����-���.c=(�}�ںb=8�={�Y��!:�/%����?��>U�>�>?/TW�2S8��'3�g:�ec��$>
ݢ>N�>�>p��;~�$��:㽚;˾[����|꽺}v>�Ec?�K?\Wn?hW �v�1��^���!���.���ekA>m8>�҉>�UV�*/�N&��>���r�(���A���
��u�=�\2?i{�>��>��?ؤ?w\	��J����w���0��`�<���>q%i?�&�>tq�>([ν�� �GG�>)"f?*0�>�b�>�>/�
���T��FV�3q�>���>�:�>��>i�ýs�B�E������z2��7>o�K?-|���@��7x>jo ?����� {=�D�>��ټ�������� Y�8�|>?D?�@�=X�:> ���>��Ѐ���w�IN)?�A?����X�*�P~>�"?܀�>>�>�-�?B�>Zqþ~�s�ի?^�^?d?J?�MA?�,�>�4=�߱��DȽt�&�L�,=�s�>��Z>{m=�|�=r���J\��Q�#�D=Ϲ�=�μԝ����<!ڴ���J<���<��3>�5�3,F�o��o�n����m��~�{]�]�5�� +����04[��y���M���޽�'�ᛏ�zG������h�?��?�={���e̔�!�����[�>�3���ҽ�����t�0!��PB��:s��o �G]c�k*���}u�R�'?�����ǿ찡��:ܾ8! ?�A ?8�y?��9�"���8�� >yD�<�*��|�뾦����οO�����^?���>��k/����>���>*�X>�Hq>����螾�2�<��?2�-?��>��r�'�ɿc����¤<���?+�@�vA?�B(��,쾹SY=���>B�	?��@>G0��O�߰��=�>V�?���?PD=lX���	�b�e?m�><��F�ZA��w��=Ť=�j=j��k�I>c��>Z��'A���ܽ7|4>m�>s�����F)_�E��<��Z>��׽%��I�?��T��gD���*��@���=b"d?���>�p+>-4Q?H�4�R#ҿB�R��vV?^ �?t"�?߾%?��ؾzԀ>h㾂�&?�?C�>�j;�s�s�82M>t�_=}s'>=����4g��`>���>���EH�͡��P�(�L��/>n����ƿ�B(����}*#�f�<��-���'��4��Ö�凞�C�0�� ����<���=]�U>tHu>��m>�u[>�Y?Q)f?��>�T�><�#��p���˾�F��PE��}Ͻ������H��ѐ��^뾰�پ������{���Sʾ�Q=�|��=s�Q������� ���b�j�F��.?�%>r˾��M�b�*<O=ʾɧ���-��l����̾#�1�l/n��Ο?SB?�ⅿPW�������*U����W?B�������� �=7h���#=��>�n�=���m3�CeS�Q0?%+?�m��m����5>r���re=&�(?7�>H���6�>n]$?�C9����">��>�б>h�>i">�ݯ����_�?��H?���S ����>��at�e{R=t�	>Y�)��ץ�B\[>=�f�톣��Q����˽��K<?VV?���>pZ'�����Ɗ�T��M�U= v?I�?���>�}m?��C?_ר<�S��oW��M��=�fY?>je?D2�=�g�VʾX����<2?�Pd?�F>�j�"�x�(���?�Yo?�?b���S~�T���3?cwv?�e[�w������J�O�>�d�>��>M"9�N��>H�??����)��ƿ���4����?j�@�G�?��z<��]�=b?��>��H�UA���X��
U��* [=�.�>m^��
�p���_~)�tc2?�d�?T��>,��a0� ��=�Օ��W�??�?�����e<���ll��e����<=r ��I"����7�j�ƾV�
�餜�c������>TY@8i��-�>4/8�n3�RϿ'���YоNOq���?�s�>��Ƚ%���}�j�Ru���G���H���>���=����۩ľ/π���L��D��}��>� �<4Av>�������]ﾐ�4=�C�>��>̽�>=���Sy��rr�?�u9�]�ƿ۲��ǣ��j?�ϡ?�y?/�?��������M����<�c?ج�?�*�?h�8��l���]=�j?3_��FU`���4�7HE��U>�"3?�B�>P�-���|=�>���>�f>�#/�w�Ŀsٶ�����`��?���?�o���>N��?Hs+?�i��7���[����*�L�+��<A?�2>�����!�0=�sҒ�a�
?�}0?�{�W.�6;Z?Yx������|wo��j��>�>Cئ�u��<�V�>V�ɾ����H�� �4��S�?��?!�?[옾z���KL?Ʈ>!>ؾ����x�<>��?E*#?�M.>��=$?�>�?�������8>{�?�-�?�;/?�H��	����^)��ه?Ս>�:�?z�M>��>1�$>
7E�7��<�{�=A�����=M�?h�~?
��>�횽����s`���G��,A�ê
���N��Z�>�L?�`,?ZB�>�Ĳ�'_�͸�]���h����-�=J��Q���.�����>;>���=Q*��������?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji�$	?���U���W~����3�7�/��=��7?��#�z>���>~c�=�vv�������s�e��>�6�?u�?���>��l?C�o��C�.H1=]L�>ϑk?�p?W}q�D�ŪB>�? ��o����4��0f?��
@:t@6�^?sܢ�D=տz��(ޤ��{;ͺ'=sdF=�>�F�J9�=�==�!&<~�ɼ� >Z'�>��Y>��U>>�;>�P:>�p>������ �h��°��Z'I��n"��$	��w^��E�}�y���	��¾a�Ծ���:���I���F�Z��!��~h�=HUT?-�O?�n?�2?�j��Q�>�t���6=�� �V6s=���>Nz1?!lL?��)?>O�=RZ��J�c�����'��J�����>��J>e��>M�>�c�>����.H>)L?>�:�>��>ˠ(=鵢;��.=4�R>�l�>�&�>���>�C<>�>,ϴ��1���h�Zw��̽�?O���#�J��1���9��v���j�=(b.?{>����>п3����2H?���� )�׹+�H�>��0?ZcW?��>
����T�P:>M��?�j��`>o* ��~l���)�&Q>2l?�i>��v>�3���5�O�K��0��@�t>S6?����H6���t���E�-u׾��S>�A�>�¼/�#�|$���rz�e�e�a.;=��:?��?���2����c|�������L>�}W>%r'=+��=�qM>�3���n�>�V{'=O��=��T>�?�[G>��=�N�>�u�:2;��ߨ>��R>��><1?��)?&��<�v��ß���M����F>9Z�>���>�		>�z_����=�#�>ؙR>0q��Q����Uj;��D>ϲH�ŮL��|���<�=�P��u�=um׼yHW��d���=�rw?Gj���^��,	꾱���[�G?�[?�W�>�wL>I���h���už��?�:@�
�?H��'[�ݺ�>7G�?m��k�I>8o"?�>"7��=��)?����N���I�{g��Ò?{�?6��-�n��T#��?J>�?��ξOh�>ux��Z�������u�$�#=J��>�8H?�V����O�i>��v
?�?�^�ީ����ȿ6|v����>V�?���?j�m��A���@����>:��?�gY?joi>�g۾7`Z����>ϻ@?�R?�>�9�n�'���?�޶?կ�?�XI>�{�?�7s?�M�>L�v��/�J���`��$��=M{;d�>��>ݎ��BF������`���j�����tb>�#=θ>4%�3"��F��=�����맾�d��@�>��p>�I>rK�>�� ?3j�>[��>�=�捽��������K?���?���)n��3�<!�=J�^��'?�C4?W[���Ͼ�Ш>
�\?���?��Z?:M�>����:���޿�t��0�<��K>�-�>�O�>춈�K><�Ծ/D�2l�>�ԗ>R ��4ھe��C��/H�>�c!?���>���=�� ?��#?�uj>�'�>UE��;���E���>	��>�H?��~?I�?Qй�P3����䡿w�[��(N><�x?�I?)͕>����}���D�>uI�9Ē�䙂?gg?=4���?�*�?/�??��A?[f>����ؾX���O�>��!?���4�A�Z�%�5����?4�?�1�>����ӽ}P�u������?��[?hT%?�t��a�w���lv�<�D��ͺ��;��-�~�>�*>����I�=`�>o�=�Lj�t5���s<N��=v��>��=��5�X葽�+?���t�����=Y�r�>$E��o�>#�L>�T��g|_?��;�V|��������\S����?�o�?ɇ�?
��Tg���=?�?o�?8N�>Ѡ���C�*"�~W���h��#��.l>��>P�����ţ�F7���0��t6�\����>���>�?f� ?��?>��>$�����%����n��<�\�Tj�#�5�v-�
�b��'��	��)����w��/ؚ>Kɋ�3;�>?(a>��u>{`�>��ӻ��>�	V>��>��>�@^>��5>�,�=��P<�{ս��Q?��Ⱦ�]%�~�������;?�,g?�,�>q�{�O���1���?���?(S�?���>o.c��*�Q?��?���r?�n=bp��{0��O�����&䪶����>�����
3��M��~���t?�?��(��|ľȩ��̬��/�=���?��$?�a-�@�S��to��TV�ʸK���N�v�h����5�!��Dm�V���]=��� ���!.��W�<x-?x׉?) �_����X��Mrh�[�>��n>@U�>Ɛ>˸�>�X5> �\�,��R[�+>*�ۈ�9�>�v?���>�eI?��;?�lP?�tL?N��>Uɨ>�H���[�>�I�;w٠>���>��9?	.?�60?�X?X2+?�=c>����|���̬ؾm$?��?�-?�2?�v?�7����ýku���Z��z�Ǣ��j]�=��<�Uֽ�sp�9V=2ST>�?�MϽ6�~��r]o>e�?���>���>;���9kd�|_�����>�H?cǑ>\I��Z_p�����>F�}?�!�6�0��b4>�R�=��e<?�><u�=����w�.=ħ��+�VZ=��=s!�=��=�{�� �X�/�#;�%����?�#?f�W>⹈>n�!�/YѾ<ܳ�7>�y=Z��=i"�>�k� �{�Pz������bF>_��?���?��<#�+=�&>�Ѕ�k8�����޴Ⱦ�����>-�
?\{H?ń?]�0?��'?��>��r����M��9������>� ,?���>����ʾb�3���?�Z?b8a�ű��;)��¾��Խ��>W/��-~�+��D�Z��������_��?f��?��@�X�6��~�����7X��ےC?�%�>�Y�>��>��)�0�g�5 ��?;>���>�	R?���>T�?4r?��x?M��>�(�t���{񥿃��_�#><�3?�YI?�t?�?���>��B>���v.¾
�ƾ�P��
)���S�>�G=eȣ>M��>7h>���<z�ϽF�8=�<޾ ��=&��>�|�>���>�?]�/>N��;x�9?�LD>E�z���$�-���l��*�><��?Ͳ�?
��?q�+=����+;��,�Bz�>ܘ�?С�?Q�?-�ѽ���=Th����2p�mÕ>��N>[��>���=ip���>��>>?Ƽ&qC�ؔg�9w���:?�a?�I>�ſ�nq���p�����4c<`e��ae�|��1�Z���=<ǘ��G�k���f[�O���=�������Ü��h{�1��>\��=m�=�i�=���<��ɼ�a�<�=J=�܎<,&=yp���m<#H8��{»yx��A�$�|�S<��I=�.����&��c�?�cE?���>�t?��?8>c�B����������?�@?��>��*��| ��>Ͻ������9���1-��v���W���=�V>�$�=�M���=�9�f���R+�_$��#�=��)>���>D5c>��4>|�'>��v?Du���b���R��󽒰8?��>���=;Dľ��>?_Y5>xq��Jɹ�f�
��~?�0�?
|�?yl?��g�pk�>
��b;��R�=E^��+j:>���=�"/�ƹ>�D>^'�"���ާ�)��?�@��A?�����UϿ�3>ú;>]">��Q�6�.��Q��v���Y��!?3g8���ɾ�=�>�ĺ=�~پ������+=�'>,��<i���X�p�=tї�(uf=M�d=�C�>�L>^&�=�7��a��=�?=E��=�$X>��K�'Q	��zܼ��A=�ѿ=�sg>�>�m�>�ۿ>?�iq?>sQ޽U��w����rƎ=��>oĝ�m���^�>�w5?o�Y?��>?P�>��"����>�<�>�}�S�����d��J-?�5�? �?8�?�A��HE��z�d�S�Â���2	?�f?��	?�7�>����2߿:�(��,�_��g =:�[=�H��g�t���U�Y/��9��>篙>���>0�>�q>��T>c�O>5�>-T�=Fi�<�>+u�o�r��\���Ip=�_\<��=>d��8T�$ȇ<>�q�[��Eٿ�*�K~�����;l>h��>�,>�\�>�v�=�7��5��=�=˾�XV����=�z��C�;m�
j�`�����:S�>"E2>[�:�����?��O>���>��?�L�?e���ȭ�q���}��󟨽�-��)����x>Nӽne/��2Y��T����ҹ�>�N�>�>3�l>e�+�Q�>���v=�Ά65�{�>Dŋ�^����q��6��� ���i�i�ʺ)GD?T=���B�=�	~?�uI?ƴ�?���>�虽�ؾ�/>�	��>�=X���p�����?b�&?���>�I�Y�D���ƾ�IF:#�[>#s�ҷd�Mf����L�<�ݼ��?��Ʀ>b@�������?��#q�-a���Z�@ǝ��#�>�*?�p�?o�ʾ}����4� �ݾ(��:`�>WtB?��K>�a?O��>�
`�]���G�o�.>��y?��?���?@�>Y��=i��e%�>�	?ү�?���?ps?Z�>��p�>[;�">���\��=+�	>���=|��=��?��
?c�
?���;�	����\��^��<�=IQ�>BY�>�q>��=�"h=,�=$�[>��>lc�>XJd>Bͣ>�-�>�w�r�����?�{�=+�>#�	?�v�=�gX=�7�뱀=�ܽ�Δ���EP;�s-����`�$� �I=젢<u8�>^g¿DΚ?�6�>�ݾ�.?���}B��<>��d>�A9<-I�>#AT>h[�>�x�>)��>(+�>��>��\>?����zR>*6Ǿ+'���U�7�Y�N�b>��>���i�w� �v���X��s\���p��w��RMN�5����O�?+���oe���E�)ؽ���>��>��-?������]<c?>P��>`N>�?&���U���z��?��?Z-�?�=c>ė�>��V?�?+�h�,��|\�h�x�ǒC���d�>^�Í��N���q	�}����(`?f�x?�|>?.��;o<x>�?�x%�xw���>0�-��[:�*N:==8�>W}��2�b�b�ҾR�ľ���"�E>�Wn?C�?j?�6U������=*>YW:?ݤ0?zut?{�2?K�;?��#?�C/>�?�?��4?�R-?V�	?�02>���=/�\���!=Q����!�ѽ��Ƚ��케�A=I3|=�-��JW<��=���<S���8ؼT{N;�}���ٻ<�3==(X�=ւ�=��>ML?m{�>w�>b):?"╽_�8��aѾaw?q,�<0}�����˾cG�	�=��k?&i�?�4R?�v�=��F�K�.���> ��>HD)>$�o>�e�>�$���n���h���>�5>ԯ^=jp�G��<��A����ż���=|i?��=��$�=�û��e� ��=E�Z���0�=���V�7���q���J�>�#5?5�?��=E&���UB��=��R?!�
?C�|?��?D��=�?�~|S���I��񶾎U?uq�<�%\�=���5���1�Z��M�P>_���U��ݬ>j&C�,��mI�p�|����L����r������$x���(�-�=�C=NB��}F��N��ٻ����5?8��=c����1���Ǿ�כ=mC�>,�> /�=gC^�2:��9���<>���>��X>X���������J�� !��<�>�<E?oB_?�D�?|+��T�r��B�\�������(hƼ�?���>K?�~A>L׭=~±��)�r�d��$G�!��>�>���e�G�Q��?S����$��-�>j:?n>ɚ?p�R??�
?�`?�*?�d?=B�>�������	B&?��?��=9�Խm�T�4�8��F���>�)?��B�>��>�?h�?��&?��Q?D�?j�>� �L@@�̓�><Z�>��W��b����_>��J?w��>�>Y?�Ճ?�=>��5�F뢾n֩�$Y�=,>"�2?�4#?��?y��>~��>С��m�=5o�>;c?��?E�o?j��=�v?�^/>��>~��=%�>�V�>:]?-�O?�s?6J?���>y݅<����V��/Xx�6�`���;H�B<��y=���Hs��
�_��<VSL;�|������.�1�=��c����;�
�>��a>�1��y<#>?&¾�˅��B>Ѻ3�ꔗ�f��BLH��O=ώ�>x	?l��>	��4��=C�>�<�>1��(�&?��?j�?��e<�{c���о�RT���>�F?�u>�ai�2����o���>=_~k?%x^?#�T�����#�b?��]?
h�=���þĵb��龌�O?��
?��G��>7�~?a�q?���>��e��9n����Cb�D�j�Wж=!r�>3X�Y�d�t?�>3�7?�O�>��b>�)�=$u۾ �w��q��I?[�?��?���?0**>-�n�4���8���Z?���>�̞�.�?㙨�E�Ӿ�{������{�o���9��Ȫ���~��,�Y䃾|�ӽ&��=��?Ty?Ċs?�D[?�w�ff�,_��P���S�@����<�mrG��4C�wRA��/n��e��=��ŗ��[:=�	Q�Ͱ=�SG�?S�?@J�0\�>����]��*O޾�8>����nϽ@�>rd���_=�Mr=h�w��>�䅌�G�?�rx>��>��C?4�C�ʴ0�_kG���C�����x�=�(�>Οt> \?��>����u��͜�_GT�tS@=�mu>�vb?T.J?�}j?����.�?p��?6!�L�o������=>��> "�>!m^�~�s7'�^B@�p�q��������8���=��/?W#>�|�>w��?2?���te���~���-�?��<�T�>�Fh?���>�׆>��ҽ]��4��>E�`?���>�}�>�I��l��I�z�s�н�|�>)��>.�>�#�>�u-��0]�8Ȓ��:����/�>o>�;H?����K���8v>��3?޸ü���<�>8ͮ��"�Ͼ�:�\W>���>"�=�=>J_���03�5W���؎� +)?���>�t���,��p�>�v%?|V�>Ť>��}?swg>�����y��?5�k?�R?�3D?w�>N�D=�":��Sڽ73.�l(<�Hh>�<$>pO=~+�=t�6�;����|I=�R=��v�p���]��<��j�>�<�W�<�e>��ݿ6�4�3p�����qUþw�"������jT��H��@�����ž�����)i�j�(��/�z���u�� ���N㽽	�?��?�o��u��E嘿���ө��X�>[vq�q�G;�����M��I��H+;a$���G��O�;�[�y_\�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���}¤<���?0�@�yA?5�(�!��{PV=���>��	?�?>Hi1��J�����r\�>�4�?��?�M=-�W�l	��ye?:P<��F���ܻt��=��=��=�����J>,�>��;@A��:ܽn�4>ԅ>{� ��S�P�^�cپ<�|]>��ս����w?TZ���j���4�T���؅>2�}?�>�j��l?�F�[FͿ�#L��lg?���?ju�?�8?�,׾�}�>��վ�{3?x)?�3�>L�S���
0=g��=�5J�(¢���V��K�=�?�.>�:��T-�w���������>8��-ÿ��"����}��='C'�c���A�����<ٜv�[�����.�J�ɽ_%)=��=`>� l>2�H>�c�>�N?�{?���>ǘ>
uȽ���~ݾ�߱�΀{�Z=�W!��C3j�ښ���J��>���J��	��f��U=��ލ=�R� ���2� ���b���F�.�.?�j%>��ʾO�M��I3<�Cʾ%�������Ǧ��X̾4�1��m��?��A?�䅿_�V�O��j?�>&��n�W?�%�;��%��O�=p,����=�>�J�=[�⾌3��sS��`0?	?>S���d���&+>܃��v~.=��,?S' ?��*<��>��#?�j1�l^�-I\>S6>Q��>���>?�>I��(8Խ��?A1U?V���L2����>����0x�
��=��
>�+�;L����Y>�b�;����Θ7��<��k3�< W?C��>1/)�1���6z"��f4=oXx?B?84�>��k?z�B?UD�<P~���T��+��J�= X?��h?�k>lmz�C�ϾX���~�4?/vd?��I>�j��辟).����?8�n?�e?Z����F~�	z�����q%6?�r?ާ_�-U��	���5��z
�>�? ,�>�E,��ƚ>4�B?"������X����3��^�?'�@�W�?���<���8�<�f�>}q�>���0���'�o��W̾
È=�4�>�l�������(�c<���JL?�h�?1�?�A���<
���=�֕��Y�?E�?s���ɏg<����l��n��}��<�ƫ=��S"�7��-�7�>�ƾ6�
� ����￼ޠ�>iY@�N轭#�>�E8�4⿆RϿl���^о/Pq���?w��>¥Ƚ���j�Su��G��H�����[�>S��=�?M�������~��Y3�?d�=ډ�>@@�Z�>�\c�9�ھD���T=|�>��>�^�>��qϲ�Qڌ?0M���)ʿ�����T4�*�N?I"�?x�?@�I?p>7����6������?�b?��6?��ѽL�"�XGҼ$�j?�_��sU`��4�qHE��U>�"3?�B�>Q�-�v�|=�>���>g>�#/�y�Ŀ�ٶ�5���Z��?��?�o���>o��?rs+?�i�8���[����*���+��<A?�2>���C�!�>0=�YҒ���
?K~0?5{�b.��u_?�a��-p�~�,���½2�>��5��c�����&)��Fe��b��8o�E�?���?s��?Ķ�[�!���&?5�>�꓾��Ⱦ9I�<E��>�q�>8V>^|>�
!~>\��* ;���>.��?���?�?Y����n���>`�|?�r�>���?@�>Sw.?���>	U���i�.��>���\�=c�?�Q?
e?K]��Fe���\\�b�D��]�A3���G�O�?>ؘ??1?�֓>t�������ʾ�����H=������="��@�M>U�U>�>�^9��c��?o���ؿ�/���U�u�1?*��>c% ?%����d���Gh?[�>e��ܰ��������B�?���?��?�F�A����=�Ȱ>s�>{ه���PY���>IvD?���:���
k���>Z��?�@�<�?�;j���?޳�2�������2`��䢽3">{� ? wƾ�W>k��>�%|>Zr�6ܫ�(wx�;к>m]�?~^�?tX?�t`?�/u�':���+��ܳ>칂?�B?���W1��}��=��?���N���e�s�g?Ծ
@u�@�[Y?t~��S�޿5���X��6�ξ�e=��<B��=)�-���>y�s=Yh^=l��=�+>/�>RzU>
~D>��>t�>��>=����k�h瞿�N����A�~�!��{�B>��l޾G�����P���x���r����������c��@-�ͨ����=$�T?��R?lp?Ig?�-|��V>�3��N��<�#��=�ņ>�1?�LK?�)?��=I���Qd�1��_���:��v�>�dG>)��>��>�"�>�o�j�D>��8>��z>�t>[y=�R;�-=��S>-)�>G�>4��>�C<>��>Dϴ��1��n�h��
w�E̽0�?y���K�J��1���9��Ӧ���h�=Hb.?|>���?пd����2H?&���z)��+���>{�0?�cW?.�>��c�T�.:>5����j�!`>�+ ��l���)��%Q>tl?��j>�7o>�y2�`�7��QN�'�����y>��1?�����4��-t���G�$.׾�%J>���>��g��.���|�vf���V=��<?<�?����ö��f��M����Q>��c>�t6=�\�=pO>��?�H��
h4�u�]=���=�U>�Q?��,>p�=�ޡ>�t���PK�)_�>�D>8L#>�>?�%?�	���/��j0�@eq>��>���>���=�}L����=9�>v�a>$� �ƌ���w�8{D��VS>�_��S^��$K�u��=������=�W�=����B��*&=R.|?c���^���
��d��I!E?�?5��=���<&(�!Ƨ�8�����?�z@��?���YoT�]q?�ɏ?�������=��>J�>о��;���?�?��8������0�	��?���?"?[�8N����d�Ȑ>��?�Ӿ��>">�����򥂿����^1�:���>)�D?�x���5=6+���?q��>QY�u,�������l���>��?]B�?敆������W����>�?�^c?z
>����g0 ���>6�Y?wP(?��F>���8�;s�1?���?i+�?�VI>2��?�q?��>�M��,-��"��K)���bJ=���;���>@�>����XwF�􆒿�f���l��)� BW>$=ec�>`@۽dE��8e�=��������Nl�C�>�ek>�RD>.g�>�� ?��>��>�=�����w��z|��\�K?Y��?���2n�K�<���=��^�j&?�H4?�g[���Ͼ�Ԩ>��\?4?�[?�c�>I��&>��迿�}����<#�K>�4�>�H�>�'��EGK>�Ծ04D��p�>�ϗ>���?ھT,��|M���B�>�e!?>��>�Ѯ=̙ ?��#?��j>�(�>�`E��9����E�X��>g��>�H?��~?��?:Թ��Z3�����桿ё[��<N>�x?�T?�˕>厏�Y����yE��?I�������?�sg?�Q�4?�1�?��??�A?i(f>����	ؾ³��y�>B�!?S3g�2�h�c�2�����?�� ?d��>k��\���郄��64�v���W*?�u?TC1?G����=�X�"�/�_;&��L��;߇`=���[u<k��=hV���=�:u>�?>{�������G����=W#�>�=>��G���%��5,?s��C��L��=�vn�%nB��J}>�dT>)���]?$D)�d�v��Ы�c���Lfc�m#�?W�?�X�?\ݳ���f�̵;?�a�?��?1��>>ⱾNi�P�z`k�%vq�;?��=>�.�>
|�UK��!��|ª��������N�s}?��>��?�Y�>E^>}+�>盾[.�#AҾڙ����J��;�]�7��*�z�"�kR��D�8�hD��+8ƾLyu�:
�>�I��1�>���>�}>"<Y><A�>��"�u�>��r>��>�E�>D�\>�J/>\�=�Uz�!��L?gվ��-�k�۾HX��8?>�??^,�>���.��sn!��I�>�?\�?4p�>K�'���$�J��>,�-?Z�p�<e?0����o;�:�=��B�|��=�`>��a>���>��S���<�nL8��	2�Σ?h?�=I�Kk��������os=�/�?��(?L�)�6�Q�m�o�k�W���R�'���h��_���$�xKp�����ON��� ��<n(���'=�1*?x�?�"�G��<~��#�j���>�|�e>���>���>�@�>pJ>��	���1���]�t�'�Z������>=�z?���>�0?n�C?�%h?�`P?��V>J�>lR��]�>�Eλ�Ɩ>��>�3?ƅA?�{6?�5&?V�.?�:->��ٽ������̾�D ?Ix ?�!?r��>��>^����&� ꕽj6=��ۣ�IS�=��ݚ�����<X$��?�6>1=?kA��8�2��	Yj>,i7?��>��>v��5k��:L�<i�>��
?�o�>�����q�5�����>%\�?û��z�<�(>N��=� ��E�Q��
�=����H7�=N΂���>��'<�=,��=L,��:�k�:�;H;N�<,~?��
?�p�>�y�>��Ľiy�������>=��=6�K>z�?C�P̃�]���/ri�
�_>h�?& �?2�;�M+=n	>(k��~_����w�ܾ��t�s�}>�2?�tL?Ռ/?��-?9D?~�H>iX���������|����?^!,?��>�����ʾ��3�d�?�Z?Z:a�;��|;)�,�¾�Խ��>!V/��)~�����D��������jy��u��?���?%�@���6��s�-���s[��_�C?n'�>�W�>.�>]�)�E�g�d"�_8;>��>3R?%H�>��?�]?`V?�d>h�*�H�����Tq;�2%���N?��f?;��?]�?[��>z�H>]�)�}�� �i��:�|+�\����=��E>���>���>\+�>��>�z��-�ܽ����.G>�6�>LH?G��>�4�>��b>��%>�%8?�M>�����,�c �I�*��Y�>���?��^?���>OO>�r0�����A���{�>Ǹ�?��?ғ??򫾓S�=GƧ=�a��)�F��U�>v�>��>��	>N?�� �[u2?�:?o@��R:��d��� �z�	?��u?m��;�!ڿJ j�~������J):����8E̾��q��Z>�k�=�H�>P33�M�$����>{ξBJ����>%��_?y>�4%<�P>�Ͻ<r�4�J$�<^g�=�>�Ɏ��b�Xdɽ.�̽�0�H6B�w�������b���ͷ����?�W?ݩh?Y��?��>�R{=��>��@�J"�s�?w�>hB�=r]���B��/���U���߾%-�~(��乩���.=�.���o:>�a>w�n>s����볻6z������b�-���$٭=��@>U&�>��(>F�a>[#>�o?Đ��'Y��q8d��A^���z?���>�N��oc��/?E�j>��q�W���o �"�n?�n�?��?@4?:;!�8�u>���to��x��=)���!.>�=Zj����>��>- 0�'�������?�p@��:?��.�ҿ��0>/pI>�]�=%�J�4��|\��KP�~l;�|i#?H;��|�A��>9�=���pؾT�=�=,>�J�=e`���q^�C׌=�N�픂=͞�=���>z�B>�w�=~���=�$ =�">?�>�x�<6.��c(]�J�b=��=ȕ�>�X1>��>�M�>�^6?�q?���>X|�`���j.ᾚ��=�G9=Н�>�S���>V��>��8?�HU?aBY?&�O>�$=�+�>=�e>��5����4�1������>��?�߄?���>>a������Q���L��-�>��?�h�>j��>	s��O�3�&��F.�C���u�û_]=N.u�F��d���$�YUƽ��=[�>E�>;�>��r>L�5>$P>�(�>^/>g��<��=���l�<�Σ��g�=D�>��F�<F�pl�dz��*X,�z���;f˃;�b<�H< n>?=O:>Y��>�=�D��S��=�j��7@��$>*g���j%�SHO�&�v��@������F�=�9/>����Ok����"?�\>7UC>c�? 8~?�IS>_/뽷��;���HJK�.�%�%m�=Є�=���4F�oq��BY�d�ݾ$��>��>�7�>mn>�+�Ʀ>�*r=�$�^(5��?�>����/*����m"q�kQ�������h�i��M'D?#J���q�=�}?0�I?ҏ?���>@Ք��׾��,>�=�
=��p����?F&?Tm�>�<���D��=Ǿ^֭��Ӳ>dcI��rV������+0�V�!<�+����>A�������ϻ+��;��o���B�^���)̲>$MR?䃶?�>��j��}pS����fxr�(�?�a?�΍>d�?��?oμŅ�P���[s=��p?Vd�?�?�E>���=���*��>�N?��?@y�?@s?H�?�]��>5�����>~�����=/%>F@�=K1�=��?�
?ژ?oS���g	�Y��A��{�_�n=6^�=��>ă�>�qt>>��=�MX=X�=6�Y>q��>�c�>�Dd>��>wȇ>�����;�K�-?�4u=�l>S�?��l>������1|`=���oܽ�����ݽ)��		8��ý��<s�h�0��>��ȿ�Y�?�ݐ>�ɾ��>$x
�aQ�5S>�>H�(��>Vի>&�>q�>��>���>1��>�v�>
 �ur�>:t��
�T�O�E�v�Q{�d�u>*J;�L~���`��ڵ��z�����P� ��.q��T����T�~���M��?֋��O ��[���A�?D>�>��=?�������=��w>8�?n4z>������=i��v~�7�?�_ @E<c>��>1�W?�?�1�u3��uZ�o�u�(A��e��`�7፿����}�
������_?��x?�xA?DW�<j:z>ˢ�?��%�tҏ��)�>z/��';�G7<=R*�>�*���`�m�Ӿ*�þ�4��IF>{�o?0%�?zY?�PV��W�^�>|�A?��??y?�X'?��6?"w/��=?L>+D?�X?��/?��8?��?�gZ>��>�6�H&=吥�#���=����Y޽�S�[�:=��9=Ə�5,��~�<�=Р��P��P��:-���V�<7�=�(E=Hȹ= y�>s�\?j��>�R�>c�7?Xn��T6�J6��h.?7&0=�Uz�-���e3���C��`�>uij?�*�?Z7\?v_a>ɔA���@�#x>Ύ�>M�'>�CZ>�O�>}x��ED���=��>�
>���=�O��9���*	����b��<H� >�?��=���+e>q�����Z�{\Y>�7�dW��c�"�pE��I��U��=�>~�K?L�*?�:�=HB��]:�;��T��W2?�2d?�_?�;�?��D=w��`U��� �IK����>�lz>���'@������ͯB�`�߽�U>�Ӿ�_i>Ԅ�ݭ��<B�C�����V���fd��'}�=�R?��U:�PY�f�H>�.>h4�����ӳ��胡�cy7?Bh>aڣ��˱�%��b��=[f~>�:�>�~�wS��z�T��4޾xЍ�G_�>�X�=\/�C�C�U��]ľ{�>�pK?��d?~��?��p��5r�o�7�fB��A�H��:)��C?ie~>fG�>t䠼iF3>� `��D��w4�`��y? �>O�/�բT�[��#����=��do>�=?Kru>�V/?h�U?%d"?��?�?s�?���>��P<���!�1?p�?ư0>z�!��{F���+��2P��^�>�W?+�~�?s?�qF?�?ZX?JI`?WZ"?�=�M��q�8���>؅>��7�����>��>�Q?��>Ҏ#?��j?tg>���	0�%ђ=�|�>Ð�>�@K?�K�>�5?l�=���>�ڔ���>��>�k?m�w?q�q?�ס=_r�>i�>4y�>�>�:d>�ֶ>� ?��A?�{x?C89?�4�>�|��*�?n��o5n���;R�L=��=;s=�|?��n�������I=z�=�Z���G��s��f�� ��Qh�=@[�>ris>쬕��1>U�ľ�K��?[A>�����̜�(Ɗ���:����=�i�>�?M�>p�#����=��>K�>7���1(?��?A�?@;:�b�';۾�K�Z�>"�A?f��=7�l�ʁ��
v�Pxf=��m?�R^?�vW�(���7�b?�^?��m=��fþ�b����O?�?o�E�'��>�q?9�q?�o�>�Ib��m�؜�Lta��6l�d��=Yz�>��ze���>��7?\��>��a>�\�=N�ھ�Pw�����Q?�͌?yޯ?��?�(>nn���������U^?+��>�ܦ�u"?��4��Ͼ1f��#������թ�໨�>ߒ�᧾�'�v�� �ս�ݾ=�D?Ps?so?��_?����@d�4w^����܁T�}��7����E�ƉE���C� �o��}�hr��-$����M=��:���R�ˇ�?l/?�OO�I0�>9ǽ������@r>�?���$ڽ���>j#+�[�#<e��<򫱽H�������?��>R%�>N???5=�ry.�`.���#��t�U�r=7��>A�>n��>v��=�d��_X�Y�ʾ:�]�����s>�Z^?4<;?��?ɮ�=n\B�`K��ر�`��<!F��١>5�=�YZ���"����i��V6�I�R�.�	�����K�|x�>Q�1?ֵ�=cm~>ݩ�?���>�	�%妾�§���-�  ����=ŭb?裵>�=��Ͻ)7����>�l?�a�>u��>Ǯ���Z!���{�:1ͽ��>4�>ξ�>Co>�-�$�[��b���^���8��l�=eh?�����`�M=�>�R?�S~9��H<��>��x��!�;y�1U(��>�%?�S�=`�<>}�ž�'��M{�F����+?�X?�8*�x�8�j�}>�]?��>&y�>8�?�B�>x����=�$1?y?�GX?�^?2m�><ӹ=��r���~����s=D=`>cX>9a@=�T'=1� ���W�j]�ɏ!�u`U<��h=�H/�IֽOq=����$f��v
>�N�צ[��������M���|�J��+��p��7^�3ݽ�s���U�f�:�)��=����3�����l����)�?jB�?N^��ze}�y���<Y��Ǖ
�>~�>�	��Q,��̿�� #�S���h���&����m!���2�c�k���h� ~'?�����ǿ����&�۾`� ?�? z?��t�"�m�8�$� >��<h󯼲�贚�bϿ;���Z_?ܠ�>~(����1�>Or�>��\>sr>+������$��< �?	�-?~��>b`q�!cɿ�Z����<���?|@��:?�{3�4^�����=��>�x?�S�>q7��:�������>q�?fɑ?x��=�O���{���f?�8<-�7��{�v�>���<���=9�l\%>7��>B�6�k�x�x���,�>]��>�\9��O��`����>��l>�����`�5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�򉤻{���&V�}��=[��>c�>,������O��I��U��=�<�Szſ,H)�=�Fh�{�ֻT-f��Y �Ä�����"k��\�t��(����G=��/>��{>\��>E�>��>��]?��v?���>#�>@������i�ʾl�<ϮK��-�9����.������۾ѽ�>��0�
�;�V3Ͼ�$D�J�_=�~T�6؏���"��`��A���.?w@>N�ξ�,O��U�r�ž�+��yE�<P�|��þ�=6�x�m�
�?ÅE?-:��:�K��(���;�����P?�s���:���"�=������W=��>.�e=�Vݾ�r0���R�;;0?�?d	��3��x�+>���l��<�/+?�?�G<S_�>$%?�*�j}޽��Z>�5>�;�>��>[/>���4�۽L-?ɟT?`�����nT�>�|���D|�
�Q=�3>T�7���:�X>8��<1���F}�yؒ�!�<x(W?#��>T�)����a��R���Y==>�x?5�?�.�>#{k?��B?:ܤ<�g����S���kew=��W?�)i?�> ���R	оK����5?�e?g�N>�ch�����.�U�e$?��n?<_?e���4w}�f��R���n6?�w?R�[���<����g�Fc�>���>&�>��9�⎧>�9?�)�⥕� &���5���?l�@`��?�>S<r�3�w��=��?Ě�>X�mTҾ�u���7��k=Ln?�
����z�� ���,�P12?`׃?�?�>�"��-��+�>���Wh�??̌?f����xm<ʾ@�`�h�-�lX[��.v=�(��=Ʒ��e1D��۾{� �����g��<'%f>h�@��F���>QȽ�!ۿ9�ʿ�y��y�b띾%�? X>�`�2׾���yn���L�Q�.�0�K�zN�>��>��������X�{��q;�@��K�>���C	�>�S�T%��ݙ��q�5<��>Ȯ�>ĵ�>�'���潾�ę?�b��v?ο����)��\�X?�f�?�m�?�r?K�9<�v���{��I��/G?��s?�Z?`%��9]�`�7�x�u?KǾ mp� �a�h�e���>�,W?n?{W/��a��Ɇ��!�>��U;�8�W"����bw�T��?�O�?/־
�?X��?u(?%�K�����E��<���Ek?��=�U��T)�V%�J���ri ?�[?:q~�\r:�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?n�>��?���=k��>�%�=� ���5��E#>�\�=!@�c�?9�M?��>qC�=4�8��/��>F�3R��"���C���>��a?dyL?��a>q���Ѕ-��� �wͽ�L1�-�케~@�l8.�"��I�5>9�=>�>��D�;�Ҿ�C2?.�8�Ǿݿ1������!�?.�>C~&?�!��m���ɡ�X�^?X��>D�\M�������g�I��?|@5�?�����/�=.�=,+�=��v>4
>�Wm�����}=�;-?�Q0�]�|�k3��`}>%��?34@<��?��^��	?���P��Za~����7����=��7?�0���z>���>��=�nv�ܻ��Y�s����>�B�?�{�?��>�l?��o�E�B���1=*M�>��k?�s?Lo��󾆲B>��?(������L��f?
�
@|u@[�^?+��⿝����3���C�����=��P>!�v>K�]��D�=�Z�<������;� @>#-�>���>�@�>�q>���=\�:>���Ŭ ��������*kb�Q� ��pKo��EǾe(��I
����M���J+�_pP�i�;<�ư��I�\l���N�='V?bQ?�p?Aj?�����>~���/=|�(����=":�>�,?dJ?�9+??��=>a��)d�zM��N5������1�>��M>m��>���>��>�7���<7>�DC>��x>ck�=�u�<d���w =9A:>��>}��>���>�;>jg>�˴��*��{�h��Jw��f̽<��?7����J��0���Q�������S�=Bp.?ؙ>���`:п(񭿳:H?I͔���[:+��>ٮ0?%W?S>��T�v�>���ҍj���>t �c�l�v)�	#Q>�J?��E>��e>�n5���6��*P�iɲ�~5i>��3?)��I;;�L~u�X
G�ӻؾ�ZQ>,q�>����龖������X�U�n=R�8?��?�ؖ��K��>.��������G>p�h>�1�<�
�=�L>C ��Hнb�L��SY=%�=o�N>rl?�S>
��=���>�a���N����>dy8>�>>�??��?��!�%������ŝ*���p>��>vsw>��=�uG�^0�=T�>R�b>����q��W���$�0�9>��MR�*AQ�yZ�=a*���t>7�=���_:��2=�~?���(䈿��e���lD?T+?g �=؝F<��"�D ���H��G�?q�@m�?��	�ߢV�B�?�@�?��J��=}�>׫>�ξ�L��?��Ž6Ǣ�ɔ	�,)#�hS�?��?��/�Yʋ�:l��6>�^%?�Ӿ�Q�>���"r������jDB��Ο>EH�>O�}?���~p2�O'v��q�>�2)?<!�+)��!�ʿ}���<?��?��?�A���M���73��,?�?eV?@`�>���!��
�>�uk?|IB?鴭>�f$������?J)�?��?��V>���?2i?���>u-|<K?��5��%y�9#�=���=�X�>Z��>`z���S�/�5�m(U�5���m�>�bg=Ql�>�t�o6��-��=���]�׾�����B?��>@��>��> �?�[?���>�P>�h�<Rn�������ZF?8X�?���7b_��؎=���ֿ����>7�M?����T���>Վk?"�l?ݗT?��?��$�����r+��#.��⾢< *�=w�<?v?��t�.�>/r��9
���Ų=A�=��ѽ���@��?*h�d��>?��=�V>��?a?.��>"�>�}�yϚ�_lC��"�>`��>�t?��o?l"?���l��`��[˟�}�8�ZhZ>XLw?$?d��>����$1���׬=����Yu���G[?B
�?V��=h�2?�Ӕ?��?T�4?���>��=�I�������B>0�!?t����A��W&����u?�+?���>#/��Ӏս�Ѽ���%���?s5\?�Y&?ը�
a�w+þCW�<��!�øQ�c��;�D���>�^>�q��*�=��>���=i�m�S�5���c<V�=>��>ô�=:7��Ŏ�3t-?�s=�,����O=�u��!@����>�f>��¾VZ?�fD�y$~�iӬ�����	i����?"��?���?5=��sf��;?�׈?��?�N�>03��X�ھ�w�64y��^H��B�e��=���>�����4���'���j��!��� y����>���>t2?$	�>%<>zħ>dg��"d�C�+FݾaTQ���&�oE�]��X��8w���$/��������Ӂi����>�,����>�V?l��>�V�>��>P���ʥ>�'5>���>Tuu>���>v�_>�(}=K��<��Z���R?�¾>�(����B찾w�C?��d?�9�>�q�� ��L���Q?�Y�?�5�?r�q>��h��6*���?�o ?YF���
?@IJ=MY��-�;Z���2������"M��=�>>�ٽ��9��M�^�g�˭	?��?ٿL���̾8�0~z�+�=��?��@?�L���Q�5�D�*8@���k�x�Ƚ�YG�4��þ��O{��雿�Ɇ��@n� �2��=Ċ?#�?������뾃�~�m�~�9�f�t�>L�?��>T��>��*>i�*�s Y�<�F�K�&���>����>p�l?X)�>�O?�R6?��S?SSp?�Z>y�>�1����>qP����>��>�K�>h�?)75?��3?��?z�=�U������+��???E&?�1?t'��B����,=�����>����~��<Nϕ=˱�U�A>�a�>�: >Y?Ǚ��8�*����j>{�7?��>$��>����'��8��<��>�
?�F�> �h~r�Qb�W�>���?��=��)>� �=����x�Һ�S�=` ¼��=�
���z;��<���=N �=
s��������:	3�;�^�<ʃ�>��?j�>h�>|��� �y�oz�=�2X>��R>�>?�پ�|��S'��Zh�y�x>Vb�?�r�?��h=��=`�=����ʾ�$���S���3�<�d?+>#?ԖT?�?�=?6:#??~>��}0���P��8����?�3?N�|>��l;�C���m �p�&?{��>e�a��]л>��U�J��C̾=��W�?�o� ��|�
�-�>�l��%�����?�̬?�:5��I0�`�־�r���B��t7r?B��>���>Z?.���g�~�5���=��>��V?kA�>�FZ?�Gc?J�Q?�̕>4=?�¿��4��,`>��>vG\?o�?�w?�'j?J{�>��=>�xI=�־��E8�/=.�	ӑ��S�=��I>�o�>���>��>|�<=����������*>ŏ�>��>L<�>|�>�1J>5c��6�G? ��>nN��_���社{�����<�6�u?햐?��+?=����E�G��3H�>m�?���?�0*?��S����=n
׼�ݶ�6�q��#�>�ع>�6�>��=��E=�M>�
�>���>N�U_��n8�uyM�6�?�F?Q��=����]��Q�� ���΂��2&��M9���pE��3f<9�t="R����&)X���q�OG��v��Ө�6-���y�>! >��>�,>ڷ>�=�=�!�)�8|,���=��(�N��j�;�U]=�j�P�潈��<�����4(Ⱦ��r?g K?��%?�hQ?~�>T�F>����^B�>tv˽t�?a�>��轨]о���E[��E3o�K�̾��¾�`�^��=3�?�l)>�G>8=�=�᝹���=@(=��q=8�c��f�;�Z�=�ȋ=8��= �=��>�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>}y2>>��R�^!1�b�]��'c�]s\�X� ?��9���˾�G�>4r�=�N޾�ľ\[==��7>�En=ls��\���=7�|���A=��t=�d�>m�E>)�=���LB�=�UR=���=0N> �a�"�/���7��X.=�@�=��`>�h$>��>X�?�f0?MTd?TG�>RWn�xϾ���&C�>>��=�j�>���=��A>aK�>��7?4�D?`�K?`i�>�M�=��>���>pu,���m�Z�۱��/�<���??���>�cS<GA����7S>��\Ľ�f?�B1?�X?��>�����*�q
)��޽��<�ޅ<�푾
`�<F�2<1�P������
>ܡ>F��>���>kΊ>�~�=%��=<a�>��(>@���/�@=��<���`��%�y^Q=iJ=@n�=�,9<�K�Ǯ���� �i��%3�ѐ5=�߄���4�4��=���>$E>&��>&��=}���C/>T���C�L�Tѿ=�F���*B�n3d�'F~�P/��X6�M�B>]8X>i~���2����?{�Y>�m?>���?>u?��>^���վbP���Ee��OS�wǸ=/�>�<��v;��W`�X�M��zҾ]��>I�M>4��>(��>�p�&����`>�$��<K�lG?#m���JL�qqν/������R����8�[Ű=�~E?�+u�`�s�ʮ�?�R3?�?"�>Y6��
��Y�>S�%����4 �ܯ^��ц=i�`?�)?j0�>����DQ��˾���y0�>)�F�S�O��ӕ�ŀ0��R�zm��c�>���о	63��������b�B�4�q����>y�O?���?�9`�/��*BO�S������V?�{g?3�>��?9�?]���{�
�z�=�tn?k�?���?Q_>���=�	w��E�>HG	?�u�?O��?$�q?+LA��5�>�׼���$>�LE�nv=�b�=��=^>M4?�O?�7�>:���"�
���	��9�]��;=�S�=��>�x>�T>���=<#�=#��=p�C>��>�t>��x>l8�>ku�>��i�t��
�7?H�$>� >8�(?Ҫ�>pq��-T�lG�>�	7�<_e�Z�/�}�������;��}=ԵO=�QT�?�>m۽�o��?��T>ށ�&q?d��j��=,��=�)�<�I3�6��>T�>�'|=�Q�>��>�2`>պ5>�=�޾k>v>�'�V�5�ǝ1��!;�S�׾8��=hSC�C`2�^�4�	1Ⱦ�\��ڢ�;B�۩g�����;N� Ώ��r�?���\���# ����Ԇ?LG�>\&s?5�ʾ��ɽ�y�>��"?���>�7�tT���,���{ྸ��?M��?};c>6�>��W?��?1��/3��qZ�Ŧu��*A�#e�ֶ`�Dߍ�%����
�vG��r�_?_�x?�vA?
Ԓ<�3z>���?J�%�~֏�?-�>!/�0-;��<=�6�>���T�`�s�ӾC�þ�K�OdF>��o?k#�??V?YHV�x+��"m>>P�??�$?.��?L$? C?|��5�?7Q�=��>��!??d?E�?ƈ?��?> y�>"�#<z+5=򟾽V����������B�vg>�ߨ=�%��e[=
��<L�<�1�;����������Z�m�μ,=��C>�y�>`�[?���>�ϗ>�KK?Ń!�C["������^"? G�<cA��w�s�ھ5�޾�;>EZc?��?�yF?�>�EY��=h���>�^>w�>%g>�v�>B�Ž�U���[;�؟=L^H>/��=E v��Q����$�7��=j�N>���>
�{>;�����(>�!��4#z�e>��Q�E��=�S�̵G�F�1�t�u��a�>�K?^�?���=DR�e���7*f��)?�#<?rDM?��?�Г=~۾��9�)�J�}T���>!�<A	��������b�:�b`�:� t>���S���-�o>#���T���]���Q������@�W�پ��D<��:�����_�`�=��f>L�p��	F����6��� I?�
�=f��1�&����ud>s��>�ϱ=�K�'��<"&��q�k9�m�>Y���E��8��p�(��>���>$qM?uT?b��?�Y4���^��?6�so�8���&�uP?�k> #�>!k>�ҟ=�����_�fQ[���<�*�?�G�>P-��Zi��eԾ��ƾ��-���>л)?_�>m
?�
H?P3%?"�V?�	?��?��>	Ž���DE(?n)�?��=�;�A��%�dCJ��t�>�"@?3���G՘>,?F?�3?��/?4k?���=vX�5	 �M;�>c s>��C�ؾ����>D6?Z�>�d?�?ް�>l.���4��$��!]�=��H=b[3?z�?`�?��>A�q>�Kᾁ9�>�H�>�;�?P�?=]�?��)=��>/7>H�>󱷽�+"?Z?M�f?�_�?��?��3?S5>d�˼�[:����7C=j2=t>�0�<����d�/�X�U-��$s��;�=Mm�;�9���= rV=�������F��>���>m��PK>�Ф����*�>P<=Ko������;�����a=�	g>�&�>�r�>�v�^�x=���>R��>��/��[?��*?,?����k������\,�5E�>"�'?�N<�=i�3R��cqp��v�=o�l?�Ye?�@7���0�a?'�e?�a�C�%���z�a��.��T?%�?�V?����>�J{?h?��>�Nf���f�����y�Z���7��2=�8�>jR��p]��9�>�^*?�	�>�I>&�Y=����q�s��a?�#?��?g�?�g>S�s�p�ۿ��.����_?�n�>J����?1��;־����	���~�Ծ*���㖨��]��g믾�-���y�K�׽�U�=�?�q?ph?��^?y��_��7]��<~�� V���9 ���=���D�#�>�l(u��F�a���zU����=M�i��<D�n��?F)?�	R���>b@������ݾ�T>Y������.�=Jj��k�<�{=��U�+�����V??�>�ϼ>y;?LM�S4:���0� 8�����>9Y�>�,�>\��>zo<	�O�$+���̾�؃�uuý!�>�4n?OH?��|?w�<�[0����M9��=:��1��J�>F��<*"|����}Cj��	
��Yi�
k�N��W!ɾ�<�� ,���>?�,�>�Z�>0��?��3>7d���Fڔ���%�U6�L�>V�N?PDn>�>,�k��	���>n�d?�d�>9��>�bǾX��Ob�'�!����>uN�>�>��F>�1�<�h��@�����m-�K2>s�a?l���'u���>X�T?����9=��>����)�_,�Lb/�#�>�D?��<F>>��Ǿ�������,b���&?K�?B���G�)���>xk?��>t�>>τ?���>s ����<��?�s]?�WI?.�A?7e�>�#'=)�������K+�h0=^��>��U>�
p=c��=��P�S�86�<�"�=FK；н�Aͻ�vƼc�P<��<�/>�߿�p\�s
��7$�bMܾ:_!��h��/��=)y2�rV�����Z���:���1�ۼ%��=�%��\���i��C���?b��?*����w� o��A����$�N��>9����E<:8�����=ި�E���R) ���9�U��q�Uf���'?�����ǿ߰���:ܾ�  ?~A ?W�y?��Ҟ"���8�� >�B�<o5��˝뾤���	�ο������^?P��>��4��U��>��>Q�X>MHq>����螾%�<��?�-?��>'�r�X�ɿ|���=��<���?K�@��@?��)��M�.u=�o�>L�?T�E>�t7�x� 髾�o�>���?���?o�$=A%X��	�2d?f�;�\F�%QY���=A��=��0=�����F>~;�>A"�@H���轸+<>�ˇ>�6������k����<��U>��۽`S��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=ǚ�+Xѿ@� �J� ��A=����S��<�����ID}��v��?ھ�	Q��
>�u�=��i>1�>�L>`G�=7/a?P�q?2H>zq�9�
�����ƾ��C>/��˽s�����/� ����)�K����y���0,�}c��T��%/E���t=��a��Ɏ���"�\s���E�;?:>�f�vac�h~f������gz�R��=��W���ž|h6���w�?��?�F[?]P����;������db>�1�6?�$ƽCT��ޯ�*҇=.�̼?!<���>E�E=N����V�0jY��=?�,?�c��+�����/=\���D6��97?7:J?8�f>y{�>
�$?@���ɼ{�=�q>�8�>ߊ�>`�>��}���A����>=�S?#�������$�>ʻ��'zt���=ת�>\�-�ؤ��[�>SY >fO�R��=��=��=��[?���>\z�հ�}ʾ����m�
=���?+�)?��>�'w?��4?ը��u��9:��!�Sny=� N?��q?!a<���=��uu��AJ?�RM?j(<�V,���
���J����	�?5�V?�}�>'���R�撿�����?k�|?WQ������ /�b�D��D?P	?�+?6U�w=��O?{�k�#������o)�N�?��@.)@�t=H�V�[>%Y?�7?E�����	��cL=�Zľ4L��H?t/��~���U�̋轃�?��N?,Z?���{��vD>&�����?�4�?Q���sj<K��jo����Vm=xq>s�/=y��M���M�}�ܾ����\G��7-���0>�@8�:���>XP��1dҿ^ǿ\�{�@þ��я��C?�4�>��U�HK���}���{��}E�_A�$��"Q�>z�>M���/�n�{��m;�������>r����>1�S��%��˚����5<@�>���>�>�?���὾�ę?�Y��<ο�������\�X?�a�?8o�?x?5;<�v�d{{����+G?�s?�Z?Z�$�6]��r7�0�j?Pe��X`�L�4�>BE��CU>�"3?7C�>�-��E|=X>��>-O>�(/�ΊĿ�ж�N������?9��?�o�A��>�~�?v+?op�^4��D7��o�*���@��7A?32>�����!�3%=��ǒ��
?΃0?�}�H2�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?��>�Ċ?2��<��>��J> �ɾ�"����>�S_>퐽?�?@�@?��>�x>�lӽ���M8��SA�5�پ�Y��G�=�jO?ot?߄�>����R�<g���!��dy���)��u���DW���.�샹>0��>e�?>0�T�bD��V@?�#4�Pۿ�����C�=z�?��p=�-?���c$��U�\�{?]�>�,�'����F���,��?�G�?W��>�)Ӿ�%�=Fn�=	L�>u�{>#��<Cn���b��>s>�;A?�����g����"�h��>��?�a�?�ȭ?� m�z�?��	�v���P���}�K;��}��=�M;?�T��!4>:��>�k	>��q�HJ��|�o��>�>]f�?��?�~�>j`]?6�_��9�ӷ�=��b>	MZ?5�!?� �`��R�L>�?g�
��8��X����_?.�@"�@^\?�Τ��-�{���Ǡ�g!��_�=��=)�W>M�K�ss?;�L�>������=<��>��L>��Z>W)I>��>��=���� �'����h���M=���Z��[�E��.���r������J��b�"�)��`o��W�9���������b�=�S?'_T?%�o?.l?R���i>/�Ѿǌ,=@�4�;n�=�p>�*?5�C?�0?*>g2|�4v[�	F�����������>�1>	��>E`�>r��><�l��+_>t�f>C|>��
>5S~=�o=�wL=TPK>3@�>�_�>��>�>��#>�����kd�%O���b&�?|���J��ʚ��啾�M����=��4?��>�ސ���ѿb���4�H?j�w��
�/���">;.?��=?�,U=����]G��di>k�"����3zW=��}9S�B%7��R�=1?X��=v�}>�H��)��:��u%�<��?X���_>M�����9XI�����t(>���>���=d�2��n������*��FL=��M?j�?��.�46@�����n���>�,�>uv�=�J =u-<[�N��D�v�"�����p�<�M>�0
?�B=]BJ>s��>�����.��Z�>0>m63=IJ?|�?<��;2\��P��U�q����=s3�>��]><d�=tFp�x<�;%K�>.�2>t�z=$K��A�B���L��X�=�����)>���y��kx0=��=��V=]�GV�gc2��~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ$�>�K޽�訿�3���a`��t>@�f>k�O?�q�����𙕾�3?�)?��5�������п�����s�>�	�?�̨?����D䒿$�Q�]�>�Y�?��6?3=�>
+ﾩp�=>��Z?=�7?P�>Q�
�b����?��?ō?�&�>	&�?��R?�+?3x�p�2�⩤�?�c�*��=�>>SĹ>��>	�T�13'��x�����ZA^��A��5a>^(=�� ?�y����ž=`3i���Xl�=�}?w�>/�=��>�?H�>@9�>5�>��s�M���q U���K?���?����/n�f��<4K�=�^��-?^L4?��[���Ͼs�>��\?6��?A�Z?�_�>B��8��Dٿ�͛���ؔ<,�K>g�>�P�>,ډ��JK>��Ծ#�D��R�>���>f��h6ھ/������K�>ua!?�}�>�ڭ=�x ?$�#?�{k>��>�D� ����D�`п>:��>�? ~?�!?�~2������
���Z��|K>�8x?Xd?#K�>d��������»o�V������?a�g?i�L?+��?y\<?�~??'�m>����)پ����9�>��!?l��9�A�jN&��`z?�F?d��>������ս�Qּ?���u����?g\?�@&?�S(a���¾��<�#�xU���;xrE���>��>�X��Qմ=:>�Ű=B5m�nG6��7g<�Z�=vw�>e�=@7��=��j#5?c?��lȟ�Kl;�A�����	�>�2>;���W?d��U���u���ڙ�߽ɾ��h?4T�? ?�PI�o�b�^�3?}��?$1?Ss=x��$�Ӿ�����t>�L�5�#>���>�^��m���ש�����+���vf�;N����>}��>��?�>i�;>��>�c���2%���,����X��i��8�~K*�����<���+:��No���[y����>�y���J�>&� ?/�r>�H�>���>ô�;�DS>�mM>�k>�a�>Ko>�>���=ϖ�<�3�ePR?A���Η'�-�ذ�,�A?)d?"��>�*c�X���i�t?�X�?�i�?:�u>�zh��+�p_?@��>�{����
?��5='(�7�<�%���l�!���+�l��>.�ؽ=�9��L�hh�1@
?�U?����~;�ؽ�*z�<��<J3�?��:?#���=��T�\�_�0Fk��bo��³���v�E5�_p��'������[.k��� �]r=P�?�s�?q���Y�-'����]�@�=�kR>�|?�/*>��>j�/>�:��0�&�9�I�;�A���_
�>�)p?O?>xi;?EH?��G?k2Z?n=�o�>�ҽ1��>�Z"<��>���>��#?�b?p�@?2�(?�/?Y>鲍��P�nx�]?���>��?�<?�}�>O������;��>��%=�h(����<t2>�d�=`��xP��퐻=�tw>^?�q�g�8�C���T�j>Xt7?�z�>��>�⏾������<I�>f�
?S_�>`����|r��X��X�>���?�)���=_�)>h��=���Ѻ�N�=v+�����=� ���#;��3<(W�=Z5�=�gr��Y߹-�:�݉;R��<�y�>��?���>�=�>�[��X� �4��k4�=Y>'ES>��>jGپ}y��&����g��Dy>�s�?�v�? g=&��=ir�=�i��;=��M��,�Ld�<��?QB#?hMT?֍�?q�=?6h#?��>�%�K���\���&����?�,?��>�� �ʾ��.�3�h�?S?�:a�p���<)��¾F�Խ�>�[/�~+~����D�^M��A��!������?���?�A��6��i�ƾ��`����C?[�>�i�>3�>9�)���g��#�5;>o�>S	R?d9�>�P?!2{?!�[?ɐS>#�8��I��ɮ���'��">8@?;�?���?
�x?���>Ź>iw+�gྟ������r��(���-�V=xLX>�^�>*G�>Oi�>?��=�Y̽�	����>�L�=��b>%J�>�Y�>��>0*w>r��<�H?Μ�>*������T+���B����M��au?X*�??,?v=^���D�.����%�>��?���?��(?�.N����=�t缙ൾ�p���>�P�>vq�>&`�=�=a=�,>���>U{�>NX�7z��7��WQ��?vVF?��=HϿSW��h�\��ˌ��;�M4���93����Ð��@�ԺS��>�g�P���qC>��`��79���������厈�W��>IvO�S�=�=�=���<X&P�W9%;���=�q!=��;#��ti�<��=J$�=�᪽���
�=��>�����:ƾu~|?U�G?��.?\D?�yo>�s>�n��X��>�_����?��E>�&���񽾎�9���Ƴ���Aھ!kԾ"Ca��u��\�>Wl����>R|->���=c�<J��=iw�= 6=��:��=�Z�=��=�;�=�]�=w�>�x>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��7>�7>0�R�>1�)�\�n�b�>�Z���!?60;�?'̾��>e�=�߾��ƾy.=��6>�Oa=O���S\�V�=��z�
L<=��k=e��>:�C>��=�Z���Ƕ=��I=���= �O>������7��:-�e3=���=��b> %&>XZ�>��?�0.?f�\?��>��h�c Ծ�T���U�>1��=4F�>�i=^�=>�^�>��0?�A?K�C?W-�>��=!v�>n"�>Dt)���t�e꾜#���x���Z�?�?���>�/<K�����9�v��s�?�2?�.?�5�>�)���+��l��u���3E<�L�=^���j��T�^������T]�5x�>b�>��>ds>�t�>=fl>�
�=@5�>�ױ=e�ѽ�Jk�˧<��ڼO����>7.=�<<_b=ϼ�=�ۍ=A��<�?=lT�;�n>�ٽ=�\� �=I��>rp!>���>��'=������:>���� O��[�=|֡��=�Α`����C21��m@��7A> �S>+����Ő���>#.Y>�8L>��?@q?˗#>R����پ�(����`��{4�Bu�=@��=\aF�ٞ9�$_�D�O��ɾ��>�Mc>�>�#�>��T��M"��FY>����J�M��>dd����<�j߽p)��=Y��3����C�I�ܼD�??�M}��FS�:�?�I?��?��>
á��{�����=䔾!�K=y�־���]�=a�?Kx?���>d��l�<�G̾���$߷>�=I�s�O�/��0����̷�-��>������оU$3�Mg��������B�Nr���>N�O?e�?�8b�bW���UO����&��zp?+}g?��>WK?�@?"���w�q��@t�=�n?���?�<�?�>�D�=e*轢t�>6)?댙?�1�?�cy?J�<��u�>���I4>vݟ�8�4>�X>&~>wx5>�[?�T?���>�מ�)������򾣋l�}1M=Ou�=E�>���>�
z>���=�N=sI�=��f>�V�>;!�>�>f>��>$�>�@��`^�k�(?Et*>�>��*?Ԩ�>tB=�O�ꑉ=����##�nl�P�"��Y ���μk��<ā=B�����>l�ſ��?pI>�����?�M��(����T>8b>�|��C_�>��0>#4�>1g�>���>��>-Њ>�ď=�mɾ���>�(��� �k
B��[G�w�۾(��˞���l�}��"�1���I�AϾx��z�T��\����T�랓��;�?M�O��肿L�A���^?���>Tx]?֖�R���̑>�>���>�-�~v��~�������Nt�?�@�;c>��>8�W?:�?v�1�H3��uZ�,�u�Y(A��e��`�p፿�����
�V����_?��x?�xA?�P�<r:z>G��?��%��ӏ�g)�>�/�#';��C<=�+�>�)����`��ӾR�þ�7�IF>m�o?8%�?SY?�SV����j�=��S?�1�>�t?OE?2�>?�h=>!YO?�?�?�	'?�K?�aL?��R?���>�[�>'V�=+1��1ZὨ��,ﶽ����[ƽx�v>r�j>sO��9O��]:=����0�%=�G�<ﲰ=m{�<�]<�J�=�`�=�F	>��>R�]?Ű�>���>��7?A�i8����G�/?_�G=�n��?k������f����>"�j?X��?�Y?B�d>W�@�Q�C��j>��>��$>|�[>Ď�>uq�oB�H.�=�(>"�>��=�FP��<����	�+8�����<&@>P�>� }>n��B	+>u�����~�+Wc>D�M��񺾞JT��F��!1���u�^(�>fpK?\?�i�=�o�6ߠ���f��'?O�=?(�M?��~?�=ɡؾ79���J��M�>d~�<?��.��JL��|�8��޳;pr>T���M���<��>���NR뾢9_���U���C  �A
�(��=\�6��R����ƽJ�d>�B�>��"4��J��{���/E?/C'>>n��`*�v����>�|> ��=�=����()<��I��m�>�ݾ>Bj�<`�3�
��Y:�H��'a�> kD?��^?z�?�J��
ir�B�ke��g���s߼�?ݙ�>��?v�9>}��=X����/���c��E�a��>\'�>�|��:I�����:��B�&���>ݛ?��#>�N?LjQ?��?��^?�D(?�?(�>������I?'?5ۃ?d�=�pƽC!/���6���E�� �>��4?�7S�vݕ>B:?=�?�R ?#�I?��?ą�=�9ᾫ�6���>�J�>eNQ�К���<>��J?r��>��Y?���?3GU>J�(�b΢��DT�"#�=�(�=՚7?)�?wv?���>��>���}��=��>2�]?>-x?Oom?$��=U��>?�s>���>E�=���>G�?�$'?�^U?��|?��F?I��>?�<LS��,餽t� �!��}�
<��V<jt�<l g�����	ȼ�rW�c������׵� 閼hHݻ1��<D��;�X�>�(n>�F��P�R>R�ܾ����^[>I�7�(���Qi��QW�t��=��>=��>�Ȍ>&�B�=[��>�r�>����?wy?�i?r��<��X�Zb־ukU�
�>;<?OJ�=3d�[�����|�^�=?o?�+T?$�^�)��B�b?��]?!h��=���þ��b����r�O?>�
?6�G���>��~?P�q?6��>��e�:n����Cb��j��ж=?r�>-X�N�d��?�>i�7?�N�>��b>}%�=>u۾�w��q��j?|�?�?���?�**>��n�N4���VW��W:h?y)�>U���N� ?�$=�ݾ�i���������Cۤ�v����睾h ��eg�򧉾����e�=��?߄d? �j?~�a?�ݾ�$`��:S�H%z��oZ�Q���NY���>��:��X:��m����`���9��6=����P�a��?�jP?8��R��>��<�]�H]���9>�����Dѽ�F >�.2� ���<!����}0�\���+��>�>��>�qT?�n
��U7��]�4 ��.2���=UIj>E��>���>�Q�<�K��_��9t��:�Ǿ�kѽM,w>Qb?��Q?K}?��s<��s�l���G������s����>�O_>��5�Y)žpp(��%�$�^�Q O��ξ����޾�s�=�TH?�"k>x$>�݋?��>��=��x����=�nuL����>��u?�%�>�Ja>��A>�z�x�>�rl? {�>Mq�>ر��h� ��
{���˽~&�>�b�>��>,p>W�-��v[��B���0��:�8��z�=V�h?������`���>]�R?��Ѻ�N<���>����]!�U �4+��	>8\?k	�=�M?>�ľ<���z��ʉ��8'?aI?~䋾�j)��@�>��?�}�>h�>�.�?>T/���V�R�?'^?�$M?SXC?�>�bA=�����dɽ�(�`u#=u�>�8X>�m=N��=c!���g������V=���=Y$ܼ�9����(<TЏ���<��=|�.>f"ҿDjC�>������`k�:��+:�<ާ��@��S��������/��ٽ�a=_���%νUI��>p�����? g�?s�k��,��������S�7�p��>qkC�!���zξ��½Z�������w��N��-|�w���W�|0?�T���¿ ����ɾ�OT?Z�+?��?4{�,�Q�Ɉ5���> w.>p�u��H��袿�Oȿ=�����}? ��>��F��r�>�&>)�n>�Ύ>j�����5Ὡ��>ś!?�?a���h������NL=U��?&V @LEA?�(�"o辴Yt=���>�&	?N�E>A�4����S����~�>���?G��?-�F=��W�R�N
d?�<IsE�z��%��=�f�===�t�ǚH>N�>�h�]�C�6�ݽ^�1>Dن>y�(�H��u:^����<d�]>��ս�ߘ�5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=u6�􉤻{���&V�}��=[��>c�>,������O��I��U��=q �~ſm�'�,0�ac6=�܋9C��$�:������a�ch��f����V�6e>.>���>F�>�;8>�L >	>^?��p?Xr�>_�=�r�d��q���P!����$�>�ut�������1þ����in澛� ���!�������:�8��=?�N�ɏ�S!��e�LQ�O�1?��>pҾ��$P��;�����|���|u=~�I���о�l=�`�r�ח�?��O?��x�w�J�4����A ���B?<���f��S]ž���=b,+<�~�=�I�>�3�<�v	��<=��[��"?�M,?�:���Xj��"�>�������>c?�}?>�ٽ�{�>��?�W����4~>�&�>E5;>yd?�1>��þ��I��?{�7?��Ѿp]j���?Ư6�#"_�|4E��1 >=��o>��(>��Z>{u����a=�ϓ��Dd�:V?�c�>.�(�+��m�v�i�;�^��<Ւx?M=?u�>u�f?r�??\�;?J��N�����=a�Z?�g?�>Ƀ���׾V�����4?F�^?ZJ>>IT�=\�2�2y�a?�po?j�?ݗؼC�y�Vݔ��
��o6?��v?s^�xs�����P�V�f=�>�[�>���>��9��k�>�>?�#��G������zY4�%Þ?��@���?��;<  �T��=�;?m\�>�O��>ƾ�z������1�q=�"�>���~ev����R,�f�8?ݠ�?���>�������C>P���N�?g�??f���g�;����k����LVH<0j=��~�e޼]Q�]>�2Ҿ/
�G����n��Sk�>P�@r�rd�>��=�L|ݿ��ʿ0�}�MyϾk�u�(�?l(�>M"��-���Cf�t8z��e9�&*A�B���PM�>��>Ѭ���瑾��{�0p;�6�� ��>������>X�S�x������}55<��>���>`��>����齾�Ù?`O��;ο������r�X?�`�?�n�?�}?�:<N�v�V{��!��&G?�qs?x!Z?�X%��]��6��o?�����(]��<��:W����>��C?2#?,B6�<�����>�a�>�~7>JJ��u���Y��nC����?��?��߾4 ?�F�?{�D?��>��v������������<��q?VX�>����O�#N��s��!=$?��B?��	O&�T�_? �a�I�p���-���ƽ}ۡ>,�0��e\��M�����Xe����@y����?N^�?g�?��� #�U6%?#�>O����8ǾE�<���>�(�>�)N>;I_���u>����:��h	>���?�~�?Hj?��������U>��}? �>Y��?}��=��>E�=����/a)�w$>��=��>�J�?ʵM?�A�>�@�=�"7�׮.�zF�_�Q�z��,�C���>��a?�<L?�Nb>T淽.�!���̽g�0����yd?��C+�
$޽�7>��>>w�>�=E�H�Ҿ��&?�9%�zcԿ�����p?��X?���>�	?�~	�8�Ѿ��
�pkk?Ŀ�>����ʭ�����F�3��ɤ?�L�?x�?�<¾J��L8�=�{>}�=>i�ɽi���< }�:�W>J�@?�!�L����y�rOH>�o�?�t�?{��?Tug��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?mQo���i�B>��?"������L��f?�
@u@a�^?*zٿ3�����h�|��>�&��WoY>G�=��=�~U>��=H�Y�aL>9f�>^�>�d�>LO�>���=��ܼ�c�� ������c��=�4�L�5�.�&�`���Oھ�����2
��aY��X�<�ж�Ǯ�~R�}Ui����=��S?��Q?#&l?��?b���Uy#>~����"=r����=xɈ>G1?^RL?c�.?�3�=j���{ic�1�����������w�>�RK>u��>x�>R�>���$�<>�N>c,�>���=�%#=aK�<P"=�U>2:�>���>˴>��:>�
>�u��x�
Jh��uy�{�ӽ�t�?ٜ����I�n��B���絾e��=�.?�>?#��8NпR ���H?���)��p�*��%>r�0?��V?*}>h����Q��m>�v���h��5>���]�o��)��<P>�?��+>���>U)�t}3��GE��ݾzj�=!�?������O��8P�I�����>B��>6�X�֊1�����Ë��96��6�=�.$?�	�>� Y�n��s�@�g����`w>��Q>��ؼ�r?=\l>�y��On�����@G��7�=�6>�?r/>I>��>������2�43�>DO->Ǖ�=�� ?g�?�x��4���WW�>&L�=�9>f��>p��>�bK>3�e�-���?4��>Z =��)�����z眾AI>?�J<��˾Kc�<��>���>Gz>m2�=�1���j��&�~?z��*䈿��Ed��'nD?�+?]�=��F<��"�	 ��zF��D�?1�@�l�?_�	���V���?-A�?.��0��=�|�>�׫>�ξޒL�(�?��Ž�Ǣ���	��)#�	S�?��?��/�ʋ��l�;7>_%?~�ӾT��>�n��R���UO��6�>��>zkM?;�E�������G>?� '?Qz޾0�����ο)��%ȑ>���?kh�?�ō�=���$o����>V�? &�?��>Us�:��k]#>��0?�F?�.�>Z����rz�>Ղ�?`��?��c>�|?��b?Ɔ�>9T�=S����^D����Q>�z4>�&>���>��V�n������Rd�C�M��G�*@>���<��>n`ܽ���3W\>l�=7�ʾw�˽�H�>��f>���>M[d>�^�>Ƌ�>�C�>��>�J�w����@B�l�K?ׯ�?I��{,n�'��<k0�=b�^���?�J4?�aX�' оI��>\�\?���?��Z?f[�>���qA���翿�Y��$D�<�K>��>"0�>n:��elK>yվ�6D���>X�>�U���&ھ�U��zή��<�>�e!?�s�>���=��?��?�Vz>#6�>'@�f���A�v{�>n�>3�?}�q?H�?��˾��5�#��lע�_�U���8>ʉs?? R�>�掿w���=5�O�Vd� F|?�u?H>���?*��?`�>?[�6?q:[>ݢҽ�X־����fr>�!?����LA��-&�_��:?GS?���>�y���Aӽ1ϼk���'���.?�\?�f&?v:�u�`��\þ�:�<�p&���F�{6	<�XL���>��>ì����=�n>���=H�n��6��D{<]Q�=2��>�#�=86�2���>,?r�F��ǃ��)�=��r�0kD��>>@L>��ڛ^?� =���{�^���i��'KU���?ޙ�?�h�?yc���h�}=?�!�?n"?e��>(8��\޾���WEw�x8x�����>@��>�l����.���Ǔ��y?����Ž�Dӽ��>Ƀ�>NU?��>k�W>��>���ư!���(��vL���TLA��S$�o:��4��"'߽��ƼY������X�>��v��>��>41h>rFk>� �>����}>&!>цw>#ٚ>=J->K�.>�	�=�������R?����'�'J龱�����D?`�d?ш�>�|�Ŕ������ ?ْ?阛?V\s>��i�|D+���?r?�2}�s4?�==��ûծJ<G���������]a���>wc۽��8�hK���m�c<	?[�?�^��XTɾ��Խg�1��)����?�e^?��)�B�A����0R��W���C��h���J�ý�N0��i�"���f��[Y����t{=��?ԉ?\u(�����3�]�P�3k���t>�m/?�q>B+�>o�}>J�]�#�Ж,��P'�����_.�>)vR?o�Z>��0?��:?��?�sG?U�>���>����{�>K�>�V�>Ƨ�>+?s-?U�r?!�+?��%?=o>�d�p�վ�	?q?��><��>�T�>܉���O�_mq>ԥ=`�׾�ot���>�>}_�=���=ͯ==�7�=ʟ?�y��8�I`��X�i>�8?_X�>Ȝ�>D֐�1Z���y�<[L�>�p?^�>�����s�#����>� �?;����<�)>=��=\�������(�=�μ���=N�����9���%<W�=��=�����9�(!;�a�;"#�<1��>�?�k�>S�>є��� ����%��=VQZ>��R>Z>�ؾfu��C	����g�;\z>�T�?�}�?8�h=�p�=�(�= ����L���������mM�<.�?�*#?"+T?0{�?��=?�p#?�T>�-��$��_O����?�2,?��>�s�6sɾ�P���3�D�? ?03a�M����'�dQ¾J�Խ[>Y�/�Q�}��T��sC�����ճ��"��՝�?��?�N�/&6�Z2�8���^b�C?G�>��>P��>�e)��Mf�B��(9>���>�Q?c��>��O? �z?z�Z?KX>�h7�����ͳ���(���#>�@?���?�%�?A]v?Mu�>�>`�-�ӭᾊQ��?a�pb�����kq=��U>�H�>m�>�q�>_��=��Ͻ����[=��ח=q�d>ւ�>瑤>���>�>���<mkI?�-�>�G����
�rDo��y�����o?m_�?��?���=M�� jF��<�L=�>r��?\Þ?;>?�'�Ӟ�=$e��6��Sn��Ƨ�>�+�>�:t>8�=i�A=�?d>[��>͑>Z$����	���,��C�c+?83=?�Z�=_�ſ?�q���p��r��U<�Ӓ��d��F����Z��;�=����d���R��r�Z��d��������X>���N|��w�>��=ĝ�=#�=Bq�<H]Ƽֿ<�LI=0ƌ<=OXn��o<�V8�.�û�9���.�&&]<�[H=�-���Z˾c�}?/DI?S�+?s�C?&�y>��>��5����>�5���J?$PV>S�趼�uv;�����M��[�ؾ�O׾�c�̽���i>R�G��>�3>T��=��<M��=��q=j�=��`��=�$�=�$�=>5�=8[�=�N>�.>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>e�7>�z>�R�|1�TU\�l�b��VZ�	�!?�;�|(̾��>^Q�=��޾8sƾ�0=e�6>}2b=�o�3T\��i�=�t{�9I==��j=Ӊ>o8D>�ƺ=�尽�#�=�J=7�=.P>�f��s'8���*�)�4=c��=��a>B�%>�f�>(s!?�z?m^?jC�>�w��SS޾iQ���6�>�$S�\$j>�n�=r�����>~�1?�QE?�$?	�>B M=è�>t2�>�*�r؅�����av�{3�ZÐ?P��?���>]3>���ض��u
������@?P�?�,*?��>D��`���R��S�il&�������=4Խ\=W��>t���'/���>��N?oQ�>I�>"�,?�>-:�Rd�>� 
>ܨ>]su���I�/�,>s��=Ai}=�ۼ^�нr���϶=�3�=�Y���&��"�;6 �<��h�hLu�Q�=���>js#>���>�Շ=;���M5>U蘾�L���=C���t�@��c��#~�I/���5��M?>�X>1
��ң���� ?�kY>x�B>8��?�ds?��>U>��b־�6��1@d��QS�ν=jR
>4?�n�:�n2`��yN��`Ѿc��>�B�>�f�>\L�>��D�_�/�Rq>��6�=�>ܰ��s<�X�B�X�����YG��X�Q�%06=��H?�����А=�g�?�<E?�$�?���>$Ľ���[>E�b��.�j����0��� �;�!?�K+?5�>�.��yC�8<̾d.��3�>)I�J�O�	�����0�n��H�܇�>�����оm!3��f��>����B�Hr���>��O?I�?zb��X��UO�e��H@���e?zg?�#�>�E?�??�������6s���w�=��n?��?�8�?v>���=sU��*Y�>'	?豖?%��?^hs?y+?�hh�>lȢ;9@!>�옽	��=1c>V9�=��=A�?)�
?�
?�M��r�	�Y��ª�+^�0*�<�ȡ=W�>8�>�;s>l��=�c=���={�\>���>}��>�e>\1�>��>��b�c&�???�S^>��<��.?Wc�>�K]����P<B��<��N��a�+�U}
��=��ٻ
��=b��<��>XP�����?�=~�¾O?&�Ӿ�=X��]>|�M>ID�����>�K">�h�=�#�>�Y�>]�= E>R�4=@Q�����>(@��|:�Up.���n���E�,�&����;.s���(�y`>v5��(���M��"���|�IR��x�?>+���U���,�G&ҽ�H?��>O�F?�嫾:�O�EV�>��C?a>r�#�`k��|:������Xn?�8�?�\>+f�>]�R?�&.?�Z���M�a�R�ht�c:�sCh��gd��t����S9�rƈ9a>J?�uZ?�Y7??�����>�Fl??�6��1����>=�$�383���>:��>(�Ǿ�����������BsZ��?>��m?��??˝f���m�K5'>��:?�01?y�s?X>1?�~;?�s��N$?�7>��?>�
?��4?�K/?] ?=5>���=�?��4	=P����Ċ��Ͻ�ƽ�*��H5=Q>{=��&�ި�;�F#=T$�<	s����2�l;�_�����<gD=g�=���=���>��o?:/�>U��;�6X?�|��{P�;��a?'y?>�K���������Ȝ����>5z?��?*�?�l�>�H^��^+�J���f��=���>�'�=�g>j\��R���@϶=1�*=!>��=z�C�����'���]�)�;�o$>���>��{>Sۊ���(>�y����y���d>@S�Pʺ�МS��,H�ƪ1��Hu�{�>׎K?̦?�'�=���B�����e���(?��<?��L?��?z�=gm۾$�9�TVJ�'��o��>��<��gˢ�G���d:��|�9$�r>����p��Ia>q`2��2��P�#���J�I����U�־��>��C�r��s� >��>�۟>c�te:�����Y���d?�r�>�6���O�#����=g_�:�|`>��>��=�I�v��>�>���>G(#>=���T���j�o̾qQ�>��;?z�Z?u؇?�N;���q��zL��Ȑ�J����?��>Nž>З�=�$�<@M�����V���1���>���>�3��C�ݧ��J3۾�'���>��?d�T>�m?�XK?z6�>�W?��??� ?Me�>\�׮��&?y�?2-�=O�ܽ�T���5��nE��Y�>=6*?,�L�Z�>h�?��?B� ?��K?"?=v>+W��0;�v��> ��>�X�oY���iC>�F?��>��Y?�ł?5�V>��2������*��+��=��>4�0?w'??ޘ�>���>h���>�H>g�>�i?H��?d?��i=��?�'.>���>�w�=��t>�a�>я2?3�N?��?�/?��>�e�ϒ�7�*�9������<�Y=��<VfP=�/��Ss�������Ud=�!�=O��<�� �Z���ƽ�����X��{�>r�s>�񔾺*3>dƾ�A���@>�_���ߜ��.����8�� �=��~>�� ?�ɒ>.�%�qk�=L�>�:�>ԍ�S�'?�?�J?��;�b��TܾOJ��r�>&JB? �=��k�A���$�u�B&|=^n?d^?�DZ�i���N�b?��]?=h��=��þx�b����g�O?=�
?/�G���>��~?d�q?R��> �e�(:n�(��Db���j�Ѷ=Xr�>KX�R�d��?�>n�7?�N�>(�b>%�=iu۾�w��q��i?��?�?���?
+*>��n�X4࿎�Ծ�ؔ�O�j?��>ܸ��FT?b�`=0/ᾪ��Vd�:wξ���u����m��Ҟ����(����B�=,?�j?.1V?a�f?��߾�u`���\�v�u��\������.��)?���>�3�I��\k�̣��־����Bm�<0�[��vK���?~�'?%V_�Ċ�>�AX�����1ݾ�kI>�������� �=[!���P���'=�C����3��}���O?�-�>�I�>~A?%C��	7��2�G%4�Ax	��'>��>�q�>��>�G��](����j��񷗾X��]~o>� g?;�=?;�}?��O�q�C�¨����ul�i��V	�>��^=���;�̾��y�"��HV�{`��v�����\���^��=r$ ?���>?��>�˃?�'�>�Mؾ�۾7N���:F�e���{�>n�:?��?�I=>c�{�2 #�v��>��l?P��>���>/�����)� �~�$��wú>Kb�>=�?u)�>؉g�>�[�����p��&D>���=�,e?#0x�)�>���d>xgJ?�ػ+P�;��>=��#�(����� �Bn�=ER�>bn�<(kC>m��im�}�l��:��}m!?q[?�L|�x�&�ju�>�Z?Fm�>L��>E�?W�>�˭����<�� ?� Q?�J?�:?OU�> ȋ=:��"�z�7�Xh=�yB>��>34�=�0>� 5�t��N��	 �=�i5>�} =���c{^<�!=:p=��i�!>��ۿ��G��K��m���о~�
��B��)�߽����?���Ǿ\É�<�O�_"׽�Q�K��ݕ[��i��m���"��?q�?+u���� �$��JV��S�b�>`x�Qߖ�?ʫ�g����{�Y�ϾNL�����Q�M��&p���m�(�*?��?ο�����}˾�wN?��?�S�?<���MD���4��|�>@�>|
B>��������u�ƿOYu�7�|?���>t���e�=���>n�=7�>��>@��ƾG���6�?��4?q �>�z�� ���Ѹ��G�<H��?�/	@�mA?)����W=y�>7u	?��@>B�1�I�ʼ����>�+�?��?8�N=1�W���
��$e?�<�F�s"�W�=�j�=�=H��`J>�>���B�F�ܽ75>�Ѕ>f�"�:�T^���<�e]>�qֽ�O��5Մ?,{\��f���/��T��U>��T?�*�>T:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=v6�����{���&V�|��=[��>c�>,������O��I��T��=M����Ŀ�$�l�,�z��=� :�-C�]�ݽ��ǽ�Խұ��0rN�p P�:��=Y>��>l(v>Β>��>��\?��v?g��>�g0>t��@�����ݏ��-,���/2���L��H���+ξH8ɾ 5������$��뾛<�Ċ�=��U��R��L�bc���H�h&&?D�->�ʿ���T������؝������Yl��,�Ծݎ6���q�R0�?��??8A��!ZS�N�6D��̺��k]?A�形$�%絾�S>߶�;��<�*�>y�?=l�ѾQ�1��6M�b'?�2?���������	�>(�?��5f��L?��?�d�=���>V��>ӑb��y�鴢>Q�_>���>�s�>�W=�ֿ�୊��>?G`?�_��6(����>���Hɛ�n"��b>�E��ޚ�=}�_>Q�m=1�d��&��a�������Q]?R��>��"�D��pkf��
Ƚ���S�?0�'?�>V�j? TK?,�q���7�Y�eO>�K?��\?�$�=4���{�ƾe6]�}�P?9A?��>I���^s����D��j(��� ?f3~?"&�> ��=��Z�۟����+?:?��v?Rr^�;s�����n�V��<�>�Z�>r��>�9��k�>�>?�#��G��񺿿aY4�Þ?p�@L��?��;<����=�;?�[�>��O�U>ƾ~��B���d�q=�"�>����%ev����P,�`�8?Ӡ�?m��>�������4�>���ݧ�?~4�?�k���Eʼ����n�A���@=m��=�����`���==�,ʾ-�
��ҥ�����s>�0@v\��>`8)�1\ۿ��ſL-���5޾*��M{?1��>��ڽ�B����t��*���<<���D��h�9��>!�>�#���}��M6z�r�:���ܼQt�>�z�>q�X�!��bϛ���u<1�>9^�>��>���S���zę?V���bο����/���qX?ٞ?��?��?5�;<��x���s����AE?	p?�*W?�ＢdY��{�c~k?����u_�1�1������	�>��b?���>#�N��Z��M�>���>���>{���fƿ���E�վ[��?�3�?�O;�t*?�B�?D�W?�@8�-㾿T7پC`��<"=�Zo?%�8>s('�8�.�E�u�m�`=[?�?TY�O�0�[�_?'�a�N�p���-�{�ƽ�ۡ>	�0��e\��M�����Xe����@y����?M^�?h�?ٵ�� #�d6%?�>^����8Ǿ��<���>�(�> *N>TH_���u>����:��h	>���?�~�?Pj?���� ����U>�}?}�>;�?���=�|�>���=�<��5�7�}�#>r�=>�2�?z�M?ß�>D��=��8��/��bF��)R������C���>��a?]L?� b>�฽eg0�%!�u�ν�l1���缚�@���-��὇>5>�T>>�]>��D�8 Ӿ�~?F��DLؿ;���R@0�� 8?�@�>aG?���W��qK1���`?��>�<����h��r��d��?���?��?�վ����j>���>d�~>�B½7㧽Z���9>4EC?o&��Z��;�p��Ԃ>���?�@@I��?�Vi�<	?�%L��W^~�Q���	7�՗�=A�7?G�S�z>i��>ڪ=Ckv�����Ҿs�w��>�?�?�v�?B��>��l?~o���B��1=�O�>�k?�f?Q`i����1�B>6�?�������I��f?��
@�t@O�^?�ꢿ�t��7��5����r�����=�}j>�[�>3���,�:�4s'=��V�^q,�Ǧ&>+�e>׃>��>�i�>�Z=�K�=�o�����ea���恿6E��g�G��#-�����MV����hꦾH���]w�V�݅�̑G�tDֽ,����E�=�U?��Q?�qo?� ?�jv�� >t���;�=�$���=gP�>�A2?`RL?��*?EF�=����p�d��E��[\��>����>&�J>�H�>�)�>��>�r'�_(I>� >>�V�>��>'=����C='IP>ϫ>3U�>S=�>�<>i$> �����1h���v�n�ѽT��?CI��gWJ�Ě��R����ش��s�=��-?,� >����gOпU䭿2�H?zo��0��}a.���>�d1?RW?��">�x��U�a��>����i����=�v�n���(���Q>a?ͮf>ju>A�3��c8���P��~��@f|>m/6?�綾�A9���u���H��\ݾ2OM>ƾ>pkC��j����7��hi�N�{=�u:?"�?+O��/ⰾ��u�AL��|GR>G\>�Y=�c�=�cM>_Mc���ƽhH��D.=Ƨ�=r�^>�=?�>*��=���>�u���X�̱>� D>�79>�;?k�?��ּ���F����(P�ϳi>5��>vV�>$�)>�06��U=g��>[�?>��=��l���`�h1>O=��S�D�*�!�EoM=��W���>/V�=뛶���c�c<�\}?<N��B�������F[d?B�?j��=MM	���:�9��Hv�(,�?��@���?�v$�<�S�(?�s�?��_��b�=Wd�>�>
��K��?��
���8���L�<3�?י?>n���ˇ���e��_K>s�0?�̾���>�K��Ω�]C��e�X�ޑU>�n�>k"X?پﾊP@�!|���?~U?���������ʿ��y��)�>���?� �?�p���sn��9���>��?�+�?��a>����Ч����>ǕJ?�?���>�^���7��8��>���?4��?��N>�?�\?��?J q=#|S��j��1Y?��1�<PF=vD?�XA>J)�UdN��Gc�:����c���h��>А=L��>�F�u���Y��=�㗼Õ�ӑC�k:\>��=:�>5%>���>���>��>Ɉ>�1����޽����K?P��?����1n�ʧ�<��=Ʀ^�s(?I4?�E[���Ͼب>e�\?1��?�[?�f�>?��U;��.濿�~���S�<��K>�+�>�@�>����NK>��ԾsED�k�>�̗>�T���3ھ�,��=k��DJ�>0f!?4��>�ˮ=B�?�/!?-s>�ּ>��@��c��VE�ap�>�L�>P;?I�|?n?��¾t4��둿�z���X�.�=>��v?0,?�,�>eэ�U����~<��d��YԽ!$�?��l?����W�?H�?��2?:	>?��>\d�!Ͼ���?zv>��!?>D�+�A��?&����v\?�D?}�>Tȑ��sսWռ��ad��7�?K\?'/&?�{�r�`�4�¾I��<5�&���K��}�;;�M�k>2�>`���s��=�
>�o�=)Cl���5��a<T>�=)��>��=J�7�����wE.?~�; ���\a�=5f�d�E��b>��>����,�[?\�6���n�Id���ٛ�;����?+��?�z�?WP���"i�ξ=?��?qS?�C?����3ܾ�ؾX�����m���Z�=z�>5@Ƽp�о�X��6V�� �~�綷�i������> �>%P(?���>Q��=�I>p4�����Վ�E=���cd�.�)���J��.�����~�����F;<��ژ�C�>��@���>�?��1>���>�/�>��`����=�`>q��>y��>��=��w>a�>/�=v7��R�R?HMƾv�)���'��"�H?��f?���>���`���_��'#?���?�j�?�k>�m�Q�*�V	?,m?��y��8?Fa=�8�;����Y����� ��
�1��w�>����i9�+zJ�~q�T�?v,?{����þ�����k�7t��jf�?�OG?�#.��V��>;�%KZ�}�r�y��~n*��5��R����k����R����z���%���>I?��?���C4پc25���]�hT;� ח>'��>�~">L�>�L>�V�o#�4LM��<�h�V��K�>cdn?Wj5>0?BW0?(?CpL?�\�>�R�>�p�Ĝ�>Ƶ����t>�E.?�l?�_�>h�b?Q\F?tB?m*>�Mg����Ռ��j!?�W?���>�>+��>�ճ�W�k���XX==s�`�>�
��\�<�>>�չ��&	>m�5;�~$>�I?�u���7������h>Z"7?��>�>1+��ϙ��m��<&�>�
?=U�>$ ��7r��|�2�>y��?���	� =;�)>;�=p�k�#0��xS�=ۗüK`�=}���6���&<X�=Zd�=ho@��`,����:��c;�[�<Hz�>	q?0��>q��>�j��� ���1Ա=�g[>�XL>��>��۾������Ag�]^y>�~�?�W�?�.g=��=���=�ԡ�(����9	�@���=t?2o#?0#U?�ڑ?�c=?��#?�x>U"����c惿���.�?9#,?!��>����ɾ�@���q3��?R?�a������(��_þ�Nӽ%�>E�/��}�Կ���:C�ͺ���u��� ��?&��?�dD�G�6���qט�n����C?7��>�|�>�3�>�'*�6g��(��V9>���>�Q?��>��O?5{?��[?HUT>��8�)��������5��!>i)@?���?mԎ?I�x?T�>�~>� *��ྱ���� ��6傾k�V=�Z>��>��>���>�9�=�5Ƚ����?�+K�=�Sb>���>K��>���>��w> $�<�cY?W�?�ц��6�op���Y�����/t?���?�FL?�>�>���]�g о�]>���?ޓ�?��L?��ӽb">e-� �ž�+���>y�e>UY>��>vY>+^�>���>z�>�W��_Vp��ξV���~.?y�>2��<�]���os���M�r���>��k��x�C�����H\`�T��=�j���/�0ɟ��]L�Zˤ����<���9ꚾ�fi�o��>lYn=>��=ݭ�=��C=��ż{(<�&=��һ�� =Դ&�/��<O()�X�U<�!\�3��ʭ<R�=x��:˾��}?,$I?zh+?#�C?0y>9#>Wd/�cږ>����z+?V>�-R��B��Y�:�!{������@Tؾg׾% d�۬��zn>ҺL�'�>ߢ3>Gq�=[��<z�=Gs=l�=���=4=T�=I�=X��=��=��>Y >�6w?W�������4Q��Z罥�:?�8�>i{�=��ƾr@?��>>�2������xb��-?���?�T�??�??ti��d�>M���㎽�q�=I����=2>u��=w�2�T��>��J>���K��E����4�?��@��??�ዿТϿ5a/>��:>�k
>�kQ��s1��x[�ɮb��ZZ��2"?j�8��ʾ�>��=�޾�Ǿ{-,=�j8>�0m=xZ��[��&�=?ւ�R39=\�a=�>LC>���=�&��z�=J�O=���=�mR>w_�0E>�RM'�2�G=��=�-]>��">[��>,(?��%???�S�>I"M�7�龒<���y�>9����3�>�5�!)
>"�g>D�?�-?f?Ҏ�>)��=P��>_=�>Ew6������ �L���*>_��?���?i�?��9�A��
���L$��v��X�>�M?[.�>���>��<�;���#��V��M"�=I��=����;���v'_�<>.������2>�J>��>�>���>%�2>QNx=^	�>f�>g�=>�<lEn=�*��4���;$>���=RĽ�۽�W��=D+�<h�<S&������ƞټ4?>x�뼁#>c��>�k�=��>ٟ>��ƾY��=1�.�Bx.�u�=���9[5�~l\���|�
��1	��XI>D�m>���#���L?��b>m�F>N{�?��i?��*>�)�,���Q��d�G���X>�p<>E��N6��bu��5��Z޾
�>;Rc>S��>d��>�\���B�u>t⾋5����>�	�����H��bu�)�����i�U�=�8=��R?8Pk��2�Y�?6�O?8��?U�>��ֽ����Ʈ>F���ѽ����|�����*���A?��4?��>���G,���ʾ�2���Q�>:F���N�R���0��h�����v�>�0����Ҿ��2�;��e�����A��Tt�:̻>��N?i��?�f^�v<���O���O����?mug?���>g?L�?=���#��Z~��*�=�m?L��?N�?Y1>�8�=���[U�>v?�[�?鸐?0�q?��:�6��>0�;��>ط��4�=Fb>��=aG�=��?�~?�r?%��pT
�2���ֲ�3�Z��=P|�=W��>6�>lg>��=[ǔ=%A�=A*[>���>���>]�X>���>���>Ov~�+��^�4?ͯM>p��=��?>�>MK�:��彋��=WR�[��g�m��wMP�1K�<������i=Ԇ=&�>B���i��?�/�=�W����?�׾p�;��"I>ז!>xaݽ5��>�E>l!�>dܿ>�m�>j{�=�6C>�s�=׍����>n[�+�-�6�)��X4�p����t>���z�B8h�ָL�YHS>G��L��p�m�ji�*�o��RA�F�?�I_�R󅿱iF�C�����A?*��>�?'���{�r�p>i�(?*��>�0����~���dpa�#Xw?(��?j,c>o��>��W?��?�.��^3���Z��u�/h@�sBf�Cw_�$��쀁���
��]ĽQ_?�Aw?�0A?���<|{>�e�?�%�h)��5U�>B.�;:�
QG=�g�>����DIa�c�Ҿ_��;U��-H>��n?5:�?g!?�$U��q�C�Ƽ��??A4?�~?6N?@lD?���Q�?��a>���>��?e�	?��?�D?�>��>HF��W?�_ZǼ�U���ѽ�
��6i;��=��>_��U�ѽǎ�=Pǔ�hە��K7=���=fh=��a����=Z��=��&��r�>�>_?���>`�V>6?���8�����]8?�=J�e��/������%޾�>&�f?G��?�}^?z:U>�:?���B���>z�q>_�>>�`>E�>�#��w�+����=�t >	[4>���=�f?�K�q����!���5ex;+r>���>z�|>�{����'>������z�[�c>�P�/��/�S�@�G���1���v�3��>��K?Y�?f��=����H��fTf�.9)?V<?�!M?C�?!Ӕ=�N۾��9���J�����u�>�~�<���.d���顿o�:��4+��:t>$����,ܾ�ݧ>��;�p&Ǿ\�
�1m���1�/�꾇����2�>V�;���A�ȳj<|�?F8?���d'�a,��v�¿�G?ObS>~Ͼ�7=	����;�ڰ>��v>b��xNŽɎ@�����N�M�Y��>��>�x��;;%��a��#w��և><�D?_? ��?�䃾�r�@�D��\���О�K%���?�)�>5�?��)>齚=
�������dc���B��7�>��>��X�F�|���N���&�Fa�>
�?��$>u�?{�P?�R?@�a?�'?P�?� �>�ܽ�w���2&?}�?���=�ֽRNS���8�k�E�jA�>:i)?s@�ꔗ>�?�?��%?^Q?�s?_>��� W?�Ha�>��>R�W�JO����Z>�/J?���>�Z?RI�?q�=>��5���������,�=�>h�2?��#??��>�O�>b\��x	V>- �>F�b?��k?um?C�;>iR?�d�=��>hJ>+9Z>.�q>! ?\?_]}?�5?9�>Jq=�����[�h�<����@=h�=���=�xj�[�J�~����<�/��ƿ����<:����\��_�ǽ�/�<9V�>|=n>�˒��4>�až#}���gC>}Ǯ�S���~��ے9�]a�=���>#�?ɭ�>Q�&��^�=�Ի>#�>HV�0k'?�`?n?6��;�;b�̏۾>M�i��>w�A?��=Hm�~ᔿ�0t��Cb=N�l?-)^?��S���K�b?��]?'h��=��þu�b����`�O?+�
?5�G���>��~?m�q?I��> �e�-:n�)���Cb���j�Ѷ=Kr�>=X�N�d��?�>n�7?�N�>'�b>%%�=iu۾�w��q��`?��?�?���?+*>x�n�Y4�J�Ӿ$쒿��f?��
?�G����?d�d=�S۾@�Ծ�1���Užp���:��ef����]u����kL��7q�=�?��h?�\?y�s?��վ��i��CU�P4r���J���徐��QN�cN`�p5�M/t�1*���ľ��b�i
ʺ��q��9D���?�c+?qk8�N�>���,��ݾ�H;>6�������W�='�l�z� =�"�<��x��,��ꧾ�?�:�>�ܿ>��A?R�Q�4<>��h1���6�.����'7>��>v�>���>R�.<��6�H��sǿ�G�t�5���tl�>��i?�M`?Ӟt?FY���;��rx��3����������?���>�$Žz����R�u���L�#�Y�R�������D��n���/?�R�>��>8�?�+�>�v:�"e���j���<�UG�N
x>J�d?�K>ѐ�<�)L=�־]�>��j?# �>��>OU��!���w�k�н�m�>[{�>��>s�n>oO(�Щ]�d���a�����8���=mpi?k����f���>ZR?�@{;�5<v��>{�����"�t�ﾩ/�7�	>۰?�4�=��D>c¾����q{��߇��+?X?���5-��f�>�;$?���>V�>�?p�>�Ḿ�5:���?+�[?J?p�C?д�>I��=�����н���3��<b'u>ιs>��:=�>�=i���^�&��Ut=a��=M`��穽Jk�Kdu��0	<���<�=/>��ڿ�qR��z̾U��Tc��/�哾����ir�}�ݽ�T��3�y�秒�L9ֽL
=8���1Gg�ܠ��(��^��?��?]�
��|پ h���c���Z,��a�>�翽��.��㸾�I ����z}��ߞ���
�q[J�Ǣu�]��4:?��ؾ�Ͽ�������-3�?�k,?���?�]�� #h��e8��.�>�k.>ͮ�>�����������[ž�;_?xd�>ڰ��Э<-��>d�_>��k>ɗ�>y0��#'澭,D��i�>b�C?�>	��EĽ�B,���%q�;�?��@|SA?�)�-S��Z=Gy�>�\	?�A>CP1��������[�>��?h�?��L=h�W�M|���d?�]�;�=F�5���R�=�r�=�= ���J>Њ�>a��l
A��ܽ��5>��>y)�
��(\�<:�<�i]>�Wӽ����5Մ?,{\��f���/��T��U>��T?�*�>U:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?8ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=k6����{���&V�~��=[��>b�>,������O��I��U��=���eƿ������T�=B�=>u1��/	�lH��;V��Ч���\��^�����=�+>�zj>:b�>5>>��3>��Y?x�j?��x>P�=$����h����@�%<H�b��t �:�w�����:y��lپA-ξ�D���AA��6Ѿ[�F� ��=|S�������+6]�Q.W�PN?��P>y=����W�QN7� [�C}���B=�gQ�Ν̾�R>��g���՞?JNX?�#����N�6�꾌׎��+o�4k3?��1����􈧾�%�<�SD�-0>��>d�>⳾$�=�˧e�y�?F�;?сʾ�"���
�>Fܽ�=ȼ�@?�?,�����>@��>�yk��~E����>�~]>���>r7?�V�=����Tཛ@2?�?�V���ߨ�.̴>D���k���j��'v�<��yUI��lL>w|�=�ᵾm��` (� ���l�T?���>?�-���0%>�ȩ���V�<��?DD?_�>��n?Y#6?��;ī�oCG��㾃Y�=��Z?ehh?���=��g�9?Ҿ�Ҏ��88?�V?�UB> )F�}��j!@��e�[�
?�l?wh	?SS�;}y��7��e����1?��v?�g^�Eo�����?�V�m1�>SK�>��>d�9��u�>u�>?�#�I������S4�|��?Ԕ@3��?
<<t�Ř�=�1?Q�>�mO�?-ƾݲ������)tq=A.�>����
nv�i��u.,���8?%��?��>)z��c�����=�k��� �?g�?����?�;��D]k��o�u��<
m�=	�J��>�a��ݽ9��N;�7��*��殼���>�'@ۧݽ�D�>��7�3�˭̿Q"����;'�o��C?դ>O*��᧾P�l���t�$*B��RD�^���B)�>��5>Y����X��f4:�c{Q����>���zcT>�3���(Ǿ�ǀ�q��=��>���>��5>�����ؾ�C�?���_�ǿС�����1\q?�?�?��?~�?E�h��1�f��ǽ<��C?L�G?M�U?^�e=�8���7�ck?����`��H�FE���>9�o?��?y�:��宾�I�==�-?"�:>Б��ʿ�轿��� ��?Q�?zþ��%?�
�?��W?���BJ��T��� �IM�s��?$�>�b�����P��%���I�>v�?�jq��O���^?�`��q��d-�M�ǽ��>��1�@s_�au��'k�W�e������w�b��? Z�?uʲ?FG��{#�v$?�^�>]u��L�Ǿ��<���>x�>
kN> y[�ޡv>c9�/<���>�p�?B�?q�?����1I����>��}?s �>��?��=m?�>��=�԰��/��Z#>�F�=[+?�g�?�M?k$�>��=A�8��/��HF��0R���b�C����>��a?�uL?�a>h���0�z� ��_ͽ�_1�
��r�?��T,�mF߽kD5>U>>�>��D��Ӿv ?���0�ؿ�v��|(���4?k�>$?��L�v��w&�l�_?7��>����(��4:��2����?�?�?"�?�@׾��¼.L>�E�>���>gnӽ�\��}��q(8>ĤB?���*���o��͆>J��?�@��?y�h�U	?��I���J~�P��`7����=8�7?����{>���>=�=>rv�����ߴs����>�C�?
u�?��>֤l?`uo�Z�B�KL2=�e�> �k?�]?r�z�J���B>,�?�������r6�~f?�
@�r@��^?}颿�Eܿ�	��9����	��V�>i��>n�|>�@�������=��ҽ��J;��L>��>d^�>-�>i�>ȯA=q�=v����"��▿���7V/��}����&������' ��@����D:��>����5��*�]�V�B���Ƽe4�=ϢU?��Q?(�o?c� ?��x��|>����=�#���=HE�>�U2?��L?��*?d�=�I����d�ni���0���Ӈ�ť�>��I>hh�>��>�4�>,
.9�=I>;2?>᐀>XX>�'=�>�w^=ƕO>�W�>���>jV�>�_>��S>�ѻ��/���~�_�ѽ����?V�@���[�x��U���!����>3�,?d�-=�g����˿4w���<c?k������g�羄Q�=L{�?��c?-��>
����43�`��>+>c/��>�,����+ǯ�Ա�>��I?��^>�v>6�3�ܕ8��M��y���n>�c2?븳��15�.�t��#I���پ	�W>���>�# �*��IT�������?d�р=t9?B?�����a���Co�R`���vJ>B#c>z!<=�e�=�b?>�eC�{�����B���3=���=U�Z>�	?��>>�y�=��>�\��hV�Li�>%�v>�_>��<?'?s4��ҽ�چ�@�-���m>���>䇍>W}>=%2�É=��>��|>�1���J~�Qe�OO<�g�V>q�(��.F���Ͻ��<<�5��>#�=Q�`�>%&�.�<�~?����䈿�뾩p���oD?�,?��=/^F<Ć"�G ���A����?��@)k�?I�	���V�?�?BA�?d�����=a�>�׫>�ξ>�L�%�?��Ž$Ȣ�۔	��)#��R�?�
�?�0��ɋ�}l��7>Qa%?e�ӾI��>�C�jt��t.���u��}-=S{�>}}H?�����4V��>�k
?�K?8���x����ȿxMv�`��>y��?���?G=n�����z@���>���?i�Y?��i>�۾�nZ��b�>��@?��Q?Ӽ�>���-l'���?U��?��?��z>��?+�v?�a�>qǽ�� ��Ӿ��ca��)@>=>�?��>�����T������V�Z�9�S�$���>~�=�k�>|3=����h>�q"<wc̾�c��\�>�(k>���>)2�>�>�k?�f�>W��>L�7<�Ʋ���i�q�K?���?'���2n��P�<E��=7�^��&?�I4?�k[�q�Ͼ�ը>ܺ\?h?�[?"d�>-��J>��G迿.~���<��K>.4�>�H�>%���FK>��Ծ�4D�dp�>З>�����?ھ�,��_M��eB�>�e!?���>_Ү=��?�b?�P�>y��>G�=�������:�<��>t�>��>)�h?�l?a����[�{.��Ŋ��GPS�q�u>��g?TX?6�>�Ə����Z�ּڠx��ⷾ�;{?�5�?��L=�?0\t?c�.??�x�>:�=�⊾��5�
�>k�!?���I�A��Q&��]��V?�?�R�>�����Nս�׼����;��'?S*\?�Z&?B}�[Ca�օþ�9�<�%!���N��o<`F���>r�>c���\�=+�>�,�=�Zm�%7�;,o<gn�=Б�>��=�`7�n���F<,?V�7�r-��xЗ=�r��zD��">�BN>�L���^?E#<���{�K�U����T�I�?F��?]m�?|��E�h�W�<?��?!?�l�>"~��_D޾��߾��w��uz��j���> �>^C}�?��p������P���Ľ�{�I��>�<�>�)?C�?��D>t��>�#��e.(�m�ݾߖྙ4W���!��*7��]!���'��9����;w浾�I~����>���C��>��?�~z>�-s>���>���<:Y>o,7>i�>P�>��Z>�?>�>g�=��d�Q?4�¾�&�- 羽f��{3B?��d?�>g���x����t�?ϛ�?kś?ZTp>J�h��+�{�?�:�>b���q	?��J=vK��ʥ<�ܶ��#�GƊ�����f�>C˽{t:�#�M��`� Z
?~X?�/���Ⱦ~7��b��p��Ԑ�?�Jo?]4+�S�_�n+�Z�E�r|�{�����m����-���\�C���D���m�9���7�=�?�T�?�&ɾU�cε��~E�b�B�ܔ�>c 
?9>L��>.2�>�!G�0�[�S[.�Û �ZX����>�q?H�T>.�A?��:?�!?!�N?�ia>�=�>�2����>@��ӟ>վ?#T$?_��>��4?ם5?�;?�M�>��z���������I?!�?	?��>�3�>�;W��ʦ������s��\���f��H�=��m=��?<�H�=>�X?e���8����y�j>v�7?É�>���>6��4@��W)�<F�>�
?�D�>w �	�r��b�`T�>���?y#��w=��)>���=k+���`ֺ�p�=�;¼�ܐ=���*;��v<+]�=���=��r�������:^��;�n�<�Q ?�>?F�>/��>�+���= �����=O"b>��T>�(>�qվ��W�����f�):x>�ŏ?Q�?��y=���=��=q裾���1:
�������<��?&%?��R?.h�?��<?j�"?�u	>���8���'�����_q?e.,?�x�>��0�ɾM���r3���?�/?l�a�iL�=)��n¾��ҽ��>��/��3~�_����C�R熺�������C��?<ٝ?��?�>y6����е��O%����C?�>�ɤ>��>GP*���f�Eu�i29>O��>��Q?&2�>
�S?��?;uZ?hm?> �3�6W��%����ݠ<c�5>E�K?���?9��?'k?ȭ�>��*>cM/�������5�8)ܽ�s���p=}vO>8M�>]�>{j�>��A=o5佗Z���)/��Y=r%]>� �>\_�>�Ƭ>D��>��<:mV?�?�@ʾ�� ��6����b�k��_?���?�x?�d>�&@���W�L��xj�>�̒?�?�}?j����<0
=M���ց�g�)?d8s>��$>�E�=����>�>."/>X�/�=���@{¾A�[>���>d�?&T�=e�ƿts�Cj������<���6�`�76���*[����=�ꚾ�&��\��0,X�ঝ�v���U岾�&��V��G��>lr�=��=��=}J�<C<��ن�<w�P= ��<�%={e�V�<�..�KEֻ	���O�˅<�<=�����ʾa}?�UI?<�+?��C?M�w>�k>��D��5�>����V?�ZU>7�k�-N���8�B���ǿ��f�׾*@վ��b�܈��߷>�W�q�>��5>���=��<0�="�=fg�=��ֻ�=u<�=�Ի=6��=�)�=5R>!�>�6w?,�������4Q�5X�m�:?�8�>�}�=�ƾ�@?)�>>�2������Zb��-?���?�T�?g�?�si�qd�>%��}䎽xr�=,���!=2>O��=A�2�	��>"�J>����J�����O4�?��@��??�ዿǢϿ�a/>�3>Ҡ>
�R���1�"W�Ƹc��`���?��9���ʾP�>��=�ݾ��¾�@<=�;>�h=�����]�Bb�=�v�Y�@=�x=�	�>rB>"�=����Wu�=n�Y=���=�3N>x3���%����&>=���=�?_>|j#>�h�>O�?}/?�@?�X�>�V���[�ž�̈>��9>O��> P�<�<7��GF>g6"?�/,?�8?6ݸ>��#>%��>\0�>��0��~��8��׉�+�D�i��?�[�?y��>����ơ������7E��e?�T?S?/^�>ˢ�hT���˾8�ܾ�<	=H��<��(>+��g�/���~��Q�+i�>�/�>�G�>봫>¬>מ=-��ϵ�>�x>���=Y��=^�2=�Y���W����>P�Z=���镽X(�gV�M ��k8���|k=~�)�yQ�=������=�(�>�`>�w�>Ho�=1����.>W��Y�L�v	�=�%��X"B��d�5<~�8�.���5���B>.�X>{m�� ��U�?i�Z>��>>�>�?�Qu?* >|��z!־V:��if�cuS��V�=u�>��<���;�:O`�'�M���Ҿ�
�>�Z�=eq�>G�>�`Z��K����>ҺȾw܀��K�>��˾m/^=&Lu>�iu�f��~S���ff��}��b�e?'>c�FN6�J3�?�2-?
�}?�'�>-8ý��оؚ,=���A��ɾ����);N>�5?1@�>i>H����?�s��'��,u�>өQ�%oL�'璿��-��M <;
��ė�>����#�ƾ��2������q���=�q�m���>O?
ҭ?�d�7���J�y��s�����>�>n?V��>!
?k�?#뀽��޾�m�;��=�h?���?���?�C>���=j맽���>z(	?�p�?s�?Jr?�D���>ǒK;��)>R���h�=PO�=5�=w?�=j
?"�	?�	?B���R	��ﾦ>��Y���=$��=x��>&�>cx>��=��K=��=��X>4�>ӏ>g�d>�>�ֈ>�j���^���&?���=��>r<1?j��>�T= 3��	�<ͷO�v�;��K$������Q�O�<���p�S=�&��Dt�>�@ƿ��?��U>�3�Y�?N��Gr2�2UR>�R>6�ν���>D�@>�؁>�ٯ>��>a�>pX�>�>��Ͼ�>����"�&CD�@�N���о
�>�t��Ά-��-	� �]�?�P��D�;�h��΁�B*>�w��<�~�?	�
�~�j��3,��H��G?l��>o06?���r��y>z�>���>�����疿ό��^ݾ4��?+a�?�Gc>U!�>�W?I�?�r1�t3��lZ� �u��A�]�d�F�`�{ߍ�v�����
�L/�_?��x?�uA?�+�<jIz>]��?�%����>j/�&;�A�<=�K�>��k#a���Ӿ��þ�,�/4F>�o?�%�?Ga?UV���Ƚ�>(x??h?��r?�E!?��7?P±���$?�]�=O[?�?��?��??;?��>2r>���=?K@��ѽ�������%�-Yν��h=#��=���;�mU=��=r�=@�0�ȑ����>���g�o/�Cl=�h����=ϱ>/2\?�m�>,�Q>��C?�`�~5����S8?��=�P��������c⾥V#>�o?�]�?)�e?k�m>�FP�p�.�x�>�px>��@>�P>ơ�>�����S�w=��=�>���=�f���o����o����V��f>���>M;|>����'>ˢ�jz�md>�UQ��ƺ��T���G�N�1�/v��>�K?��?�`�=���V���{)f�Q)?�^<?�(M?e�?H�=!�۾9):���J��;��ȟ>p֣<H	�U���:	��N;�N�:�s>8���7㑾&��>��	��:⾦Qd�i�;������;��d�=�S�4�߾����݈�=�>iȶ�T�G����~���oG?�/�<����/)]�˪Ӿ|V>�Ҧ>��>�`�q�m��\<�k���p�=B��>�w�=�5��n�n�:����l��>"�1?�>3?E��?Z����a�S�N�!�����p>c�9?
��>-��>F�[>C>�>[�f�{���4�W�^��e�>a��>*$g�
"��Ǿ�A��y+����>�#(?����/?̡R?�B�>m�?�<?�>�>Ⱦ�>�3<�~�̾��#?�0?Z@=;���)O��J�m�T���>fv;?����>:`?��?�<?Da??�u#>=�R1Q��C�>��>iNK��㫿���>�lI?�A�>�3?| d?ϳ0>�/��������<�y�=*�/?��??�
?���>���>�ޖ����=չ>17f?���?(�l?��=�?�GZ>=�?��=�I�>�Y�>%?k�N?��t?�O?��>�@�<NM��0 齕�w���0;>�M<��O��(:=�8ļ,EV�S��˚K=��<�m	���:��f�_�r�BT���H?����>.@s>�_��v�0>#�ž/C��u�=>CZ�������Y��.�7�;N�=�,|>�� ?�	�>�)&��߉=��>(�>č���(?q�?�?�<фb�[�۾f L�,&�>�B?�r�=�<l� ����7s�_p=o?��_?�7[�8���i�b?��]?�i�J=�2�þ��b�����O?d�
?m�G�2��>��~?S�q?���>��e��4n�d��Cb�4�j����=/p�>uU��d��@�>Q�7?E�>�b>.5�=Cz۾��w�r��C?f�?� �?���?�3*>�n��1�O���M���]^?���>٦�3#?����ϾH������w/�lV��v���U��"M��v�#��	��x�ӽ�ļ=��?�Fs?��p?"`?n���c�I^�
���lV�r���.�E��:E�L�C�5n�W�tL��掙�\�C=�8���E�p{�?��?a��f�?wf��b�s�Ⱦ஌>�S��uԼ��i>cx���X=���=#`��\~��B�����?� ?��a>�Z?Y�r��r.��\>�A�:������0�>�E�>�b&>,�p>���B=�Ê.�hTǾ�ײ�.Z��;v>yc?G�K?��n?�D�? 1�X��:�!�i�/��R��y�B>�Q>���>JW�5v�(&�jC>���r�.��n�����	���~=x�2?K,�>=��>�G�?�?y	��u��=ix��}1�C �<�,�>1i?�3�>0�>��Ͻ)� ����>�-l?{��>A�>K犾.!!��{�i�ƽ���>�o�>��>�<q>F/.�(\�!M��o3��d38��`�=Jdh?H
���`��>�XQ?���:�S<{�>�hs���!�)�񾩬#�:>�R??��=
�8>X?ľU���Sz����)??�?7���0*�r�~>�""?I�>��>���?{p�>��¾\Tں?9�^?OJ?�8A?���>��=@O��m�Ƚ�&��"+=虇>��Z>0zj=^��=����\�و��H=�	�=��Լ�Q��g��;8����Y<��<�}3>L�Ŀm�F�q׾��� �����vR�w�>vB��p��*����Ӹ�-/���+��6<�^%�|�ܼ��ཧ@M���@}��?K���)��������.��"� ��>�����X+=�p��Xŝ��FҾ̿�_L��rV������ϋ���L��.?�7��sƿ"�������?�K?&��?�ʾ! -��)N�{�>j>'��Ä��]��B�˿�q��(_?�f�>�����Խo%�>:��>a�>�LJ>5?W������5��G�>��+?~?\��ɿ�㭿�ڔ=�h�?6�@�PA?��(�5�"L=�B�>�l	???>2���㦰�){�>��?݊?�kK=w�W� ��ֿd?I�'<�DF�=;�����=Ħ=b=����%K>���>jW�
B�ؽ8�3>��>j������8^�2��<_�[>Sֽ���5Մ?,{\��f���/��T��U>��T?�*�>R:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�鉤�{���&V�}��=[��>c�>,������O��I��U��=� ��~ƿ�����W<��=���]\7��)��d����(|��qL�J5�W۱=��>{��>oˬ>���>nM>�$j?�	`?Oo�>�OK>M�ȉ��I���s>�;���X1�_dy�fpO������K����#N�l��=���2���o7���=k>S�]6���b(�w2a�ӀO�ۈ3?��=�.�� �M�����@2žra���Bݼ�_��[�ʾ~�2��"j�Ǳ�?ӖE?�>���Y�{��]?��E-��I?�."��#��񛰾���=ټ�f�<���>�M�m���:�t�N��1?��?�x����\���4>?��I�|��?) ?��^<Co>��?S��� z��>;/�=�'�>��>�4W>G�������߻?c�a?dn��{����l>4���x���!�=s�p>'!f���ԽZm�>P3C=�PQ�1v�=�>;���$�}W?��>c*���� Ȑ��T��W<=�x? �?I�>�Bj?p�B?I��<�d��>IT�����s=9W?��h?��>�F���4Ͼj ��h5?ڣd?,�N>p�e����t//����1�?)?n?��?�t���#}�~���$N��J7?��v?s^�xs�����L�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?{�;<��V��=�;?l\�>��O��>ƾ�z������,�q=�"�>���ev����R,�f�8?ݠ�?���>��������>縑��c�?��?u���,��=����3l�a���%y>e6,=�4һo��<�7�jK"�����3}��*��1z�����>yM@�[����?�|��%.�x\ʿ���M�������&?	��>$�m�������?��c�c2�Y:N������U�>�>lj��^��A�{��d;����j	�>���<�>%�S�"��1�����/<��>�f�>ni�>ݯ������ę?�U��w<οT��������X?l�?�]�?j? �8<y�v���z��� 1G?Hus?��Y?��'�,/]���6���f?�8Ծ��p��*O�XgJ��#A>;� ?�e�>[��)���W���=?�gM>�*F��B��L���1Y����?��?�����?��?e�.?T#�yǚ��ɐ�Q�-���I��/N?���>����X�T�Y&��E경ћ#?�G"?��[��	U�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?-�>��?W��=7��>K��=�M��h�ϼ��>���=�&���?��J?.�>"I�=;�?�L(��SC��FS��$�`�J��ݕ>��h?WL?N�>�q���yؼ��Y���--��>D�X$�^K�;���"�$>�+d>��->��A�d ̾��?Uq��ؿNj���q'�>54?c��>T�?R����t�����<_?�}�>�7�,���&��7Q����?�G�?�?H�׾�>̼�>Z�>�G�>��Խ\�������7>E�B?��6D���o��>d��?w�@�Ԯ?�i��	?���P��Va~����7�c��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*�hֿ����_N��R������=���=�2>��ٽ_�=��7=�8��=����=��> �d>Mq>n(O>�a;>�)>���J�!�r��P���Q�C�������Z�>�� Xv�Wz� 4������q?���3ý�x���Q��1&�<?`��u>%�Z?CNG?u]x?�d�>I����6�=/��{��=�&��(W�=>I>h\?a�Y?g�-?��=��M��tj�v��^��� Lz�n�>�D{>
2�>_,�>��>S�(=^p>�
�=�Q><�>��h=D��<!��L�B>��>���>C�>E�G>�0:>ȫ�����z�������2����?IBѾ�0�}��{�����$�?,?^<=��r�Ϳ���\�[?�ʓ�2��w�]���=�l-?�y{?;4�=,�����w�=������I��>�ǽ����LM�T�4>�?p�f>O�w>��2��8�.�O����t6~>��4?p㷾4d8�̒u�6I�	P޾��K>P־>n=(����O����~�0!i���y=�:?b>?�<������
v����e�S>E#]>�r=c��=��L>H�c�o2Ƚ��I��,5=dr�=yt^>V`?��">q�V=�Ү>�	��{�T�W��>��>.V>~'7?I�?놝����䕾a>��Z?>���>�w>? >ZX����=1��>%|>$����������G*�BT$>�X��
������]�==x<�}D�=+��==c�Y�2��q=�~?���)䈿��)e���lD?R+? �=�F<��"�E ���H��F�?q�@m�?��	��V�@�?�@�?��/��=
}�>׫>�ξ�L��?��Ž+Ǣ�̔	�/)#�iS�?��?��/�[ʋ�<l��6>�^%?��Ӿ�v�>cQ*�뚜�q0��cv��o�W=���>�\?��ݾ�����,��h?��?%�%M��	�ȿiY��T��>���?���?�0}�$|��(z,��?�o�?��R?aЊ>�Џ��̾�>�yY?z/b?���>�5�s�P���?{��?,��?�I>b��?#�s?�d�>�	x�GU/��4������`{=^;L\�>SP>����hF��Փ��e���j������a>z�$=��>>G�92���=8����B����f����>�,q>��I>EP�>�� ?W�>)��>�/=X[���߀�ԯ����I?��?���W^� ��<	x =:���X�>|a9?g[D<s�Ǿ�R�>�hV?�/�?#a? $�>���i������������<�<>��>(��>��ɼm�W>t�澙�p����>�}�>���i���	���>�e?���>�'�=˝ ?C�#?�0j>��>0dE��/����E�
p�>��>�:?L�~?��?gι�IU3�Q��}桿�s[��	N>M�x?�M?��>���� s����G��DJ��p��n��?`g?&�?�(�?Y�??�A?1je>���*�׾=���W�>� ?����c�>���$�����	?�`?���>�С�����߃����=)����?�!Z?&?q.�hIc���Ⱦ	�<�{I�zݦ��:��ż��$>r�>���1��=�`>��=��n���8����.��=߀�>���=�!6��L~�-=,?�G�\ۃ���=��r�xD�y�>�HL>��i�^?�k=���{�����x��Z	U�� �? �?8k�?
��0�h��$=?��?Z	?s"�>HJ��}޾;��`Sw�|}x��v���>n��>�l�"�Ϗ������YF��I�Ž{4彲X@?h?���>�9?Cb)?~@?��ľ�cw������������M�,���f2�����Dz��%��hG8��9�� ���;�>PG�>>Z �>c�A>��c>G��>(>M
M>tz>YE�>�tj>+Jk>�K�=C�>Br<?�}�}RR?�/����'�L'�w����,B?Bd?|��>��d����k��إ?'��?!G�?��t>G�h��K+�=f?���>���<;
?��9=���	q�<�2�����Dȇ��Z�K�>��ֽ�:�X�L�.�f�5+
?E?���j̾28սm ��Q2q=��?��(?�)�̘Q��o���W��R����7eh�������$�Q�p�K׏��I�� ����(��&=~*?zڈ?����p���� k���>���f>H��>bɕ>��>M�I>o�	�P�1�?2^�{�'�e����R�>[~{?��X>ZX?�U?��y?��]?��>(O�>�戾�@�>�R�ᝣ>Н>�w�>DZ6?�<?�K?�E=?��A>Fu��&���׾�(?Gz?�&?�>�&�>c��K�q ��1���N0��+>��h=!|N���齙����>��>e34?�ӄ���/��
�f	<?��>J��>�H>E��</I����g�>y�=yv����W��F����Ao�>@��?��FkR�DJ>�ݑ=��>c�1=c=�7�u,�=gd�������"=\���N��W�=��0=�C����=��Z>���>�?�]�>�"�>X��$� ����%�=~Y>Z-S>��>�4پ�t��[����g���x>k�?	_�?[�e=#`�=�f�=Vz���:��p������B�<z�?�=#?�$T?+��?n�=?6n#?p�>H��N��QM���4�?F,?��>���{�ʾc쨿K�3���?B`? :a����#9)��¾��ԽN�>�]/��)~����(D��������<t�����?<��?��@��6��k�޸��=X��D�C?S�>�`�>�$�>��)�n�g��$��/;>��>~R?���>rz3?o?IȆ?�L�����6_��H Y�T��>�M�>�J?xFa?)h?9��?A??/�C>�X<&/��SN�qf���8��UV�I�l����>�l&>�!�>òD> ��=���M���Od���h����>@
�>A�v>4�>�h=32-���G?� �>�U������Ť�����Ou>��[u??�+?�=?���E�^)���U�>�e�?p�?�*?�>T�(��=�-׼�߶��r�I��>���>^@�>�G�=kE=yV>���>A}�>U�x�#�8�>QN���?uF?��=I�ſB�q���p�̗���`<>���� e��O��J�Z�rn�=]���z}�༩���[��ˠ�ڞ���ĵ�ȑ��d�{����>pޅ=��=w�="��<�ʼ��<2�L=1ˍ<�?=G9o�R�m<Ql8���λQc���� ���\<�I=��߻��˾7�}?�:I?�+?��C?�Zy>Gv>Hn/���>�M���/?ϝV>�uN�(���D&<��������ؾ�9׾}d����>�K��>�A3>��=뫉<�G�=�r=���=�B�/�=W��= )�=���=��=C*>�>�6w?X�������4Q��Z罥�:?�8�>d{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>t��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>۶9>��>+eR�|1�E�\�9�a�C�[�i�?i:���ʾ�s�>d;�=�߾�Ǿ1"=&3>�d=0��K�[��m�=�V��@�9=D^f=� �>ƵC>bz�=�y��#ȵ=\?=)��=�FN>훔�E@�ݟD�^�#=���=шa>@�+>A��>0�?O�/?~�d?��>o�o�ϾJ=����>���=i;�>�j�==B>�߸>�18?�}D?�K?��>[�=�r�>&��>B�,�@�l��^徍꨾q�<�e�?�?₷>�g<�?�!Q�}n=�ý*�?ss1?5�?6B�>*���ݿ\�5��S�����9�>7�m3���>�*#�q�Z��>��?�� ?]4?�?��>A�=��>)=#X�;�7>y"��O$P=��̽|�3>#�&<Y����֛��}͙=إw��>ɼ!�<s�<��$>ޡ���?0>0q�>d��=���>�OZ>�D��I0>�m;�G���=�N�/�A��#}�p�dZ��h ��ߚ=�!>V��2Ŏ�	Z!?���>@dX<V,�?�>�?�A�>,b���A�5)��D.���?��=��`>
�ý"w��;;U�Хa��]оz�>U�>�i>Z�]>��+�"/S��J�o[ʾ�.�5'�>ť$������0�F�O�����B�����f��޷�	�?�����>!��?ܯZ?ǵ�?*m�>����Ǿ�&6>�z��ָ<|����(zH=�?X�Z? '?0��k�g��D̾����۷>�@I���O�������0��&��ʷ���>������о3$3�qg������5�B��Ir��>��O?��?�?b�W��LSO�����2���q?}g?��>�H?�@?~���v�p���e�=��n?���?U<�?�>$k���j�=V�-?�,�>#N�?�Ey?3�o?�#۽D}�>&�>�0�>ݲf��9>ۮ�=->ݖ
>�5-?�?@�?l�!�.���\ ��$��
_���M�db�@]�=�3�>���>z�>j}�>�֋>�P�>�y�>c��> �7>H��>﬊>o���_���}�]?ny���.�>_�?
U�>
cU>>k��U置�7����=���>z驽+H����<N^|�S�>M�=B��>>�տ0ލ?˽�:�	�K�>?-��A�Ǿ\JD>�U>�O����>��=>�"~>mg?Kđ>�D�=D�>uՒ<Oc\�j�c>L���(��W>��0*�v%ʾk�A=^~��9a��;�������'T�}aؾF,
��*\�(DV�P!<��］��}?�L��N�����f���9�>s?NI?DU�sA��>z?� �>�����ܙ��1��>�¾��?�g�?�4c>9�>�W?ט?n\1�v�2��XZ���u�7)A���d�ɫ`�����Ǡ���
�Ŀ���_?��x?�WA?R�<�z>뙀?&�%�k���#�>z'/�@&;���<=.�>�/��}�`�ċӾ�þ��F>x�o?Y$�?[[?�OV����m<=>�D?~�?�~?T�-?<&5?6$�e�?׍�>B�0?�3?��:?�m1?:?3sN>8>mP�=ڝ�=.����k��J���<3�=�I =�:j��ں&�X<����	ʻ��m�;έ'=��:�='w<TIB=�=���>6�d?�>�c�>�F<?����%/��<��zi?��=�n��D����q����=��a?g3�?τ7?�B >x�A��[��>]�T>��=7Ry>�ѵ>�׽Bu9�ӫj=@��=��>�~�=��ӽw ������B���K$=pS>=\�>�ʸ>A�����G> ��8V��"�A=0벾��������>F(����.D���:�>�A?*C"?ڛ=����g���a���#?��2?+?�w?�`�>�0��J-�!ST�@����J>��w�Gt�կ�O`�����f}�P�)>]�B��D��Q�l>���,aھ�Vk�S�D�|c��ث<�3�'��=s�
��S׾N􀾽5�=�{>�빾�"�>��o�����H?;OK=P����+`������>���>��>��G�=@l�W\=�\��}&�=_��>"# >�9�T���MB�Hf����>��A?*[[?R�?g����%t�D?D��"���t��YD���?�ɮ>6?�E>ɝ�=ló�����`��aE���>�?�>*����?����F��"�#����>d�
?��>�?�?T?T�?�?e?�.?Q�?�H�>����Ȓ��{�&?�5}?��%=<`=;����H��I����>I 9?�������>�?��&?��H?��k?lv?ǩL>��^�kf>Ha�>�N�,����]>*2H?��>��,?|�V?��U>�k7���ckF����=m>_�(?}%?�C�>Ǧs>���>����z��=��>ـc??u�?nOn?�.�=	�?��.>�\�>	�=�ȩ>D?�>Zj?[�O?]]w?��K?���>�U�<"���+��=`k�FWn�m<-�<�~T=sm)��sC��+	����<�m<����D�.����,��M����#2<�i�>�Qt>ퟕ���1>��ľ�􈾒-A>{������d��7:�٣�=K�>��?���>�z"�ނ�=K�>.��>J���.(?,�?��?�>;
Pb�/�ھ��L�� �>��A?��=�l�#M��A2u�
�i=Ьm?�t^?l�X�ո����b?f�]?E󾸸<�0
ľΰc���龖�O?x?�KG��:�>��~?�r?��>�e�(n��ꜿ�%b�^Uk�8U�=>�E���d��F�>�7?�I�>��b>U�=�>۾#�w�����~?n�?E�?q��?�E*>Z�n�q:���9���*�j?���>G����?sӼ�$��㖾R�I�����x�I���X+��Sâ��[`������p����=ˣ?d$|?��S?&ie?L��;�U�jGd����Ѹd�H'��D!���_���V�{!I�&�o�? �}��"�Q�ͳ���<e�?�O�6��?>�?P׽�j�>��V� Ѿ2ܸ��rV>�g��(~��Q�=`�(HA="#>�T�aa���)��|�?�}�>n��> ??_`��dA�:T1�=�?�����e>�hd>��a>�^�>|PL��6���	�������V��<v>�xc?��K?��n?�m�R&1�Ӆ��ڠ!��/��S����B>�\>��>޶W���'3&��V>���r�c���u����	���~=֩2?�%�>���>�M�?�?�{	��f��Dgx���1�S�<�$�>:i?�7�>ކ>��Ͻ�� ����>�l?�w�>��>zǌ��k!�X�{�
!ʽ�!�>ǭ>��>�o>]�,�F0\�e��i}���9���=k�h?���Xt`��ׅ>_R?� �:��J<�T�>\x�$�!�x����'��o>�~?Cu�=��;>�Fžp'�q�{�{@��;')?(�?�(��M�"���n>?�8�>J�>V��?s��>�?��@����R?zea?�8N?�@?���>��<v���
�ɽL\$�| 
=��>t%\>��=��=X#��+]���S==��=dhg��4�[<'ڃ��8;�%
=^6>N�ڿ��>�M>Ⱦ�������V���~žI}:�r~����D���¾넼�vy���)T�ŬA���ͽ�xi���$�EAn� �?���?����������T�p���m��>ҏ��ὁ放�֚�W���ɾ��X��H��n��W���i�
c*?�� eϿ�!��ɒ��*0?�d?�y?��̾F�X���+��^�>V>�n�D�"�[w��w�ֿך'�XK?�b	?KT&�k��&��>Lw�>���>��N>��)*���`/�j/?�w?}��>�\��ˬ�f���U�?=��?H#�?�aA?�?)��J�	�T=Y��>^d	?
@>��/�P��������>�8�?�Ǌ?�K=�vW����?e?} <~nF��o̻t��=��=�=�a��5I>��>��
�B���ڽ�3>k�>�'����T3^�E:�<��]>�lԽ���4Մ?({\��f���/��T�� U>��T?�*�>Y:�=��,?W7H�`}Ͽ�\��*a?�0�?���?$�(?>ۿ��ؚ>��ܾ��M?^D6?���>�d&��t�օ�=�6�A���w���&V�r��=U��>c�>ǂ,�ߋ���O�J��J��=���)�¿�����/����=��=��f!"���T���= ���ds���y���;!=z�>:��>��>��x=97>�-b?��f?��>�ٚ>����<B�JN�upS�ߧ����޿�X������b-��y������߾h���D�����=���=�+e������*�E�N�g�d��G&?���=�Ǿ�$>�ܴp�}����#C=gX0�܈¾��+��Dk�0��?�C?��k;}�����%��#�}�O"l?¯&�o�ľ�ǥ�O��>�A>Gh�=���>%��n/��zS��]G���1?�?�3��B����/">1S����<�)?i?���;�d�> �#?��:�s�k�Q>�6+>`z�>��>�>����d�۽�o?-�S?����䘾�ˋ>�#��d�����9=��>��K�������W>}<�򂾄;���C��p�V<+@X?ñT>]�9B��!��r��,��;��x?{J?tHf>��Y?^A? 6��)0�,�L� ���Re=ϘZ?�Zg?>��Q�cB��m���6+4?�[?_9Q>��r��\о��-�:�*��M?�f?X��>�%=<~�g��d�������2?��v?s^�ws�����S�V�`=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�#Þ?��@���?��;< �X��=�;?k\�>��O��>ƾ�z������ �q=�"�>���~ev����	R,�e�8?ܠ�?���>��������
>�L���A�?�$x?W��Z^�<���m�e��l�>��;���:��ռ�N��q�6�����2�8�@� ���ϗ>h<@JpѾM��>3�����ڿw@ҿ~`����ž�F+���?N�$>�������s�a�>"��*�R��HS��8���`�>�>���ȑ�h�{��l;��ġ���>$��,�>�8S�����󃟾�&5<�>m��>���>e���佾1��?p��>+ο���������X?�V�?�x�?�?�6<~Fv�t�z�̗�#BG?�ss?��Y?2v#�]�i6�x�g?3
�l�q���2�f�kX�=KA?lN?T��H�o<��O>3�?�y�>�	)�w}��m�,"�5�?���?���$�
?�;�?D#V?�=2�Uի��떾����(e�m?�L�>t��=*��y$�MA��s�*?w'?4�ݽ=m>�]�_?*�a�N�p���-���ƽ�ۡ>�0�f\�#N�����Xe����@y����?N^�?i�?ص�� #�f6%?�>e����8Ǿ��<���>�(�>*N>[H_���u>����:�	i	>���?�~�?Oj?���� ����U>
�}?�m�> �?���=���>��>����<��@>(��=f����� ?�L?��>jǳ=�GV��2��oI�9KM��}�JVJ�X��>��]?��F?$v|>���R�G� �;��[#�6���c;�lF��;���!>�55>B>$�:���˾�? ?�"���ؿ�����*���5?KC�>�]?�����߃�k|��|`?x�>k�����������\�??�?��?Y�Ҿ����">YV�>��s>ȿ��	�������(�N>k??��{$��0�m�H�>3P�?(�@�c�?Peb��	?���P��Ua~����7�a��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>!�l?��o�P�B���1=8M�>Μk?�s?�Qo���h�B>��?"������L��f?�
@u@`�^?*�hֿ����]N��P�����=���=Ն2> �ٽ2_�=��7=��8�/=�����=s�>��d>"q>=(O>a;>��)>���Q�!�r��\���S�C�������Z�B��Xv�Wz��3�������?���3ý�x���Q�2&�$?`�$��=Jmf?h�=?�2x?���>����=�+�?^�=��Ǽ(�s=2�=*T�>�b?&�2?��v>��O����0��� ξ₾<1�>Dk�>��?O4�>��W>�Y�=S@>R:J=��O>ۙ
>�S>����y��<�`�>5M�>V?h�>��.>�*>m��t۴�/�i��4}�u\��o�?ux��^�C�R����� ��>ʑ=��*?Ђ�=�����oϿ_���+US?�o�����D��C�=�-?ƍ^?t6'>�⣾�0I�ŗ�=�J���.c���>f�0�"%��{�2�*A<>�w?��\>���>�1%�fe/�<C�m������>�?���e�5�0_l��'I�������D>�2�>�)�<�q��5����{��~��=D�5?;�?�����¾�ҕ�D)���W�>u�g>hc�<O*�=<>����˽��7����=�Ӄ=�*>��?$ �<��&=���>��վ�7��ryB>�'�>g��>�M?ν*?��\=ڟ��K��j�m�U��<l��>�C�>�t>W�?�^�=���>��]>.b =�3��B����9P>��d�}c��oK��=e=���(�=�8"=���!��B��=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ~9�>+� ������ w���8=���>aNH?YW�|v�D���
?EF?=t𾖡��X�ȿ�x��a�>��?6 �?�}o��㙿��=���>[�?=pY?�i>�GپG�c�k��>��>?��P?�>�>9�x�0�i?�ն?��?jI>���?/�s?�k�>40x��Y/�i6��:���
o=	7\;�c�>"V>�����gF�;ד�h��W�j������a>a�$=�>F��4���6�=틽�G��{�f�<��>�,q>3�I>nV�>�� ?\`�>1��>;p=�s��E��������nI?��?5�b5U���2���C<y��N^�>��4?O�e=�¾�>�>�W?���?��f?$��>U���x���Ŀ�ױ�E��<�t8>���>��>7�,�7@>:�ܾ�_�!(�>�]�>I'�ބ�Jǎ��d���%�>�?|i�>'=�=`�&?f)?B��=���>T�F#����J�[�>���>��?��?�?������O;��`����H��c>άQ?C?�c	>㲃�a�x�ǽ� �����d�?��?zK�3fC?#ڎ?��7?$�u?S'�>�Jh�败��	���e�>�?���.�/�������^	?&?D��>��I��������k+��2���>��W?�f$?@�
��Ec�0�ʾ���:�/;%�<��߼*����<>���=V-��)q�=��M>��>íN�a�[���'����=K��>�=��L�#�e��<,?Q�L��􃾗8�=��r�(�D�/|>�tL>������^?�<���{�/����o����U�~ۍ?��?�f�?J�����h��,=?��?�?�c�>����{޾u��~�w��x��h�<�>���>��j���侙w��ߎ���H��7�ƽu0�<*?H�>e9�>�2?Jn? 6?Fg��\y�6�W6*�,͋�bH��+Ҿw���<6z������Z�u��=1���=
�K>�������>�\�>�RK>r3
>��Z>��=�>�۾=�4/=��>�#|>@�[>Mx�=A�1�/zq��BR?������'����Bf��V@B?��d?_��>SYk�����V��KR?0m�?�k�?[�u>h}h��+�[o?lP�>a"���k
?�:=RL�ZX�<�7��}�����#j��r�>��׽��9���L��f� o
?�4?�q���̾��׽a����d=�?Ez"?7�-��I�(�n� �`���N�%D=B�y�{|������"p�FԌ��x|�� ���X��'�7�-?�?+2��¾�=ž8kt�fxF��Hx>�?�>V��>ΏL>�$�����[G� �7��/l��m�>�^z?g�c>-!T?�B?�
`?�-Y?�U�>�˞>*���,��>3V󼯤�>=�>M?ƞ)?�g,?��'?g7?�1�=G��$��`�ھ�?;?[�$?Mv ?��>��;��鰽5����d ��y����a:F�<��=�������9	�=J�>�N-?a
����"�Bk ����=��?�>MX�>hw�|�Ǿ��L�; ?+��>����
 � み�� �?�>&ي?~�����@1>�~�=t�=n=$��=�Q�c}=�5�=�)�m�|��>����9�	=n�>8i{=O롽3- > ��>�?&<�>�0�>3����� �.��B�=zY>G�S>�>�پ�{������g�#�x>�K�?b�?[g=�O�=���=35���9��{�+���*`�<,?y_#?7�S?鞒?N�=?� #?�>�V�EX����0�����?!,?��>���²ʾ�!�3�7�?MZ?�<a����:)���¾\ս�>	[/�	.~�K��ID�������}�����?���?+A�>�6��y�}���TY��H�C?�!�>8Y�>9�>`�)���g��$�:4;>{��>R?:�>�l)?D�*?&e�?׶�Ty��	����^�G�>��>P�E?kUS?��?u|�?��:?��5>�7	>,�侴�F�?=˽�[�<��Z���D<�1r>�B�>��>���=�=!��((P�8�����T=ջ5>t�?q��>�,�>�ty=�/����G?F��>�F��;{��褾�̃��G>�Bnu?X��?p}+?�=�m���E�Wy���>�>�Z�?��?*?�S����=vD׼�ն���q�R�>!ع>��>NN�=*GD=�>w��>cI�>���Z��n8�0zL��?�F?k��=<�ſڍq�IVp�M����d<	!���Be�������Y�$�=Oߘ�m��㩾�\�I���2k��d���bn����z�g��>r$�=e~�=:��=���<�GǼv	�<��H=���<]�=arq���^<�7�ȊڻR���vvºn�X<�rH=0N���پ�|?��:?�~#?��M?�I@>�N>���=U��>g���\�?�q>h���r���:������oh���ľθ�g���uz���8(>'0��*h>��3>C/�;>��<��1>a��=rՇ=�_>�x]H=���=?�2=���=:">�I>s">�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�;>�>��Q��@0�L^�Υd��^\�:� ?�-9�W=̾���>[3�=��l!ɾU+=�2>��^=N<�$DZ�Tș=��{��==�i=��>�D>\̺=ư����=�A=��=��L>D�^�[I��/��8=�5�=0�a>�7'>��>��?��/?�ld?,\�>�&o��zϾΠ��G��>Lm�=�[�>Ë�=�2C>#)�>�h8?~�D?�K?1j�>*߂=f_�>H�>l,�xm����Z���G�<�0�?�r�?���>��F<<sB�8���&>��Ľ�9?7�0?�?-�>���ܿ��4�YO�����<B��1=���F����=�_��
f����>��>d�>]��>�g�>��=�,/>5y�>��=N0U=_m|=E	�=�'�= '�[.>���ѝ�=�����O�`s�=��׽	��������s=#D�r��<��D>zd�>H��=���>��=�G���/v><���OY����<S:���B:���,�v�X���=����\�g;2��>�,�=U7���A*?9�Y>��=C��?}s?���>N�Ƚ�� ΐ� ����N�=��>*���)w�ԗ7��:�~$�����>3|>��>÷t>�52�aF��I[=�˾�Q0��\�>�~\�D�V����3�l�����~���d�4=:P??���Q�">�v?�D?Rc�?���>�i��Uھai�=�;�����<��W�L�"#J���?Ƥ?�o�>�_��IA���ľ4ý�F�>�
F�I�P�� ����.��>-��賾���>�d����;�4��ą�Y��^B���u���>�N?�I�?p@s��l~�}TM�p�����]� ?�Bl?�ɤ>G�?QB	?g���R�B�n��=�Gg?���?���?��>��ｨ��=/[?%�>��?��?��Q?]%�Z�>y��(�>�ݪ����=��">��J>�V>��"?0� ?,	?~�T�y=�.;ľo/����� ���I��<5Y�>��>���>�>��z>��>'�<>���>�)�=1�A>���>J�r>�߷����?�<?�//����>�),?�C�>���>���<�/���!�:���=F>yQ��.��햂=�p�~�J>^>Ex�>Oп*��?�=�����?'��3� �nƃ>[s�>�E���?��>�}�>��?H�?)�K>.1�>δ$<��n��GU>��,�!�'��yE��*��eϾ5V=����P=A���9���o�D�8��w[¾�lI��t��D55��z�����?��;�RE�.l��̧�v�>��?��S?��ս��-�XT>�
?���=����{������&Ͼ�h�?��?�d>О>�W?��?�(1�r2�|)Z�ږu���@�x�d��`�Gʍ������
�������_?��x?��@?0I�<��x>�{�?D�%��ώ��C�>�.��;���7=c"�>/���6�`��UԾPþ8��\�D>�Oo?��??(?��V��[���{>m�X?1i�>��q?̠?�B ?7<gN<?w(,=��%?ֵ?�=U?<Z�>� ?��>���>��=J�q>�V����6��|��\<?�^>X4>���#�.��tϼ7����/���Y=��=�Q��_
��:�>�l>�V>Α,>��X?HW?�H>��4?�xP��"/�����KVB?[>���*81�[�����h>�n?9�?�QJ?tP>�'6�2�7�̔�=�i>7v�=��(>�`�>J�����Iᶼ�g>�v>æ>��z��8�Ⱦ.r���u�d�3>���>��>v���w>S����S@�$Q�=��۾�+��gi��`0�Z�"�u���Q��>��_?Tv&?��=����.�� Z��?'�"?�(?�Hq?�`>�v��?�:�֞D����&�>��<��^"������Q �r����t>�cL��t����f>���Ҿe�k���L�s��A8=�D	�V<�=�<�;ھW%����
>� >Z0���� �Z������<&H?˩a=9C��o�O�r\��� >��>F��>�9-�Q�l�f1?�F��	��=Z0�>��7>�����J�7E�n��.C�>ɞ7?��5?E�?�����n���W�/���>���\>?�ݴ>_u?�<�>��J>	�\�G�	���[��8`��B�>���>/�d��VѾ𲒾T.5��2�)�>�S?F��=�S6?��`?��%?/ڇ?�2�?��?�g�>�J2���оk*?��|?(�?�;�<V�q��c;�� O�͛�>-#-?��\�P��>UB�>��?ϵ:?��e?�4?���=��:�U�j!�>��>$$B��ۯ�`d\>��T?� �>Q�:?q�]?�p>R%�c|���ݮ��!��=[=0?��1?Ig?�+�>�O>DS�h��>�>��e?\�b?^�n?��&>2l�>�h�=4�?3�>/��>xR�><]?�f?�ۅ?�SU?���>��=H&߽i��'��Z���U?=���<b-/�]�2 �]~��э��ev�_H�=ɲY���g²�1��������>Ϣ�>�[Y�x�>�Y|��_���ӓ>q�!��Gྰ%����!�ѕ�/S�=60?;�>,i���>��>�h�>��*��I??�0?]����y�!��[�N��>#_M?��v>�=�f���y�Q�"��=R�?�]�?�ȗ���=�b?��]?�h��=�[�þ�b�C��y�O?��
?O�G���>��~?{�q?3��>��e�9n����Db���j��϶=r�>UX���d��?�>��7?*M�>��b>�(�=�u۾��w��q��<?��?:�?<��?<+*>t�n��3࿻O�����n?��>�i��4�?��<�Lž)����啾�� �_3��MP��aF��Rޤ����P����9��:K�=��?�y?��i?��j?l��b�R�*b�ܙ���W�����2�0<U�vpK��6�ra��������c����h�̢[��oS��y�?uc?���2��>?�m��x߾h<�\<>c�Ծ/6��m�=�2��T	�<���=�t��:���v��m�?��>�ڼ>�uS?PXq��z'���;�n[�GA�y�>�F�>��=��>�b=���fY��+[־@f���:K��Wv>&sc?�zK?��n?�b�(<1�܍���!���.��5���B>�.>���>�W�0�-&��T>��r�����k��H�	���~=�2?��>~��>G�?C�?Vt	��W���rx���1���<�-�>�i?�2�>[Ն>M	н,� �7��>��k?1�>�ݠ>]u��r;!�Z�{�T0̽%x�>�Y�>w��>��o>Xk1���\�S���\��-U8� ��=�Ni?܌���z_�t��>1\Q?��:4�E<��>�����!�j4�9�'���>��?���=O�;>'ƾ��
�{�e2��o�)?�?������'�+�{>(}!?��>X�>��?+w�>��ľ�)9��?�\?�J?5�A?��>�!{<�uڽ�ǽ@�$�:}4=Hix>�t_>t��=-��=t��[^�
��a.=h޵=#���R�H8������j <#<=�A>�Mտ̜D�����(m���d��Jbþ�����5�ȽH*��;���7�A]�Gz)��ۧ��s#�恄�O/}�J��?o��?���bkܾ�Ԏ�Bnw��y�b�>zr����ͽ&|¾*ċ�ۄ���|��\ �Q7���j�����J[���2?f`�`&ԿE����!���I?'%+?")f?ex���A��[�iߘ>途>)�����"��Χ��Nؿ+���AkS?gV?X�9���=.D�>ǋ�> s�>�z>��A�Ќ!�yhg���>rW9?' 9?��������ȼ������n�?#�@�A?$�(����{V=X��>�f	?��?> _1���f���:�>�#�?�Ɗ?n�J=?�W�_��ee?���;�F���޻���=_ �=��=���fJ>�U�>eT�y�A�7�ܽ��4>���>�M%��-��^��.�<gL]>M4ս����4Մ?#{\��f���/��T��	U>��T?�*�>]:�=��,?X7H�_}Ͽ�\��*a?�0�?���?%�(?Eۿ��ؚ>��ܾ��M?^D6?���>�d&��t����=�6�׊��r���&V�v��=Q��>>�>�,�����O��I��u��=߲ ��Ŀ���:�_��<@F����Ͻ�䬽�%׽I�l���3�d�:���in =�b�=;��>?i�>ؘR>]�A>_�[?X�m?�u�>�<>(�Ľf����վ��q;,��w�.�o��p�N�O����A��QS߾)� ��=�5�jjǾ�7�`�>A&Y�#M�����Yc��]�>ED?�2μS��FH��)�-{���yо��<��������R���g��V�?_�U?�����}�ŷ��sa��҄<6V?1�������¾A�9>M0	��->��>�<���*��8b�qiI���2?�F?f跾@b��Xu">���2W�<�'?~j?�̥<3�>��"?q�R�J2��M>��>~v�>��>+�0>1N��5�ʽ>?T�N?�*������z�>�Ǿ���hr=�a>O�F�s�3��([>pA�<�R��s �:У˽���<�\?�� >Cw ���������ѽ�6=�#l?��>���>2p?^76?��|�\ھ�a��(��Z��u�J?�An?���=�Ni��䔾蕾F73?��U?d�o>�F߽��Ӿ�L���/� ?j�^?��>�`��6a��Δ���o�F�*?��v?�r^�=s��U���V�+=�>\�>��>i�9��k�>��>?�
#��G��躿�YY4��?d�@j��? �;<[ ����=d;?U\�>D�O��>ƾ�|�������q=�"�>����eev����FQ,��8?蠃?ڔ�>̔������>=4����?��}?d���5��=���s�}�k���%�=�Jp����4�@�P���3�偱�_�������Sǽ�#�>+�@�ʾ @?m��a'׿P�Կߕ���d��S�˺ֽ3?x>y>�k#���]�]�?��fi��1@���T��@���J�>>�����#����{��e;�)����>/�_
�>.�S����3����5<_��>P��>Et�>gi�� ���6ə?w���:οs�����ҾX?_l�?T\�?u�?�~6<u�v�`�z�vb�w8G?`s?��Y?J�%���\���6�e"k?������d��
4�񆆿{�>ղ\?T�>����G�M%�.�B?��> �W�Hj������۹���?$m�?��־�}?�k�?�R?���(��qC;팾�O���N>?#��>ȕ�ܡ5��w!�xѽ���"?.W ?����BP�E�_?)�a���p���-���ƽ�ء>��0��i\��.��*��2Xe���-Ay���?I^�?��?����#��4%?��>C���9Ǿ�	�<�~�>�(�>*N>�L_��u>@���:��h	>>��?	~�?�i?}��������U>��}?�#�>��?�i�=�a�>�g�=?��
-��n#>��=��>���?�M?BL�>�W�=�8��/��ZF�FR�g$���C�w�>��a?�L?�Nb>���w2�i!�mͽ�b1��m鼝T@��,�Ø߽�*5>��=>�>^�D�1Ӿ�)?�<���ӿ��������IW?��>� ?�3޾�=Ѿ�"��_|?5��>A������Qq���b���]�?��?Y)�>?���my�<c�&>��H>�#N>�A�<!cE�H�Q��dR>�:?X�7�xs����Y�^C�>�b�??N�?X��?��c��	?���P��(a~� ���7����=��7?g0�C�z>���>��=�nv�ۻ��?�s�T��>�B�?�{�?=��>�l?�o�<�B�"�1=M�>��k?�s?_\o�e��B>��?�������K��f?�
@zu@#�^?#��ޔ�������辿�b=��=5��;�U��E%>��=��z���!��2;=���>��S>/��>��>V�>;�=�������᡿� �7��H�c��9T=��⾁o
�7ܾ�0���Ǿ�s�un�̘ �(��H�;�8���m�=��T?�}L?��r?`��>Ѧ���� >���L=�W�z�p=[Mx>��.?��R?/?DΛ=ի��h�g��ӂ�n���� ��ھ>2�D>���>%��>u׮>Q�ջ�8F>)k?>�z>M��=8=����q�<Q>b#�>���>Q�>��7>��f>趻��J���wi���q�Wq
��P�?X�оo�4�_����^��V�ľ�W�=��1?ʳ=�꛿�^ٿ�|���p?��¾c�+�1��J���kL?���?4��:s�콭ꪽDE=,2y=lz�X�>U�|������!�B��>"?z�f>�-u>g�3��V8�I�P�@v���<|>6?4Ͷ���8���u���H��_ݾ]1M>7˾>P�C�"a�������3gi�.){=�k:?w?�A��rװ���u�+7��x2R>#\>@l=gE�=�M>��c�URǽpRH���-=���=r�^>��!?m�<o��=S��>�����E��܄>�Y>,��>_f-??�>��5=Gо�ؾ/_���V=(��>��~>.��>U�B��lU=Hs�>�o >ʏ��i��@��s��Ƈt>���퐾��
�����j��^�=~C�=�⫽X��L>�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ
g�>�)������J����u�[�9=���>�_H?'W��1e�p�A�?�'?�򾪭���Jɿ�w����>e�?j��?�m��m����?��7�>�#�?K�X?#�h>�I۾�*[�궋>��@?�xQ?��>�V���'���?%��?���?� I>���?Q�s?{h�>!0x�7Y/�4��Z�����=�?[;�Q�>kZ>H����kF��Փ��g����j������a>�$=5�>�H��4���4�=����F��k&g��>K%q>��I>N�>�� ?�\�>P��>]0=A_��q뀾���PDL?ɿ�?���2B��2U�iBG=�ǁ�˪�>q�/?�^>��ƾ�|e>�Y?�J{?�Ui?�A�>Y�龢+��VdĿ^ש��k~=�]>t܌>�`�>��=�N�>d;޾��l���><�m>e��#fǾ�۾���r.�>�r%?���>���=�#?��?m�V>�Ұ>d�F�񛐿�B��h�>T��>�$?.��?�Y?�Ⱦ��1��c���Ԣ��T�]YC>Q�u?'Q?��>s���ro��f�����uU��Y�?(c?�����?6@�?@�,?}:C?�^@>�<1���پW\\����>H�"?�����?��#���M/?vA?���>��t�_�ýڜ����������
?�QZ?�#?�_��Ob�����n�<� �?��W^B;4D�҆>��>i���WZ�=ݺ>�	�=�p��:�_�<���=t=�>	�=t�<������<,?�H��ۃ� �=��r�)}D���>�|L>R����^?xG=���{��
���v��~FU����?*��?bf�?�촽��h��#=?s�?q�?=6�>DI����޾���Iw��yx�k��>���>k���供���ꓪ��E��ƽ$6.��0+?#*�>\�?��D?,+
?C ?�/��5y�~�+;��0���k!���CJ!�F��<$���^���<��Ӿ���x�>"���#�>E��>
=s>Q�=B�>��=ߺ�>$�>���>"}�>��>us>�9>uG=M഻�MR?�����'�j���Ȱ��GB?�ud?>+�>E,i�쎅������?���?�^�?��u>Ðh��<+�(u?^r�>���k
?�;=�����<{Z��3���m���=�|��>�ֽ�:��M�~vf��b
?�2?���(e̾�V׽6����a=��?d,(?�*��Q��mn�,W�[Q�|d��,�`������%���o������C/��t(���,=u)*?G	�?�A��뾥ԯ���k��D>�Rt>���>E��>��>#�O>ؘ���.�4�^���(�0���E�>��|?�ց>��L?I~>?R4M?PpN?��>Uˢ>H���YT�>�\���g�>��>A64?�)?��/?�<?�</?�f>���Z� �U"վg�?�?��?���>B��>p4t������C0����|�^��<��5�<�;�<������9�=%�h>�g4?a���J����¾f9 >B?;��>�&�>p��o���K��Pb�>n��>�R��K��9��SE���"?q"�?�I���o�<�O]>H!�=g��=��D=��>E����=uv>�(����=[��=ec}��L>p{�=C>ĳ]=�@�=H�>x�?ᆊ>�D�>cI���� ����c�=�Y>!/S>�.>�9پ����!����g�G!y>4s�?�r�?'%g=	�=)2�=!v���K����O��X�<��?bG#?iAT?U��?W�=?Q#?	�>�.�hL���[��K��c�?�#,?<w�>C����ʾ������3��?qh?bCa�'��01)���¾}ս�]>zl/�"*~���� D�1�������"�����?���?��@�q�6���辦���ce���C?@3�>��>��>�)��g����;>!a�>��Q? ��>�48?? �>q��?m�=,0���¿\������>q��><k?�?�OK?�ĳ??^p?u>J>Ƒ{�8H�y�e�r��'B���c����>�|t> ّ>;C=��<N�~�sc�\b���P��N>	�>��[>�M>cՈ=�{18[�G?ѵ�>������6���/X��C�=���p?��?�
.?-+�<�
��/D�������>BЧ?�C�?d�&?�'[��u�=Px��)͵��sv���>�2�>a�>���=kT>=��>:��>c��>���Ƭ���:��e}��?'F?f%�=?ȿ�tv��m�������D�����FV��ҙ�?-D�5��=��p�]z�~+���J�-m����x�����E�������?w9�=���=c�>�C=*����ZC=ҿ�=�����';J,�O��<�X���iϼp�u�I�@;���<�?=���;Z��[�?�)]?ظ�>|�b?J�>$��=1l�=e�>���.��>&*8>�VA�V�Ҿݜ��gi���s��y�P�c�A�^�O(��:��=gH���=Ss>φ�=���<��C>���=��^8�<��;E->+s=��>��Q=�f>�;+>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�8>��>b�R�`1���\�صb��<Z�ؚ!?[;��$̾�5�>�s�=�y߾��ƾ�+=ρ5>��a=m��\�ߪ�=]M{�~�<=��j=�>��C>׵�=Xү�;
�=>mG=θ�=��O>7����7�6p+�[Z3=��=�b>?e&>L��>,6?/+7?��x?U��>r%����˽��m�N>Ү�=X�?��۽;�G���>٨(? iU?E!{?]`_>�Nd��2�=u�>>����&k��ﰾ�Y�-�Y�(5�?$"�?��>O�q=�P|<-۾�!P��<�?�")?�?T%�>QJ�t�ο����!I��u�� ��/r���C��IV���>I�t>�Ť�U�>t��>�>�>���>A>�>E�<�m<:W�>�2�=/�=�}>2\�=>y�=9�=�К>�c�Y�;l����	�<�a4=��@�����\�>=/r;ãX� ��<��f>���>���=�V�>?��=:���.> �T�}�g����<,��+�K���w��be�M�>��򟾝��=p��=u'<�c����<?fn >�>�a�?��?���>z,��/�33���?����ʾ8ZE>u��>m˄����F�F������m�w��>�i>��|>��p>�PD�k M��v�=�����<���>��l��^��H/�S`v�t̨��ܘ�w�^�� =��6?\=��j�F>��t?��>?���?�0�>@C��;�=%ze�t�=S�'�V�^��=�/?[�?��>�����F���˾����P��>��H�|�O�)���(�0��s������>�r����о�>3�
\��������B���q����>�O?2ٮ?-c��?���O�	��粇�W?��g?,�>��?�r?�U��������[�=^n?���?p5�?gf>��:�b=��?l�>�X�?�t�?ǂY?Eڝ��� ?�`��q>�#s<��>�k_=��=��S>��?��?Y4?�G��D�����|0ھ�.����w���=΄�>r��>�D�>�Wk>g9�=C��=��D>^ԙ>��>n�>�q�>�9>:���%����,?�����>1T?�l�>Gs>r|;�d)W�V�`��P>m'�=��;��?��l�y�*���>���= �>�6ڿ��?�z�=ǒԾ�>�ž�YC�6�H>�����.��M�>.�D>��t><��>��?��2>fp8>�&>[�f�>�r�:�
��R5��.����K=/ m�62�=�zܾ��/��Zz�{r˾x ���_���X�jAA��P�,�?�o¾�$L����4��{ �>�[�>t?�=��׏��˽>,�?x�u��~ľ�楿Kg���%ݾi֓?�*�?�?c>�'�>2�W?.�?v1���2��gZ��u�.+A�r e��`��⍿����4�
�'����_?T�x?[kA?O-�<Dz>x��?�%��ȏ�P�>�&/�r*;� �<=�8�>�����`�Q�Ӿ߰þ�&�SMF>�o?�*�?�M?��V�p������>��n?΀�>��v?�9?Q�6?���=�?(:�=m$?g&�>$M?�z?�m?qv?L�?�>���=�����c��?T�����`��Bɰ<�5�<��5/��8϶=!����ռK�H=�%>�5<��=|t=*�P=X�ż��P>�Yp?}:
?�i>��H?(����C'�����%?ȏ'��Щ���e��{�{_����X>?�_?r�?�9:?�%J>� t�B>���>JAʼ�0m>l�c>��>Ȱ��93��_���R�T�b>�N\>�Ӂ�.;��$��%����=آ�>ax ?y��>���Q�&>i�bZ�c�O>�v������1����G�f�3�tG`��V�>�mI?At?���=�l�e���Z�&w?`2?�<5?�t?wƲ=+�þ+a+��F�sj��T�>��<O��v��MI��Z�F�چ���~�>t�l��x��Qya>=����ݾЫn��lJ�t��J�J=E���W=&��\�Ծ�:~�|�=��>������ �����ת�*�I?H�l=g~���&U��	��0]>Q��>�W�>K9�d�v�y�@�Ӫ��⍗=N%�>3�<>�֒�p��=LG����6�>�3?jR?Z�?��������L�t�⾣�i��փ:�E'?��>�?��~>s'�=4Eܾ����b�~�9��r�>��>h�
��2�xP�������*��V�>�R?G{�=b�?�oW?
?�q?��:?�C�>锡>���^�;T�&?��?�h�=����tZ��f:�^�F�>�>�(,?|�4�+��>�?��?��)?��T?q?��>� �FB���>��>��W��s����`>��K?ȷ�>7R?+$�?�;>/>7��孾fȽS]�=n�>�0?^?&?���>��>$��bz�=�>Ac?��?��o?���=�?��1>$�>Ui�=�ҟ>�t�>�?vO?��s?��J?/�>�<�-������-�q�
�S���M;U�D<�y=e& ��q�X��8��<�N�;�+�������+E��{�����;�j�>*��>\�T���8>A���D&��=[>`���m���!����d��� �g`>g�?d��>p�:�<0�=�t�>���>���;�$?��?Cp?UHB��{Z��oҾ>\��`�>M?�{>�0[�Ӣ��8�j��!>,�z?Po?�0�C�.ca?�U?2���0��ҾH�������6zL?��?�V=��z�>�T�?��n?�?��J��Uq��u��Akc�;<z����=�P�>64��}^�ƻ�>��0?��>=�K>k��=�O־K�w�<6����	?�S�?�j�?M܉?�y/>��l��"῾������h,_?��>�K��uY"?�+�e�оzH���<��H�澙L�������6��ׇ��ڱ"�-���a�н��=h?��p?�Xo?�3`?6g ��`�{�^������S�o$ �C�!%F��XB��@�z0i�� k��L0���3=��E��c=�,x�?�`?��:�U��>-�u����w����>�Ź�����w�~=�;��L��z�t=׉����սѭž�6?�:�>��>3�D?�4a��-��D�gMN���m�>���>�i\>�a�>b��z����_���辐%���ɨ��Aw>4Rc?��J?8�n?�� �Ȗ0��s���E"��)'�����?>�!>ر�>˩Y�Q��&��>���r�x��/���3	�M�|=�X2?��>Γ�>��?�y?z���l��q�y��1���Q<a�>��g?i��>�>iɽm�.@�>1�j?W�>�V�> ˌ�yi ��P{��|ν�)�>j�>,��>BWm>b�3�MS]��ώ��0��B8�W��=)1i?�v���Q^����>��P?���;��<}ܠ>v���_,#��1���O*����=��?5٫=QT7>+ež��o�x�ē��{ ?δ?�L��-�0��D�>�I?C��>�=�>�ƃ?�|�>�!��j�<��?��U?��I?�lE?R�>sB"=mږ���̽�{/��z=�>�mn>�,=˒=RN�M=N��~7���<��=�uG����;<�i:5!Y���;�A3>��ҿ%c9�l�ھߑ�_���gu��_K�����<8�t��-�y*��d����=��ٽ>3�=���H�f��>���A�?��?J��7J�������j��x'��>�i0�q>�������h�)����������,��6V�;d��S��0?������ۿI��TK���o;?�>�>{�s?�ľ��.�K�%��o�>RG>��'=g�je��a�̿z~�<PN?2>�>	}��#>*=�>�%?|��>�t�>�?}��'�2�����>�/?�� ?���K���̛��{9�=Vw�?I�	@�}A?X�(����ĥU=���>�	?�?>^1�<�����-�>#5�?��?M=i�W���
��ie?�u<��F�֜ݻ-�=�e�=�b=����J>�J�>��ܝA�p�ܽY�4>�Å>R�!�p��ny^����<�c]>�yս���5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=�� �J{������x�U�=����p˳���T��K���Ԯ/��M<!d�=�R5>�؂>�Њ>Y �=��">@^?v[l?ٚ>���=����h����61	=�؁��#5��%w�X!�/8��Q��_Cɾ�
����l��d�ɾp}4���=s�d�閒�@�+��+V�0V�_T0?�.>�v����I���9� F���0����=TX���ξ�v;��%n�&{�?�	7?�\��bC\����X���Z�-�A?Q�������	���F�=��ؽ�P�<�t8>����~	
��z6�3+G��2?;�?W������7>L���ˉ�$�%?)�	?��9�I�>��?G�s��0�!�?>~C1><�>xú>@�Q>a:��l�ʽ�7?  Q?����j��K�>³ξ����ɟ<���=�w?�!�,<�[C>#�<r-�����[^�c�T� W?p�h>���T!��⏾�ᏽ�L�ò{?s�?��>P.j?I/??��M���S�'��Z>�9?�Ru?�� >��輶u��n�����3?u�b?�%�=5��������/�Q%�U?�\?��?���=x(z�x����uA?ѕt?�]�4���q{ ���+��}�>~k�>��$?��6�+�3>
8?e�<Pz��a����2�0Տ?eP�?;� @]��=1*��Y>� �>�?����0����cEپW�>dt9?����=�p�9�9�>�Yb?[;p?O=�>��	���3��:>}�����?�~w?N�����=����Nw�h����="�<6ϼ��I������?��iƾD��G֌�Ϸ�����>�5@J�s�?B�[�2�׿��пj���a������I?P�>:]̽�9��ivF�d���CaG�X}T�ߺJ�=O�>�>�G��K򑾞�{�l;�����>���Z�>�SS�7.������w-2<Q>���>r�>2����н�䵙?�����#ο����͖�ЉX?�[�?My�?#c?=�7<)v��O{����
G?�Ss?�Z?9#� *]��8�)�j?�x���V`�^�4��$E��UU>b3? q�>{�-�G�z=z>d��>�6>�-/���ĿYʶ�"���
 �?���?=_�8��>�x�?u+?����5���>����*�<˸
LA?{^2>���r�!��6=�������
?@�0?��C�X�_?�a�A�p�z�-��ƽ�ۡ>��0�'f\�:O�����Xe����@y����?E^�?\�?ص�� #�c6%?�>F����8Ǿ��<Ȁ�>�(�>z*N>H_�Z�u>����:�3i	>���?�~�?Kj?���������U>�}?��>2�?���=*U�>�=������-�ܒ#>�o�=[�?��?��M?��>mc�=�X9�</�QYF��8R�D���C�!�>p�a?LwL?��b>j︽�2�� ���̽�1�|C鼋H@�,�c�߽rv5>?\>>G�>��D�l�ҾH�-?��1�o2˿S���ƀ>B|]?��E>бI?�=�X���ш��F^`?�̳>���Hܥ���x@+�$d�?P*�?7��>������=�=�ގ>�{�=��ͼbżߠ׾N�=�+?��~��=��%�Q>�a�?���?:g�?��\��
?Q���&��@Oy�js��"?��(�=��9?s��0}>�_�>�5�=��v�J����r�Dض>�ׯ?V#�?��>� h?Q#s���8�ZOO<u^�>,�]?Dq?u"=$G徚�H>;?�	�CC��w� ��BZ?z@	@pS@'\?����
ؿ�Π������Co����΁�<�>�ý-�u�c��>��=G��t`	>�g�>��>N �>��)>=�=2�=�I~�5� ��/���w��"H�����Ҿ�>�3��ï��P��̾\侬��-ߚ�.�6������~�L����5�=|�R?C}P?^�q?$��>����>u���#:U=`|����=O>��3?H|N?�r/?�Ŋ=�����d�����e��6��H��>7�L>�
�>r��>:�>���;�J>�D>\�>?�>�C>=�;��	=K�W>C-�>�9�>�>��>>G >¶�޴��Ej���t��轸�?�����I�Ε�����z���K�=&�,?T��=�w���>пU���K?L?NE��ѫ��--�v>X1?�eX?ux>/���)q���>M��o}n��;>"��?�}��+��}U>��?�$g>�u>5]3��!8�ƁP��&���-{>Է5?����c�9���u�A�H���ݾ��K>�X�>-�F��r��떿�~�hi��`|=�V:?��?uֱ�Q|��`�u��O��4�Q>{�[>�=�-�=�$L>Йc���ƽB�H���.=�y�=L�^>j�?�7�=zM�=�Gc>�l��y���O>��{>֫>��%?{.
?����'��fþ�V�X�><�?v�=-�>�,����= �>R�g>��d�.Љ����Np�����=g�"�I�����ּ�>������>�J3=G���V���P=�~?�x�������s���oD?�0?ܐ=�E<ك"�M ��%N����?x�@�j�?L�	���V���?�?�?������=�t�>eի>�ξ�L���?��Ž�΢��	��*#��R�?��?��/�	ȋ��l��'>�[%?��Ӿp��>1��{w�����Hu��,=�K�>�cH?����T��>�ޤ
?�4?���񄤿Xɿ��v��
�>K��?Dє?	�m��˚�O�?�1��>Ѕ�?1Y?�j>Zܾ��Z��7�>�@?��Q?)ֶ>�	�V�&�N�?#�?u�?��L>oP�?�Bo?�?�>�n��s,����������=O<��>�v�=�nþ��F�;Q�� J��(�k�u��+pc>��=>�>|��!f��j�=�u~����_�CU�>I�l>�=>O�>��>��>[��>[�=��p�f�s�������K?���?���9)n���<���=��^�*!?�J4?�sZ��ϾeԨ>��\?��?�[?J_�>����=���濿�|��V�<��K>1.�>�H�> ��9LK>��Ծ�9D�un�>�ŗ>鮤��Dھ�4��Y"���?�>�a!?$��>���=�s ?^�?u�(>+��>N��񋿎VQ�|M�>�f�>�^?�)r?W�?k��7f��R�������j�4Î==k]?�"?'��=
����Xo�E춽����w�f �?��o?D߽Z�:?{��?��C?�z?t&�>�vt��"z�����w>��!?�	��*@���#���7t?4i?��>����Խ���?��	���
?�?Y?�i$?%N���a��+��\{�<�Ờ�v��O<�J軒g >�>ٟ���A�=�D>�=�Ov�J:���<së=���>�$�=�0�u�t��.?����l�����<w��ȕP��K>���>���k8R?!Ύ<�[h��ɮ��9��D���#?j�? ա?G56���]��N<?�_n?�?�(�>{խ��O־Q���4��t,�-���<��>��=�&&�����]G�������J�0ox=&?���>5�?-O)?;��>V'�>l����9��8%���F� p�1����Ѿ:�&��(�C�þP{�<F~Z>?Ͻ�IG�y)�>��;��>l��>M��=�U>t�p>R�T>�1}>���A�=dQ�>�R�>��k>�8�>���>!��5	N?X�����$��Bʾ��z��H?��h?���>�b��p)�����sF?�?�S�?wTN>�!p�8|0���?O9?�Qx��; ?!�=A�D�,�<�k���:� �g��`Ƚ8A}>�彐�=��H���f�;z�>��?��s�¾�ʚ��`�����=�x�?*%?n�(�}	>�}wo�SOa���E�[�f:au�����88!���p��o�����d?��F5'�O��<�N%?�i�?�l��v���\���o�B�@��W�>�o�>��>4�>n0>w_ �-���UH���4���u���>�n}?P9>�j?Z�T?�B?�3?m�>�f�>eԾ��>+���5��>���>��;?��@?M�-?$�$?�M?i@�>� ٽw|�ξ¾,��>51S>�?p�>z�?�2ս��z!y�=��=�=ZB$>,��9��]=�ꆽ]���1���ڈ>�y?����*�]�˾0ә>�}:?�. ?�I�>����Z���b���U�>�?�>�����ir���pu�>V��?���b�<o	>�S�=gߎ�¶��l�=Dj7�N��<x����n��OK�X�=t�=�<�����"���w\��d"=��>��?���>��>�o��� ���k�=�_Y>�3S>6�>4Yپ������q�g��y>	�?�l�?fg=���=ʅ�=@T���@�����m罾f��<��?~@#?�<T?2��?X�=?~:#?��>�%�l<���F���D��G�?�!,?-��>�����ʾ�𨿋�3���?�Y?�:a�^���<)���¾Uս�>C[/��.~���lD��A��W���z��R��?�?A���6�By�}����Y��ȔC?^�>KT�>��>��)��g��%��1;>ی�>m
R?j-�>p�>�:?��?�4`�||��2{���CI���>�S�>��X?��?i�?;��?DE\?���A-�^a�Ѥ[����o/<�/��E�=��s>�p�>< �>V�!>�#o=�2i=����Ji�87�=�)�=���>��>��>0BQ>;Ƚ��H?��>僗����=ξQﰾ�����G�?)ߋ??�)?7W>~���a��r�P<M>�|�?9��?��?�"�7|�=������ۢ�3��>f{�>�f)>�>���=H�u=���>|R�>��z��w���)���1�+0?�?TU>�ǿ^q���{�>���<��<�S���MX�f���3q�Ɋ�=�2��AZ�����fB��獾G�s�H���٫����>��=���=6��=���<=� �	K<c�=r��<o:���n�2��<qj'��&�;@Z`�I���>e<.�3=Xr¼'ƾM,}?,�;?�'?�yI?H��>�>V�<;D�>蟎�s�?�g>M0����ξ�RN������ ��Q�ʾ��ϾK�\�ԍ��� ,>��g��f>�G>r�>�}�<7	>��=��=���'=�/�=3K�=�>�/�=��->�>�6w?H���ز���4Q�G[�M�:?8�>	~�=ǀƾM@?��>>�2��җ���b�s-?b��?U�?��?�ri��d�>���㎽q�=P����>2>6��=��2����>��J>����J��0���U4�?��@L�??�ዿˢϿ�b/>��6>a~>1R�-10�uT��]\�dZ��!?	�:��;�i�>���=�H߾��ɾ7_=R�6>]!Q=����Z��ɔ=�!��5�I=�k=m��> hA>�ǹ=���;�=yO=$�=*lJ>fH4�|�3��o��QK=# �=m|f>��$>"��>��?B4?��a?�f�>E�^�T�¾Ǿ�ǋ>Pz�=�ϲ>ShY=��C>���>L77?�E?�P?���>�w~=�{�>�T�>C)��lm�n��Z������<Qć?N�?!��>�Y�<���̡=����
?��-?*?�
�>��ҳƿ�I��h߾)-���֡>ڽ��D)��c�?_=i��3��>.c�>�J?j3)?���=T������ū>I\b>-Av�� ���O�=�(�=+���P=
�<�Yj���h<�8>��P>4�=n���r���T=�l�����<��R>a��>q�=���>�5!=e]V��N>�s��v�>��`;e�Ǿ	�;�%�k�k�U���B��Ţ�W��=.�>�F����vz7?D��=�"Y>�B�?*j�?�T�>��ͽ��.��2��Ȳ��,�;Ġ�>��>4o��5�fTO�I�9�������>?ٍ>���>�p>�*���=���Q=�(��43���>t���HDC�^��yq�P���[����g�����.&D?�����$�= �|?$%K?:�?v��>d����پ(�/>u��G=r��u�r��	��v?6~$?�W�>q�得�D�[����y�>r����E�Hӆ�����  �E�Z����>���>��F�;�p0��8���H7)��1�Q��>AyG?]k�?����J�E^Z��|&�DF\�Ѻ?�e�?�8�>�b�>�4?�w=������R���D�G�q?"�?�H�?�D�<f��<��>y'?ƶ�>��?R��?�1�?	���V�>gkĽ���=��Ͻ�Rm>�m�>��>`r�=�y?F�?\?5�*���쾮�۾����ýx𽪪�=�!�>�>�>2��<�k/=A�n>��=?缴�m>�|�>��e=F��=jY�>�}���6���~!?���;"�>R�0?�w�>�m>V#��g5�����󕏽˷i���k�s⤾L>�b��7I>:n�v�>�6ͿÜ�? �;J8�<��>���,������>�s.>=�Q�N�>*=>�'c>��0>��>�4�=��>��z=������>�E>�i}6��gQ��>�a����>��j�p�=���ȗ���Y���]����e�8L����N�-OX����?�g��%r�vJ�����?���>ST"?:�g�c����Q>�?&8W>NHӾ�
��\����� ���?�'�?,v>2�>2~`?"Q?'�w׽�XO�dz�Y,�5�[���i�r���XM���������V>?F�n?��A?=oM>ׇt?U����i�R>h�,���$�+ �?�>�������꼾P-��������>j�e?_z�?��?����� ��ۑ>M[Q?��>��u?��?�<L?�6��#?�Z�=+W?g&?��9?]"?��?Q�>C�>�<�-��a�$����[<���Г�u�p��5=4��t��=�R�=�:�<�F ������ϼEt������"�&=��=	pn<�Gj>Vvb?L&?��=��=?G�h�- ��H>?t�����c��1ֽ鷧�Hv�%�7>(!w?��?/�*?!t�>@�7���e��d�=��>�>>��L>-0w><���rN�����<��N>���=a��%*6��iվ}O��?Q�̂�=�� ?fx�>S��k�>_�����=������i�F���A9-���"��:B����>��E???���%E���4�w�X��n:?��?A?��r?C�k>����Z��T�(���=�ė���6�x���dﱿGB4�ƭֽ~Z>Qם�UI�a��=��������t�]�p�B��ͅ���侮��=�Բ�+z���jw��(�>�@>L�����
����������L7?���=�˾rbO�@O���q>�	�>*�5>�⨽�{���jO�|�����=�p�>�Վ>�{V;?�׾	�F������>�aJ?\�]?(�?�z�U�j�9�<��� ��N�����,�?�Х>yF?�I>Z��=u}����(j�edH�8��>(��>ί���<�>��1��?$����>��?~>��?(�]?*d?�\V?��0?�?���>�������n&?T�?�)�=�ν�(V���8�m�E�?��>�)?*�?��^�>�X?oy?��&?�yP?�?A�>1B ��?�z	�>��>��W�:���c_>�(K?�>cZW?��?4`<>67��֥�d䩽vO�=@>��2?Y!?_s?�8�>'y?ơ�����=���>x�`?��v?r�J?�:�=W�)?LY�>���>���=X��>ɗ>�$?(�i?i[?��`?Z	?D�1<F&�����Fc�=�;�0r�;�c�=���=g.������-м�Y	<Q=,�-=20=}4���r�;W��=�r��o#�>#n>L@��֪4>�Mƾ����#;>8�����r<y���F�6#~=��o>u��>��>|Z.���6=���>kC�>+o��u?�;�>�?�Ǽ�^�3�ɾ��;�#��>$@?u��=��m�K��5zt���<�5i?8e?�7A�����;4_?�@>?t2��(���*���+
���J?,T?+ *��E�>i�? �[?��?�P��Qv����9�i���o����=�>�� � c��>	�2?~)�>��=��M=�߾�l���ˬ�o�	?��|?|�?P�}?�?>6>����g��������]?g��>�᣾�_!?�{�<DϾ4��A��Z��w��������Ԓ��2���J����ͽ�i�=m�?�r?�fo?#�]?� ��tb��e\�����W�����$�)�F�KE�[�B�%[o��b��b�t��e9=H2B�y�C��̹?�I?�_�L0�>�l��N�P�Ⱦ_�>�վ�\��vP�|k�}Nb;{�<�瀾A�3��g���%?��>�7>�Q?�R�F�*��u2���<�sO�{��>W�>��D>Q��>�͝={�e�paC�Pp���%���+=��u>�c?K?��n?�"���0��i��M�!��3�}g��L�B>��
>om�>�+W�-�� &��A>�~s����&���K�	�lz�=��2?��>�y�>�+�?=9?�	�E���pw�"�0��K�<iȹ>�Ci?	�>Y��>Ҭѽ�� ����>p�l?M��>��>����V!�x�{�8�ʽ&'�>�>���>��o>��,�3 \�?i��ā��
9����=��h?e���M�`��օ>�R?���:�#H<"}�>��v���!�����'�L�>]t?OW�=`�;>�zž��y�{��4�� 7*?%�	?�s��|3(�)��>�� ?��>B��>�9�?���>|Kľ�|6Uu?3�X?JJ?f�B?O��>�L=D��|�Ž�4#���(=1�>&�[><+m=�O�=���|�^�����>=Ͼ�=�W��W���(�o<w{�� j<�
'=+f+>O�޿y%H��������B�ݾ��Ҿ��	�B[���;C�K����������W��~���>J�o�n?6�l���>Zľ'� @��?�[��-ɤ�O���6u�(>1�� �>44�5��<ag��)?��u���^H�JJ�#��|F�Y4Z�M�-��0?O�Կ$����'���=?@�2?�Uf?H�ľ���=>L��G>lE?°*����<M��"��٧�:�f?5=�>b�����=5T?F��>��>���>���o=�78X�/W�>6�?��5?_����ḿ}����r>���?�f@�8@?B|0���پe�=y0�>#�>�=�cϽ���Ǘ�>?ͬ�?~?�S/>��L��˽�T?����6��F��~�=���<u�Q�&����0>*-V>�p�1�a�),�x2�=j�g>�&�+
�C-��!)�:�m>�F���)�2Մ?{\�Ef�"�/��T���T>�T?�*�>Q<�=��,?G7H�=}Ͽ��\��*a?�0�?��?�(?Oڿ��ؚ>��ܾ��M?CD6?a��>�d&��t�Ѕ�=8������㾞&V���=ë�>x�>ƃ,�����O�L��)��=$7���ǿf�������=�(�<�#��w?Ͻ�����C�<蔾�r���D����=E�k>e>co>wV>��=d�]?-�f?���>�"6>����u�B_��s�:�,M�yTؽDdv�k�J�����/�������� ��+���	��յ���5�\��=�BZ��+����,�K�[��qe��(?1�*>�����fB�l�<"Ǡ�Kء�WN6<|Ԙ�z�׾S=�U�l����?�B:?�ܙ���f���+�ŭ��V��:�8P?
�F�/���LJ>P)�Zd2=H�u>��p�s��E�8�ɝ>�̚4?%�
?~���	q`�^<P>�[�VcO���"?�?��2=��>%^?J�I�A�)�W4�>�i>U��>��>��4>(��N���?�[?×�?N��\/�>G{���������<��	>��o�@j����>�߼����� M<at���� ��2V?.d>����u�������CZ���}?W�?�Ǝ>��Y?0�(?�V#������L�6�Ѿ���=BS<?2�a?վ>@ƾ;�����˹�оW?m?��|�Ac���P����B���:�j ?��>?*t�>ņ>�Dq�__����loT?2�s?
h^�Ǜ��a����˾Dta>^� ?6��>ݫ.����>�7?oϙ������"Ŀ	g5��3�?��?���?M�����]��#K>/v?�$?�60�����E.�Һ��Y�>n'$?܅�G���:3���!��>?��}?�a�>h�9�S�n�=*(��7�?�$�?��\ݵ<s0��o�7`���)=�j�=�k0�5�9��c��6���Ǿq�
��B��!)�����>(�@j}���>�=?��W���Ϳ̄�Њ˾p�`���?���>˿��(k���Df�lu�0kF��H�P끾�b�>��> ƞ��咾9F|�m�;���ȼY�>gw��F_�>�[Q�K:��*`��i�^<��>#��>��>0���󽽾H�?�q���\ο�����/��KX?Q��?R΄?��?k	<�z��my���T�F?�[r?fMX?��8��]�w�7�e@j?����d�e��F>��wK��#a>�:5?�w�>�-���<�b>��>�x�=/:�9Q��O���З���?���?����L?</�?{D)?����ʠ�WZ����'�Vp�<��L?�UK>�ʾy�3��<����=�?�7?[���(`(�P�_?��a�=�p�Y�-���ƽ�ۡ>��0��f\��Q�����Xe����@y����?9^�?V�?��� #�b6%?��>7����8Ǿ��<ɀ�>	)�>�*N>�G_���u>����:�=i	>���?�~�?Dj?���������U>�}?^�>B4�?_��=s�>.�=�b��)�u� [">��=��.��D?Z�M?#��>���=��6�_�/���E��jR�/��� C��0�>��a?��K?�b>����j�*�n��~�Ƚ$�0��"ͼ�T>�7�/�B�ܽ��3>��=>q>�B���оOs'?h+I�pտ�������Gke?���>�n?� ��;��"޽A�o?[�?Sx(�*������>lN����?0��?��>n=��g�r���!���=���<f�*��7�emN�܍q>��D?��F��C���녿�M�>pr�?Yu�?(y�?�0��A
?a���o��ڛ����&5�ƿ�=�6?�0�i?v>���>���=A&u�V�=�s���>*�?c��?̆�>7�h?HTk�b:=��N+=�p�>ӧ_?�?~E�;��zX>-?1����і�3�a? 7
@j@��_?�����׿񘚿����)g��,�>�В=.6c>�2ѽ�e=��=�F�;G�%�r>(�>Ua�>�[�>ۨJ>�5	>1'�=9��e�"�Õ��aH��&m9�����.��xl��%�Z�O�cJ����7@ľGf��l+��t�p�Һl��16�����h=×^?��A?�t?��>�~c���=�qվx|�~F��>Jư>�S#?�;?OS=?� 
>�����y���~���Ծxm���>m��=!��>��>�\>:�>��>� >�?i>%�A>U��=�
����=��>TZ�>��?��>�<J>? >#^������_y�j�~��u����?�����y=�w/��{e��&����=^�'?��=�M��'�Ͽ_է��TU?���r��gNz�"�=�G9?� x?��>����-˽�I�=G�׽Fc*�,;�=F
6�,����:�P�i>��?2�g>��s>^�3�M�7���P�=P���Ez>q�5??i����7��u�H��ݾK]N>U��>Ҩ]��C�  �����i���z=�P:?�s?���k����t�洝��5R>,\>y=�o�=�^M>%�c�2Bǽ�G�Ko-=c��=\�^>�"?F	˼~==�8�>ۘ���Ӿ$��=�>�>P�>LA?c]G?�(�=�*��a�M�F����=-ܰ>�*>+p�=ֺ���>⠽>���=�A=;��=F
���0��0>���'Ɨ��i2��v�< �4�k-���K>��4�Aм�>��~?���2䈿H�=e��[mD?�+?!�=�yF<�"�0 ��H���?6�@�l�?�	��V��?7A�?���۶�=�|�>d׫>�ξ��L�ӱ?4�ŽnȢ�U�	��(#�DS�?a�?��/�#ʋ��l��7>�^%?��Ӿh�>;�����t���=�u��P=wO�>�0I?.t��Űs��>C��}
?��?��W�����ȿ�w�$�>s��?��?�Km�7���g<��h�> ��?{�X?
ql>3~߾i�c�(s�>��@?cQ?�u�>���W$���?w�?�0�?�I>���?��s?-o�>�xw�]?/��#��L����|=-�E;n-�>1�>�����CF��ӓ��o��?�j�:����a>lA$=��>U�㽐^���ص=0���[��=�f����>�Rq>��I>�F�>�� ?�:�>}��>��=����B���Ж���K?Я�?���+n�i��<�d�=��^��"?�G4?_rZ�%�Ͼ�ڨ>�\?�?@[?W�>K���>���翿�z�����<c�K>�2�>2G�>A���JK>��Ծ0D��o�>ϗ>9裼 :ھ�+�������@�>-b!?Ԗ�>ܮ=�
'?@�>*;->Q��>E�W���6�/�u��>��?RYL?���?IZ?N_����׾�Ay��j��ɋS���_>��?�g? �<X?l�_Cl�ȅ��M����(�ܜ?��f?7�N{?yU�?��?��?�3>�V9�6�����t��O#>]�%?[=.�m�2�FK&��p��t�>uA�>�C�>Tz�<�ܽ�����6>���	�D��>`�S?��?���o�U��H���<{�)������O=U�M=V5>e�>�
ս2�=�)G>�p{=٢��}����<����=kԵ>��=em��Lg��o.?6��放���=��u�v�B��@�>i>tì��}a?���hl�x���="��.���Zf�?�ο?u��?�F����e���H?��?�?�?y���0R��4�h����z������D=q�>=�4 �de����������E4޽�O�I�J?��X>��?!"?��>j ?.�Ϫ���;;���(�:z}�� �\���ɽ%��t3�Y���A���7�q�վ�	����>%X�٥�=O�>��=f�>5m�>�
��)Q�>�E�>K>�W�=��>3x�>O�+>	���X��H?ٙ����)����Ĕ���L?��k?���>F
K��R��j����>��?* �?��,>�v��2���?O�?�w~��}�>Wh=�t������A����z7�����૶��3|>�ĽFu4���Q�k�r��-�>��>����u�ξ�����ɋ��c=�́?h�)?=*"�ˍB�\k���b�g�L��=�����ʥ�Pf�8�l��ĉ�9͂�҆���]���=��)?�2�?Hq�u"ξ�$���n���9����>���>Sˣ>Ϙ�>&�G>���#��$Q���*�Wu��;��>:�?��>�lN?�:?}O? M?ǎ�>�A�>8����>��L��N�>�8�>y7?z�'?t�4?��?X�1?ƼC>[��g���Ӿ�?#�	?��?�p�>��>�	s����(�>�:��K�|�����17=��=�uн��~��&�=��a>F�?����;5��U��:>cM'?nY�>���>�p`�͚c��������>I� ?��n>����bi��@�<��>Q��?y��!�<�>7@t=l���r9<{��=EMi�\�'=���k̽م���=c��@�����<��=�\1=],�<a��>��?æ�>	��>o���Z ����]�=gX>��T>��>�pپbY�����3�g��x>�'�?�V�?��k=�$�=���=e���~��7�-����d�<��?�l#?OT?@��?�=?܆#?�>w��yB���6��R^����?=!,?��>���ʲʾV���3�՝?�Z?�<a����t;)�"�¾;�Խa�>�[/��/~����D�Hą����F�����?���?yA���6��x�0���;[��ܓC?{"�>PZ�>��>4�)���g�=$��3;>Q��>�R?�X�>x�?5�:?<@U?���<`�^�ζ��Gć�38p=�Æ>�MT?�u�?��s?9�?���>�Y��+��2�c���ּo
��$rA����='�]>L؜>@�>]�>I�=��~�_��(�$����=r�>u�>&��>�j�>���>:3y=��J?r~>������θ���y����ҽ`l^?�ғ? �:?�(p=�,�&�N���Q��>0k�?�?�x&?����dH�=�?������,�����>��>ﺡ>��>���=~KE>E=�>��>��;�����M�d�B>��?K?�)=5�Ŀ�n���c�����՟<??��\Ga��Ø��fW�z�=�\�����%ߦ�uTR��朾b/��E��%���c��+��>.��=���=�?�=�A�<�JѼgg�<�P=�;<�=�u��I<<j�I�WN���Ŗ�=�j�
�M<�]X=f���'��@�?Xe?���>��U?5fv>���>�9�=�>�z��r��>�m�>�����}���0����M=�TT��lʾn�1�J��?ƾ�8�=p)��.�>�-4>���=�(��m�>\�=��=��=��=��=���=���=:�)<�A=��=�6w?X���
����4Q��Z罢�:?�8�>q{�=��ƾq@?��>>�2������zb��-?���?�T�?>�?8ti��d�>K���㎽�q�=4����=2>g��=w�2�V��>��J>���K��8����4�?��@��??�ዿ΢Ͽ=a/>5q>�ʁ=bP����>E���M��eG���C?	�!��ђ�_q�><�&>�Hľӕ�����=y�l=\�=2}�~bb�~�=B_}���=�3�=!��>�wO>��=���"<�=��f=Uu�=��F>5�<HYB�����_�e=k��=);�>�Z>>���>��?V�/?�Dd?��>		h��;���/?�>��=�o�>�ܑ=��A>Ŵ�>�9?��D?��L?��>��y=#_�>�!�>O�*�#�l���ݾ���0�o<3�?r�?��>��<�e<�Oe�E�?��N����?UK1?~}	?c�>���࿉�%��.�eS��̢�:m�$=$q�ޣR�����Z����~K�=�$�>��>�O�>Xw>��5>oH>;��>	:>��<���=6껆��<��̼[��=c*u���< m��!���n���7�O>μHؓ;��;�g<�^�; �<>��>��j<��?�W>�45� y">�m�1�H�~��=5�ᾍ�q��r���<��f>��A�f>0��>�g/������;?[
>��+>��?���?���>�_k���4�󷜿��˾B��D�>�`>��<�kT���z��R��:��X��>�\�>b��>d�m>^L)���;���=H��8����>`�����I��I��>m�Ɋ��Q<��2-i�6�C�Q�A?3���
��=.8~?�I?�?DW�>c/���FϾp\<>�X~�2�A=�Q�Z�i��ޠ���?z,?�>���E�d♾�5޽��>*5C�=P�\Ϗ�G��5����d��>�����t�I�1�D����׍���9���R���>˃B?e�?�e��-f���Q�a(�]��?�~o?���>�
?��?�|��q���4~���=<)�m?���?8ڷ?�Z�<��;X��s��>���>�(�?*L�?A�o?{<��o�>�U=W>Y�����=&��=J� >j�C>�?�� ?�e ?���|��x�v�辚	
�W-Y=�lr=G#�>���>,?�>e��=�%W=���=CGn>���>	�>�f>2�>�w�>nV���|�$	J?����T'�>j?�A�>�X>l都.��X���g�,Q]�넣�@����m�up&�oM>A�=��W�>A&ҿ�ģ?��?>��̾2�?���G0��M�>�X�>�%�kӖ>�=�=��>K�	?�1�>'�E>���>ӈ>����|�	>�y&��u0�0VQ��LN�¬��у>��
�����۩�|M�������/g��y���H���Ż@�?A�6�Dz��7���I��?�8�>:+?�av���CZ�=�a�>��>�辑��}���$-��?�/�?'Gh>�>��U?c�?ԭ)�7�3�j�X��t�i�>�&b�S�^�}w��ⁿ���.ƽ��^?�rx?�B?)n<�-q>ƙ�?��$�1���r�>�@-�0�9����<@+�>�d��a`��پ1�ž56��%9>��i?ʂ?
"?�[�f�!I�>�m`?d��><��?	0?�;?�޽���>�:=�%�>O��>#?��?�W!?��?�=�>��ؽ~Z�UU(�)���_�&�ؤ[<����� �I<z���`͂=P;>�o����h��d˼z�=�ț<��#�-�=kF�=3�=��$=8�x?�?��>-X?�0��D�6=ʽy� ?�$�jfJ�Udb�$���l���>�o?��?1;-?��>l���;���X>�ZE=��>*/�=��>���!<;��]���=�Q=�_�<}�B=�Ӿ�U�zԅ��a!>�1=;� ?j~i> �d�B�}>�(���rx�}IO>EeM�K���e<���=��6�re��a��>��@?��?i<�=8鸾�����da��-?��.?F�H?|�k?��Z==Ծ-�B�K W�N*#�&#�>(e����;��'���*@��n><�CG>����ܠ��_b>|���t޾]�n��J����g�M=~��V=���־�E�b�=�$
>����� ����pժ��,J?�`j=�s��YU�Si��#�>��>�ܮ>��:���v���@�۟���[�=b��>��:>U��)��>{G�j7�v;�>�NE?jU_?�h�?x���
s���B�<����[��n�Ǽ�?ux�>�g?}#B>���=�������d��G�/�>��>o��z�G�3<���2��	�$�ǔ�>�5?��>~�?��R?>�
?F�`?b*?4C?,�>���E����A&?��?��=��Խ��T�q 9��F���>��)?V�B����>M�?߽?�&?��Q?ڵ?w�>� �yC@����>HY�>��W�zb���_>h�J?��>�=Y?�ԃ?��=>0�5��颾�թ�W�=�>g�2?6#?7�?u��>#Q�>����(��=}��>l�d?���?��p?w>	K ?G�K>6�>>Բ=���>J��>� ?guL?�q?sF?"��>\��<Sڹ�0n���2������μ<�-(<�9~=`$���b��I����<���;x����w��aѼv�>��'�7�; V�>��s>���	1>��ľ�Y���@>N����P���ي�9�:���=�{�>c�?���>*�#��t�=���>SN�>���y>(?��?�?�; �b�K
۾��K��!�>�A?��=�l�K���u�u�Lg=D�m?��^?�FW������p?T$B?�h&��Q%��ܾ��I84��SQ?)�@?
򽍊.?��?~/n?X#<?�A|�D�b�.����?s�����B2����>~U�[�C��
6>J�'?M��=�cV�a+�u�žE���7ž�?8IE?*��?�k�?�= ۃ����_i�� ���gW?���>t���8?8vO;��о0����ⅾv�߾�߬��v���#���!���Y3�q���.���Er�=6?��x?Q�h?xa?U���f��b_��M}��Q�Ҍ
���B�B�HXI��qC�θn� ����뾧o����e=Dp���A��m�?�;$?��#�E��>���?�ܾO�Ӿ�6>F������J=��ƽ�L=�:=�Hj�e�!��尾M�#?�g�>@�>j�A? �U���8���2��a;��w���Z�=D�>Um�>)�>�eu�,��PYϽFn����V�(���4v>_c?+�K?��n?@���1�ǀ��;�!�'m.�^L��hC>��>�݉>D�W��z��'&�$]>���r��������M�	�7��=�2?�K�>�؜>�X�?�?e	��p��`Px���1���~<L�>��h?��>8��>*{Ͻ� �#��>O�l?��>�>Й���T!���{��ʽ+�>ԭ>���>��o>��,��$\�7j�������9���=��h?����C�`��߅>R?f܌:��H<���>�v���!�A����'�e�>�?Ϊ=��;>�ž�)�Q�{��,��S�?u:�>��t���G��ͭ>Q�?�?5��>:�b?���>��e�=��?F�i?�IN?c�+?G��>�������I�j�Y�S���<���=<:�>��)>袔=�K��V�����9�����=����5��)Z�<�=#��'�<�i�=���='�ǿ�;R�������#��
��6�������4!=7����=����(���q�c�=���������5��Mo$��b�?�6�?�\��
��tg��v��"6��Ă>�}�P;�w���C��-ھ�%����ƾ%(#�HQ=��d�C�=�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >[C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���|¤<���?0�@eA?(���[b=p#�>R
?�wA>��4�wH�s����>w��?���?��S=:X���!���d?�2<�F���ѻ���=xR�=�K=�L��OG>-��>����J>���ٽ�,7>�n�>�))�?N�;`��Ѱ<mY\>�ؽ�1��5Մ?{\��f���/��T���T>��T?+�>�9�=��,?U7H�]}Ͽ�\��*a?�0�?���?=�(?�ڿ��ؚ>��ܾ��M?kD6?���>�d&��t����=66����y���&V����=��>!�>��,�֋�g�O��H�����=����bDƿČ�{��H�9��c=�ع<V�ɽŲ�-ij=����3
��7T��7�;o�@>'K>>âF>�A>ENW>�7f?��\?<�>}+->L��M��5쿾���!���_3������1g�1��(T�����u��X,!����}���=�E�=7R�ݔ���� �U�b�x�F��.?
r$>"�ʾZ�M��,<
nʾ�Ī� ����襽w)̾}�1�Sn�x̟?��A?����,�V����C�������W?O�����笾y��=c_��E�=�>ߞ�=����3��yS�R[0?G;?Bs��@����*>@;�=H�+?�?wd<3@�>�9%?i�*���⽯�[>L�3>p�>J��>y�	>u뮾5�۽�o?(YT?�=����s�>�ǽ��{��Bc=)I>J�4����c'\>�C�<�􌾎O��܏�x��<�W?⇍>��)���!d��YY�&�<=�qx? 3?T��>�$k?#�B?ޤ�<�w����S��w=�W?�i?t>Ƽ���Ͼ:��=�5?��e?�>P>ui�!
���.�6F�*	?��n?�?AM����}� ��S��z6?��w?;pS��X���x�ܥ�>�\�>Y��>7�:��٨>SB/?�O�����8߽�3R+�o��?iv@;a�?�컒 ]���=�?4��>uN�)޶��9ν}���[bA=��>E�����j��)�c?A���1?P�y?Kz ?��g�������=�ѕ�T�?��?�����%h<���l��|�����<]��=�X�0f"����7���ƾ�
�����>��g��>�X@�o�c(�>�K8�v6⿩QϿ����Fо�Yq���?@��>��ȽԐ���j�	Lu��G��H������v�>i�>�ܔ��ޒ�q{�;������>��v!�>Y!Q��=��w�����^<�֒>1��>(�>�[�������a�?�#����Ϳ�u��� ��W?�;�?��?F�?n�}<A�s�:�z�أ�T�G?��s?(Y?}���Y[�c�D�Q�j?3Y���S`�z�4�*DE�)U>[#3?\6�>x�-��1|=�>��>^>/���Ŀ�۶�e���s��?̈�?�k�!��>%�?�o+?ag�9��.]����*��D�9=A?�2>E�����!�y)=�^֒�(�
?S{0?���*�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?K��>̓�?Ao�=��>���=S����n���>�f>TG���?�N?}��>o
�=��6��Z-�
F�{xR��2�xC���>�:c?�K?�m>���=��#< ��Yʽ�=4��m���=���3�վֽ��+>o4>6�>��7�Fʾ
�?�o�-�ؿ�i���s'��44?(��>^�?����t�����:_?Yy�>=7��+��v%���@�U��?qG�?{�?��׾�N̼�
>��>�I�>� ս��������O�7>��B?!��D����o�r�>���?��@�ծ?Ii�D/?���Ԋ��%l��>�f-w����=� >?d:�k�>p��>��B���t�����|�o����>2�?/��?uf�>��m?�j��p5�d�����>��b?LY�>""�<���jSM>���>$��닿C�jX^?o@s�@��[?��:Mؿ%���tE¾?��mO>%��=�Ot>����z��=\y�=0�'=��z<�	A>���>F�f>g�>��(>���=[�=�~��� ��0���"���.6�+�	����ֻs��J�4V��5޾���Jh���~1��@��X��2�(���6��-���=��j?�lJ?��?���>���<�>�_���Z>pO��${c>��>��A?	{4?�$?ѯ�=�ž$
j��]w�3.Ѿ7t�g{#?��g># ?���>�?��5;�Om><�f=�V>f�=��3�1��R�7�]=�1�>͘?\	�>�C<>��>Aϴ��1��h�h�aw��̽$�?J���@�J��1��H9������i�=[b.?|>���?пl����2H?����^)�S�+�X�>��0?�cW?��>I��%�T��9>^����j�E_> + ��~l���)�V%Q>Ll?g�f>�3u>Ȋ3�b8���P��w��L|>U66?��j&9���u�:�H��tݾ�%M>���>j�D��e�%�������i��y{=t:?2�?����Ѱ��u�r@��9UR>�9\>�=���=0nM>�Zc���ƽ�G��.=X��=�^>��?~#*>Dۍ=({�>fK��6�Q�ղ�>��F>r+>n�@?2%?�3��ɕ���� V*���v>���>\7�>ʧ>M�H�)�=P��>Y]>�c뼪�}�~�-*=�kER>�Cw���_���n���u=���(��=��=�~��b_;��{=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾRh�>xx��Z�������u���#=Q��>�8H?�V����O�e>��v
?�?�^�੤���ȿ4|v����>X�?���?f�m��A���@����>:��?�gY?ooi>�g۾=`Z����>һ@?�R?�>�9���'���?�޶?կ�?II>팑?S�s?r�>�x�(P/��1��̖��7�~=,>R;�V�>�?>����aF�2ؓ��k���j������a>�$=��>3L�U5���A�=3"��sH���rf�q��>4q>�I>�_�>g� ?�i�>���>om=L|���倾8�����J?���?�#�ux*��--��9����}p�>l�-?�������e
?䇀?�l?�j�?�#�>�,;��n��!�ɿ��ݾN>�=fͻ>p3?���>�4>�\�>�'�>�=��4�>k'�>R�3�q�>Ծ-�-<��>yj?>r�>�A�=\5?a�?���<͜�>:X"�����K$�t��>���>|A�>���?��?G����?�����b��Κc��T>�p�?�� ?ԣ=���֕����}�����1��R�?!L�?��>Cބ?�ܼ?0�n?��E?�;>�6�=Ѝ���ɾHv�>G� ?��Z�@��E'�����?!?i��>sٓ��aǽ���pl��Y����?�;\?�%?�]�u�`��7��D5�<�YJ��r��$;w��h>�g>}̓�>��=`P>0@�=F�j�G^5�\�F<8B�=��>]��=��4�g0���-?�Y=Ţ��,N�H�]��;�(�M=�6�>���A
:?�κ��Ձ��[���E��	�ݽ��?p��?p#�?�!>�_#u�$�<?�u�?�+?���>A�I�5����*���U�|轖���W��n�O>,��� ���
��,Ҫ��Є����B����N?>��>g?�:�>dB�>�u�>�ڥ�v�Q�����)��p���0�3L �%�2���H�=�x�sּ�<v�+7��-aR�خg>WQǽb�>���>d�w>�g>��>+/�*2�>��>p%Z>f��>0�&��G�==��<�½�\��#R?����t'��u���tC?�jd?��>�$��<��]�0O?�Α?�K�?�=p>S,j���*�?^��>[�~��g
?�4=l/0�#$�<^ֹ�/3��o�Dj󼛡�>��˽��8�[M��[`�R/	?�k?�T��-7;��ѽ�C���G{=#	{?��&?�b1�p�S�ue�Y�V��N��Eۼ�a��h���� ��5r�Ċ�2`������+���i=?�.?c=�?#h�s-ԾPl��7n��D��j>�f�>��w>���>@I1>+�()0��4a���K�^���>9Yw?7X�>��L?�W=?v�S?�8H?�x�>o��>�=��@��>д;��>^��>��:?��+?Y+?j8?DY$?�K> �����؉Ͼ�?�W?n�?��?��?i����ȶ�7���7��4u��`����=>��:-��@�>�``�=uYg>�F?v����8��+���k>Q�7?��>���>�)���Ԁ�R��<f �>�
?�e�>���;`r��D��<�>x��?ު�0�=z�)>h��=�������=��¼���=܃����<�� <�g�=<%�=��}�hF�No�:;��<N!?4?h�T>�\�>�,���棾ނ,������:AA�8���������٫��o�>�B�?��?���"�=\��=h�y� ����������>ӡ�>�o�>�1E?7|~?��?��B?&W>��Ծ�᝿Y��I/���k-?� ,?b��>���p�ʾ�𨿦�3���?1W?]6a����u5)���¾�Խ��>�Q/�)~����RD�b]������n�����?5��?I�@�~�6��h�6���TS��דC?�&�>�L�>B�>��)�g�g��#��8;>ې�>�R?�!�>/�O?<{?¥[?iT>��8��/��6ә�H�2��!>�@?±�?��?�y?qs�>��>�)���P�����������JW=�Z>ؐ�>�)�>��>���=J�ǽ�W����>��_�= �b>��>B��>i�>��w>�N�<�	T?{w�>Ӏ��+v�����{;��.��fu?-mV?ϑ?bމ�V{<�OQ��/��ޣ>�ɩ?"h�?R+8?|�&�P>�3�9�oK��N��y�>>�>�f>���<�ў�O;�;��>���>s��ox���^<
>W'?
�,?��{�ſ�s�6o������<�d��.kN�]���IQ��v�=;���S� �ʚ��6�`�����⑾Tʴ�%-��u�(?��r=SD�=��=M�G��Լ��<#�e=Ciw<�_=bFx�Ԧ�<Q氼��Ѽ�3H�c���'�m�/=�콻�q¾�3�?�[V? ;?-�>?�q�>/1\>������>�½��?,�>ͤ�<a���2P�	ĳ�##��#�ؾң��>�t�������4>���"�h>�>� >T���O�=���<��4=�y<|X�=��%>�T�=C�=�� >n�B>�d]>�6w?H���	����4Q�4\�n�:?�8�>D|�=��ƾi@?�>>�2�������b��-?{��?�T�?J�?$ti��d�>1���⎽qp�=L��� >2>l��=��2���>J�J>����J��ف��q4�?��@��??�ዿ��Ͽ�`/>PO>��>[�S�,�2����R�w�(�d�*�#?#:�q�����y>�b=���9b˾u:@=�>[>�I�=���|�U�m��=��h���m=�=��>OK>���=,3���3�=���<��=4\>"���a�J������=���=�f>�T>�s�>O�?�X0?�7d?�3�>i�m���ξ�5���j�>�u�=iO�>&�=��B>d��>�7?]�D?�K?a�>Q�=R�>]�>��,�y�m�=h�5৾4Ů<5��?���?��>^6T<i�A�w���;>�bĽg?�[1?�c?2��>�R	�W��|����E�r�X>ޘ&>�B@>�-վ�1o<��=34N��2	�pu2>K��>*!?�ޑ>@�>l, >njͺw��>Հ>��=ThK>6w�$j?=:�=�ap=�8�;�f=a�j���=��,��{C���N���^�F:�<
��<��8>���>�P5>ʫ?�G��7t.����=�[���0j�c���2��:R�G^��{���$������>�\�>�����·�:?oyW>�ui>Q5�?�x?���>\䆾��ܕ��tB�æN��8>Ȣ�>d�?���t�Ŭl�P��5��5��>n�>7 �>�l>],��?��x=�⾻j5�q��>y������.��3q��?�������i��PĺҠD?�C��q��=�~?Q�I?��?���>f���v�ؾ�?0>ZI��.=q��.q�j���E�?k'?���>C�ѻD�Di��
����=g/_���{�ș��#�=�<����?C�>�񦾱~��4�,�<'�������%-���]���>xsN?&��?�0���o��%�	�����Mcr>�|u?;��>���>X�>�����^�9Q�׋�� z?���?�?D>L��<��>�>Y��>Ǭ�?�X{?��r?h�G��G?��=��V>k�<��4>P��>*�=�<�=��>�Ų>�?[x�����	�'	������	(Q�a��=�>�
>eܖ>~>K.�<��=���>u��>�ez>�N�>�/�>�LA>?����� �vD?��<��>,g'?kq>�]z>�1����="����T�{Ꝿvag�Ho��p�<�zf�k�={!�~h?{�ɿN=?Qy�>���G ?��¾M���}��=Ga�ȥ��u?:=r>z>�Ͼ>�D�>�Ӭ=<9�>��S>U;Ӿ��>����R!��<C��R��Ѿ	8z>m���O�%��������?I����tZ�tj��,��s@=�^��<%I�?�t��ľk�X�)��M���r?��>S6?�����̉���>
��>�~�>�J��?���꺍��1���?���?>��>$%W>f�B?�B?+����@W<�]c��Hc�S~_��B���n�\w�0���k{-���ӽ��a?L�?[5k?���>?��?2�h��)�#]q>����Q�O�l���>�������ɾP&��VA��߽�{?W=�?�3@?��N�2��)�>mdo?�\�>��?��?��e?�4���4?*�}>� ?�?>/@?NrF?e��>e�=ړ�=�Z�;n�>H}���Ӿpo>���� bX=f�<�ޑ�"�<��)�SQ+>��p�~Cڽ����JN�5}�<PS�=9`j=�=��=�`�>q#Y?�x�>�ň>�05?3��=�Q���@� ?�[F�z�������?�������Ō=�p?�j�?y
c?��>>@�>�	N8�J�>F�>m��=]_N>��>��˽y�;�Wj�=N�
>�5�=��=Co��ϊ�w�	��g���̤<�F)>B��>��~>`썽pc+>m����y�ka>K�S��举R�;�F�ܶ0�Rq��N�>��K?ξ?/��=@r꾮ʜ�Dcf�)?#�=?�BM?�?��=�Pؾ�9���I�/���k�>�}�<|�	��t���k���:�t�[;O�u>j���l����d>H��N�޾n�ϿH��$���A=�����X=����^پ���� �=:	>�迾�K!�����@����G?��u=�C����N������>�|�>ĭ>~2��Nd�=?�!��z|�=�,�>��:>{�����_JG����=�>PQE?UW_?�j�?X"��*s���B�U���|c���ȼ��?�w�>�g?bB>���=.�������d��G�j�>?��>E����G��;��c0���$�*��>U9?��>��?��R?��
?[�`?�*?,E?'�>���m��� B&?6��?��=��Խ�T�� 9�JF����>|�)?!�B�ܹ�>P�?�?��&?�Q?�?��>� ��C@��>�Y�>��W��b��=�_>��J?ؚ�>s=Y?�ԃ?w�=>]�5��颾�֩��U�=�>��2?6#?O�?���>���>᭡���=��>�c?�0�?r�o?ā�=��?:2>���>[��=&��>���>x?XO?0�s?��J?��>���<�7���:��IKs���O���;_H<��y=���/1t�L����<�׳;�o��TK�����7�D���ë�;��>�s>pv����5>R�Ǿk���=>+ü8񚾂݊�il9�F�=��|>&� ?g��>�?)�nD�=.�>�=�>�����(?��?��?�W:_�c�Y�۾��H���>�@?ĳ�=�n�����u� �\=�n?��^?�FO�.�����j?�XK?�����#��ɾ�s.˾�	�Ra?�!:?�y|���>_P�?��?�9?�\þ�}��򦿤I\������<{h�>2���������>��A?z|��JҔ����<I����|�s�l���?��?��?0�u?�F>�o�k�i�;��C�??��>%�о�w?ޛ��� ݾ[V��YF�kCžZH��+���ͨ��)��-x��0㋾꣭���=��.?D�z??6N?��a?�0�v�_��g�B�~��W6����q��dTW���_�_�H�K�h�Gk ��'��X���i�=>�u�B�E�;��?�2&?�.���>vL����XоP�J>�o��{R�h��=�驽�YR=�H=#�g�.8�����kJ"?���>�~�>�9?�R�<�3���3�K'=�*? �g/>EF�>�֎>µ�>v:�� �5��x��@�\���׽�.v>�yc?��K?��n?t��(1�D����!��/��Z����B>�[>ο�>:�W����[9&�Y\>�3�r�g��~���	�o�~=�2?R%�>���>"O�??Vx	�Ag���[x��1�-��<�1�>Oi?�:�>��>�н�� �C��>n�l?T��>���>�t���"!�f�{���˽R��>O�>dj�>�o>��,��.\��g��u��%�8��E�=Urh?�����z`��ǅ>�R?�6�:�JO<��>Fy�f�!�j��b�'��>n�?ئ�=&;;>�užy�а{�{����O)?xK?蒾��*�+5~>�$"?���>.�>K1�?K+�>:qþ$�D�ɱ?�^?1BJ?FTA?'J�>��=�����<Ƚ}�&���,=���>�Z>em=c~�=���vs\�w���D=eu�=֡μ�O��@�<k���h�J<��<��3>�Nֿ��Q��B�	��)����cmr��+ҽJ;��l���-Z��v����f�������u��`e�R㑾��V��?� �?�6��b�W�����I��s��p�>;SM�A{�[~��W�G�����K�쾼����Z&��L���_��TT�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@wA?(�Z)�X�S=��>�
?��;>�R5�2�\������>���?V,�?��;=\�W����e?�B<(G����+_�=}�=��=:��&CJ>5œ>���&B��ݽYQ4>�p�>���x��k�_�Rٴ<�\>�e׽���P��?�X��<h�PO�L���x�9fp-?Y\�>VN���>��U��ҿ��i���t?Y@�E�?�q*?K����	�>�־�4?�_M?���>"-վYDS�\I¼�g��� =���Xxx��y�=���>���=c~h�0��?<��Q����z�=1.����˿s�(����t\���=~�<�R߽���]�>-����~�|*w�V&�=M�>�G>e�l>9�*>d�?>r?�4`?��>%�0>ƽ��c�b�N�̾$孼�s��R,�雈���s�n���*N�W۾���Z����%��� =��=�6R�g���Z� �Y�b��F���.?xv$>$�ʾ��M���-<�pʾ����ۄ��ߥ�]-̾Η1��!n�W͟?��A?�����V�8��AW�Q���'�W?�P�ϻ�Yꬾ~��=ಱ� �=Y%�>���=M��� 3�~S�$y0?�I?�p��hH��7*>t= ��y=E�+?�7?��E<}̪>-/%?�y+��:���Z>a�3>��>/
�>�w>���B�ڽQk?xT?���������>䉾��{���`=�>:�5�����,\>���<���?p[�7���ӿ<�M`?��F>mT5���P����'��@�>Gf�?��?�|�>Kf�?(6B?��=�g�M�{��)&�E:��{�<?�Zz?	`>tu�u$ھ5s���S.?�MJ?���=T�}�gI��^9�u���?6�?g7'?H��<©t�.���+_!��6?�v?��\�I����y	�Pgl�'�>�{�>"�>o�8�%�>�9?v.6�	��0꾿�H/�O,�?9@���?�Zi<(�T�=^�>)f�>8�:��r����<��jr=��>O'��D~o�X#�$3��v@?�D�?c7 ?� ������=�ٕ��Z�?}�?����Eg<O���l��n��z�<�Ϋ=�F"������7���ƾ��
�����࿼ݥ�>DZ@�U轀*�>�C8�Z6�TϿ(���[о�Sq���?-��>��Ƚ����@�j��Pu�W�G�&�H�������>�g> 𗽳��8 |��;�s���%P�>�I
�K�>��S�>ֶ������3<r˒>���>�	�> ��Bc�����??�����Ϳ������X?%V�?*1�?�?ۑ%<��u�zz�hT;�bdG?qt?XZ?g ��2^�m�;�%�j?�_��xU`���4�uHE��U>�"3?�B�>S�-�f�|=�>���>g>�#/�y�Ŀ�ٶ�@���Y��?��?�o���>r��?ts+?�i�8���[����*��+��<A?�2>���G�!�B0=�SҒ�¼
?U~0?{�f.���_?� a��q�9 1�nz߽@�>qF-�e�Z���$�6%��nd�@���[������?�	 @RR�?���P!���$?ڏ�>ߥ���@þ_N =�l�>Ҵ>o�A>mar��
s>���k�=����=�??z�?��?�3������K9>B�|?��>כ�?Њ4���*?�<>N�Ҿmk��eJ:>	T>�:0
?S~H?aM?`E�>C�<���8�%yY�a�\�~��:J�A;�>��v?$"n?��>,5k���)>����F� GY�$7=�+�)k����~�M>�rF>A`H>�|��_e���?Mp�8�ؿ�i��)p'��54?-��>�?����t�����;_?Mz�>�6��+���%���B�`��?�G�??�?��׾�R̼�><�>�I�><�Խ����]�����7>0�B?Y��D��u�o�y�>���?
�@�ծ?ji�9�?��1���Dg����mw��R�=H4?8�)Y�>�O�>�IE�6�}��f���3g��R�>�a�?�W�?���>f=l? �c�K�7��9����>ɭ\?�$?��}=+����%>4��>���8g���2���h?��
@�t
@�wZ?Ӑ����Ϳ����sU��D���D>dQ>�O�>i[#��5>�q=#�=in�=P>P^�>��>�2V>�9>���=I�q>kz�m ��Ǜ�zc���8M�������c���߾�~4���	�̾ͳ��`��ܗP�t���0�J�:������~<Z,s?fP?h�?c�?+-�(�>�ɾ��>��ͽ�� >&�>�83?T?ܾ?��9�)Ⱦ�o�VWn�����]���?Eɹ=��>��>1Q�>n�*;�OL>N>Vc�>ﭕ>�5���x��'B�9��>]³>�y�>�@�>�C<>��>Fϴ��1��k�h��
w�q̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��v�T�4:>9����j�5`>�+ �~l���)��%Q>wl?��M>�́><$�kx5�#�O�Š����>�/?⺾ms-��F|���M��ھ�:>�=�>�f_��d ��떿5Ã���q��un=̾4?�7?��ƽ�k���.X�%���C�Y>L!_>|D=�<�=��^>g2�1Z���F�k�
=P��=l�E>yX?��+>���=�ڣ>�`���/P��y�>jB>	,>�@?o$%?s������&���L�-��w>V�>��>O>�ZJ�i�=�h�>��a>y?�=���ϫ���?��cW>%~�1~_�L�u���x=l�����=�=�� ��=�R�%=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾSh�>|x��Z�������u�<�#=S��>�8H?�V����O�X>��v
?�?�^�ᩤ���ȿ6|v����>X�?���?e�m��A���@����>:��?�gY?loi>�g۾A`Z����>һ@?�R?�>�9���'���?�޶?կ�?yI>p��?o�s?\k�>k-x�zY/��6�����~\=J`Z;�c�>�V>�����gF��ד�Dh��z�j����v�a>��$=^�>JE�n3���:�=X틽G��l�f�,��>�+q>��I>rV�>�� ?�b�>t��>�w=�l��‾]���4�I?���?L��|�W�:�<T��<P��#� ?!�9?��=o$��#F�>�(i?���?^O?��V>n���-�����K���&�=I>>��?���>����W�1>4FԾ�$z��O>p�>h����:�ޫC����=�X�>XV?8@�>H�=�'?\j?>/>�ޔ>�I�b��^�*�7?���>Ʒ'?~�?��?4��yZ1��h��L�����P��t>�[p?��?��n>����d┿�����A8�����ϊ?��~?/鉽�+!?(�?��L?ǁ@?{&>_�d�?��&oD�yL�>��!?K�޺A��M&����~?�O?���>�B���ս�\ּ������'�?U(\?�A&?��+a���¾�3�<E�"��U� �;2qD���>Ï>���m��=>�Ӱ=�Om�*C6� g<�j�=��>��=�07��p��E=,?x�G��ԃ��И= �r��lD�2�>�.L>���ԕ^?��=�A�{�M��,z���U�Y��?4��?�k�?�N���h�"=?��?�?^�>�<���n޾�ྣrw��kx��r���>8��>��k�s�񏤿����|G����Ž5���M?7��>�1�>)��>���>�أ>��˾�@�o� ���'� �b�W��8��$����o���E��I���ʾ����&>��&=h�x>� ?Y��>"P">���>Gq=,�>b	h>ܔ�>}ǫ>w�->��>��=�lJ�H�%��KR?����%�'��������c3B?�qd?P1�>ai�:��������?���?Rs�?=v>h��,+�}n?�>�>I��Xq
?oT:=&8�X;�<V��~��93��P�,��>E׽� :��M�2nf�xj
?�/?�����̾�;׽F���m=v<�?�v+?��-���Q���m�Y�W�CvN�A�&��(c�����3%�'�n�R���N���^��J;'���\=L�,?-߈?����  �͊����n�{�?��i>v~�>	J�>�.�>(%>�|�n�1���\�� � �u����>�#x?�X�>��I?�;?D�P?_oL?꧎>2�>Q�����>���;�&�>_)�>"�9?�
.?-0?�S?�A+?@�b> s��d���fؾ�>?��?�Z?�*?-�?�օ�2ý������d��y��܁�w[�=䮾<!�ֽxt��{T=�)T>eX?n\���8�N����k>ˑ7?�F�>�t�>�h���w�����<���>b�
?M	�> �Hir�C�/g�> ��?�$��+=��)>�=XZ�����>�=Ԋļqc�=����;��x <(ѿ=F�=Q������;��;
�<L?>T?�Y.>��8>*�4��52��T�r���.���Ӽ�O>:���7�~ș�!z���d>���?���?�~���>��D�nB��}5��P�3��1*���,>W�V?�w_?uς?{f�?��?	t?p�J>����0�����h%?W!,?��>S����ʾ����3�͝?I[?�<a�(���;)�-�¾��Խa�>�[/�D/~����>D�������3~��'��?濝?�A�*�6�gx�Ϳ���[����C?�!�>�X�>��>O�)�y�g��%��0;>���>R?*$�>��O?J;{?t�[?�gT>�8��1���ә��F3���!>�@?ձ�?��?y?�s�>(�>��)�4ྒྷU�����������W=�	Z>2��>�(�>��>��=$Ƚ�X���>�(]�=<�b>�>:��>��><�w>�T�<aH?�Y�>t뿾���R������)>�`�t?V��?�c*?��=}��ŴF�>���m�>�r�?�3�?W�*?��S����=�lμ�����9x�e�><�>���>2ʕ=�Y>=6>���>���>I	�@N�6�M�@���?��D?�`�=�:ƿ=r���p�g����i<�v���`�R���Y��[�=#���M�(����Y���zn��qµ�
֜��tz��& ?�Q�=��=F��=���<<���;"�<B�P=N)e<�`$=�u���1<O�/�d��~놽�o1��7t<�P=���M@Ѿ�݀?f�M?:[1?%G?+2�>��%>���7F�>�`���?�}>�Ӽ�楾�6�������B����˾zc��l��C<>����6�!>\C>�P
>�<wŸ=���=F�|=��h<d)=�7�=F�=:�=��>ؐ>�,>(�x?e n��I���G~����&��>[�>�>b�`s?!�>r2��-�ÿ�Z����?�B�?���?t�?��3�Ƥ�>�
��l�ս�v{�[�߼��?> ̬=��k�$qL>$=����듿��w���?��@EN?��ɿ�$>d�;>Io>�iQ�h)0���X�*�X���b�U*?Y=���Ѿt��>��=8��^(ʾd}=Q�4>�dv=����7\���=�aj��]6=��u=�<�>�H>���=�龽G �=�D=�=�J>%:���B;�[�(=�=�=�X>�)>���>1�?*0?b�c?���> >l��aϾ�������>��=	԰>\�=�A>���>��7?g�D?BL?=@�>�$�=�>u<�>�,�:�m�|v�q��j��<��?�Æ?ӷ>i}L<F�@�9���u>��qƽ�?�
1?�c?�m�>�W�n޿��d'�},��B�<Q' >����8�ͼ�+=����������'>�>���> ~>6.>��=
4>��>ZU�=��лz�>��'���$>�	�<�A�=��8H>t෽�^��J
>#v���c;��<��l=.:�=��:���=��>V�)>f�>SҖ=����[>���N���=$R��}]C�3c���}��.-��l2�Ї=>!kS>�᪽c��	,?�f>��J>M�?	nt?�_:>uS�,�ؾu���p[�*�X�e��=MY>��P�{e=��`�h1P���ھ���>D��>�
�>v�l>�,�a!?���w=�⾚b5�w�>ł��a���,�!9q��>�������i�Aֺ�D?yF��F��=1!~? �I?��?��>����#�ؾ090>�C����=��1q�i��j�?�'?0��>W��D�=���xĽԷ]>�Ӈ�a�i����/��k�i;��`��>�y�����}�9��b��M?���?�|xT����>�L?� �?ȝI��;_��F�=�
.��J�>��g?��>&��>y��>3�9�_������bg=��?���?�
�?��=��=�1��qL�> `?ϖ?��?�s?��>�$��>"��;">N����=��>\��=��=O?��?��?����)]
������ �a��<�<I��=I�>'��>�px>��=�w=n�=Fw[>�+�>���>��d>CV�>�:�>C����U��L?R >z�1>H?R��>ԓ�=�+���E=�GX�#D?��H�ܒ�WOݻj����Ƚ�c5<�4�`�?�cͿjn�?wi>x����#?���^��i>��K>Y>4�:?�";>R��=��>Z=�>�6r>��?��>�HӾ�}>���*`!��+C�*�R��Ѿ3}z>.���S&�s��d����>I�m���b��j��-���;=����<AG�?����k�k�8�)�E�����?cQ�>�6?�Ռ��
��R�>���>�Ǎ>�G��H���@ƍ�`�T�?���?S�>�j1>��U?���>��<Ѽ>leY�����&X��V���I�>Ve�	]p�6+�NɽLvl?��?�`n?l���l�>�͊?vc_�p���t6�>�'�a�0��[Լ�A�>~��|!��F�����r�/C=A�n?$Ǎ?W�
?�d(Ͼm��>4?Z?��?�ؕ?pJ/?�OW?��)�j�F?�q�>��?y�??�@B?��C?���>��;:ǂ"�hs����>�*��Y����
��þg�k��*��	u<=)_�<�P��}&>�~������8���o�׻RwV�);�= L)>Va>I��>aF?�*�>�tF>:!1?�c=H�J�J�+�>#��%�-MK���ھ<�'�W.̼�,Z?~��?2�x?r�<-w.�g� ��k�= ��>H�L=��&>�K�>.�����o�ֽ=&��=�{�="�=��N
��&���0����9&>���>��8>�b<=����現�������=F���<Ѿ�\���eu�'0L��U�����>�L?�u,?��=%�ܾ����l�֞9?��r?|�K?��m?	R4>�\}�u�+�20.�`yK���v>-�)=+���ܰ�q��3�o��r/�Z��=T:�Tj��=B\>�k�Z�ܾy�m���G�{��x�==���ƍ^=2�
���Ҿ�|p�C��='>�;����"��4��93��J�K?�E|=�C���S�� ���>O�>ʮ>��C��W�PfB����R3�=^��>@'5>�e����ﾃ�G��J���>}YB?H�_?C߂?��j���f��I�B�^T��m��Q?��>LM?{W>J�=mF���c�7Cc�|RJ��	�>�e�> �!��NH�c!��:����'��
p>���>�i>�_?��M?f$?��e?��.?pX	?<�>��潭f���D&?�y�?��=��ԽD�S�.�8�iF�h%�>�2)?v�B����>�i?&�?�0'?��Q?��?�4>�� �ZV@��y�>�x�>��W�gO����_>�hJ?�m�>�X?}��?��=>�]5�?�����<��=�>��2?�#?�i?q��>��>�������=Q��>�c?�0�?f�o?xt�=4�?22>���>O��=?��>a��>-?�WO?I�s?��J?���>���<r6���;��SFs�ّO��l�;H<��y={��Bt�B?�b��<␳;����=��$���D�吼.��;rZ�>0t>���)01>ž�S��l�@>[K��6U���Ŋ�D�:���=uo�>��?��>�#�6T�=���>�J�>6��J1(?T�?�?n� ;;�b���ھǏK���>��A?h��=l�l�����L�u�Űg=u�m?��^?�7W����[�b?�]?�g��=���þ��b������O?��
?J�G�Z�>��~?A�q?b��>Of��;n�F��eCb��j�%ζ=�r�>qW���d�X?�>�7?�J�>��b>�!�=�v۾"�w�q���?5�?!�?���?%*>��n��2����'瑿�\?R��>l9���w"?���NϾ0���3���5�a~�����u��:즾&����u����=��?@zs?0Gp?~�_?���*d�D�]�:�~�.�U��Q�ݣ�nF��F�\C�;�n�q:��.����jI=cs�^?�S^�?��'?���H_�>3�������;�38>�:�����]�=$�\����=��b=/�V��f)��Ǵ�;B!?d��>V�>�s3?�N��!0���:���?��A��j�+>�*�>�<�>��>;� =N+��'쀽Ỳ�x���c%��3v>�|c?��K?S�n?2h� )1�����?�!�00�6i���B>�R>��>3�W���9&��W>��r���{����	�	=��2?&�>���><P�?�?�z	��b��I\x�t�1��R�<.�>i?�4�>`�>�нO� ����>��l?��>���>s�;��S{�F�����>��>zV?5�~>�)��m[�S���c��!�;��*�=�n?e��s�W�t��>�N?uN�;q�<v��>Ă���< �n���&4��>��?b��=̭6>�vž5����|�l΀�X�)?q?t�W
,���~>�K ?� �>ׂ�>�
�?��>$ҿ�������	?9_?�VM?F?�u�>4��<��Ͻٌ̽����*=��>��Y>��i=���=����Z�,%��l)=po�=fפ���ƽ :��ӼMC�<�4�<(�1>8�˿g�D��ݾMj��������p�w����_��ne,������6q�v��������r}�H�Ӿ��оV�)��4�?��?�����Q�Aӧ����������>=�t���u=G$�X����ݾ�ھ�ϾS����F�[c��g�N�'?�����ǿ𰡿�:ܾ2! ?�A ?7�y?��3�"���8�� >_C�<-����뾭����οG�����^?���>��/��v��>إ�>��X>�Hq>����螾W1�<��?2�-?��>Îr�0�ɿb����¤<���?/�@٤<?� ��0þ��S>ɭ?g	1?��>ʀ��S�8�#׾ �>.��?�l?cw�k�I�����a?�Ȣ=��F�U[����=o�	=��<>Q���^>��>D/��Ŗ�~b����>'�>��8�E?���Z�넁� }f>I�=�l��B�?SO���e���>�|'����=k�I?���>+_�=�?�#9��n˿�^��V?f��?���?i�/?������>7�ݾ�LN?&j1?�C�>L��X1h�h��=����R6��!�<�Z��<>�s�>-b>v��ɒ�U1=��T���&=o> ��Aſ��"��1�)� =��k�H*�l$����?�L�5u����E���P�#�=A�>"+>*�P>#	Q>��R>�/T?uf?��>��>��佛�r�ڻþ�@Ҽ�����;�:���D]%�%)���[޾�R׾��XF�'�r�Ͼ��<�h�=�R��K���� �:b�� F��[.?{#>�Jɾ�M��,<�rȾ6���:��v��I�;:2�{bm���?:RB?�ԅ��$V����j��j���W?�o�����Z���=�ټ' =K��>E;�=�^���2�qGS��0?A�?�5���U��{9'>��C�=a�+?�?�V@<=�>�$?);-������]>*�7>��>F��>�>�9��2@ֽ^?$�T?���ش��n��>b����z���U=<�>�r0�e㼍{Z>�ٞ<#r��P�����Y~�<'"\?
�>���XX�1ݔ��T���m%>�9�? J?��0?�?�iY?��>�\���l��>��"��"T?�v�?�B�=i)395 ��*���v#?�OE?e@H��jz��\���P����>���?F�%?-[L;/�������T(���;?�v?��]�G���X���Z��F�>ɍ�>���>��8����>M�=?�%(�("���G���u4��Ξ??u@F:�?G�P<l���R�=1_?o�>�zK�_rž���մ�"n=��>ㅥ��v�� �_�+��\9?&��?Le�>a���`��=�ؕ��Z�?�?U����g<[��>l�p��qs�<�ū=�	�G"����1�7�E�ƾ�
�Ϊ��T-�����>�Y@�x�L&�>A>8��4�TϿ���]о0Tq�Y�?@��>V�Ƚ"���x�j��Ku�6�G���H����;��>9(>72���瑾��{��i;��y����>AD��8�>TeS�iQ��9���]*<�C�>j��>z��>~���$s����?8/����ͿQў����
`X?��?�-�?��?.2"<�u��|��,�@�F?p�s?U0Z?�7'���]�n�?�$�j?�_��vU`��4�tHE��U>�"3?�B�>L�-���|=�>���>#g>�#/�y�Ŀ�ٶ�C���W��?��?�o���>p��?rs+?�i�8���[����*���+��<A?�2>���F�!�>0=�TҒ���
?R~0?{�a.��_?�Ha�?�p�)�-���ý�d�>�3��^�6������w%e��ۛ�@&y��?Sb�?��?���#�V�$?�Ư>�����Ǿ|��<�e�>���>��M>;cb��Wu>�����:���>r�?�_�?s?O��Oަ��>��}?�$�>��?un�=�a�>�c�=�-�Tl#>�$�=#�>�<�?��M?oL�>�U�=��8��/�][F��GR��#�%�C�,�>\�a?��L?�Kb>c���"2��!�UvͽZd1�DV�tW@�n�,�ܝ߽�'5>L�=>�>	�D�Ӿ��?:p�*�ؿ�i���p'�z54?+��>�?��8�t����;_?)z�>�6�,���%��[B�Y��?�G�?B�?��׾�Q̼�>I�>�I�>0�Խ����4�����7>2�B?���D��m�o���>���?�@�ծ?ai�ֆ?Qn���.��Z�_�)����U�y�&>|�5?ΖҾxÍ>�4�>��5��p��㣿l�z��?�>���?&��?��>j�g?Up���8��s8�ڦ�>FTd?U?㶼׾7�5>�c?�g�I����>�=e?�@��@&�a?�+��o�ѿeE��Iѵ�����B>9���J�> �;�V>�I�<�x�2�=�~>��>>�_>�C�=R��=Rϼ<
">h�z���2!��Z��@���5�F[�T"H��<������4�c����{���
���=����'S�/��)�\=G�=:U?vvP?��m?��?��V���>����<�/&�|�|=?F�>��0? N?G�,?.'�=�X��Ėe��`��G���B<�����>�<H>5��>���>'n�>��:��H>�K=>�~>" >��*=[	<�`�<W�H>���>�Y�>���>�C<>��>Eϴ��1��m�h��
w�n̽.�?���K�J��1���9��ͦ���h�=Bb.?
|>���?пc����2H?���y)��+���>u�0?�cW?-�> ��d�T�:>O��Ϧj�/`>�+ ��l���)��%Q>tl?g>�
u>Ξ3�h~8���P�c���W<|>+)6?޶��x9�Z�u�йH�7�ݾ�JM>���>��7�87�z䖿�~�Ǐi�*"}=5n:?!�?�n���Ѱ���u��q��3R>�[>�=<��=0VM>a�c�1Yƽ^LH��u.=2�=�&^>�N?'%'>�}=m�>����_�W�1B�><�G>��2>d�??�"?6d�"��ƃ��`{4�:�>���>Ԇ>��>�E�/��=
��>��G>~c���F��b���=���Q>�8����S�UE��~MP=4����>|�=*b����@�6�<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>tx��Z�������u�d�#=M��>�8H?�V����O�e>��v
?�?�^�੤���ȿ5|v����>X�?���?f�m��A���@����>:��?�gY?roi>�g۾?`Z����>ϻ@?�R?�>�9�z�'���?�޶?կ�?@I>���?՝s?�i�>p3x�
Z/�j6��ו�� �=x];�f�>\>{���XgF�ؓ�i���j�`����a>�$=C�>�C�4���:�=��J��3�f���>�'q>s�I>cV�>� ?kb�>���>8r=�u�� 〾������K?��?��b<l�q=E�=˽r�c�>�F0?_+��XzϾ���>�)Z?�y�?{5]?`�>��VG��DJ������!�<��K>r��>)��>������O>��Ѿ�9A���>(��>C���2>׾.@��*��y�>�6 ?~~�>�ݴ=y� ?��#?,>j>��>8IE����5�E�t�>���>sl?-�~?�?-Ĺ�xw3�����ѡ�DQ[�s�N> y?�??ہ�>bv��l���X���L�y��$��?�g?#]ί?�?؟??g{A?�e>���ؾ�H���A�>{e$?h���)�<�`�+��}��!�?Tq�>eF�>�z½����o��F�!�� �x�?9c?m�6?,��|Y�"�о���<s�<��HO�K�:�[>�A >��k��ix=M'�=�.�=M$W�B!&�d�<�ڼ=�V�>Pҳ=� >�y���,?����·��o=��q���D�_�x>q�J>�o��lX?�=�!^{��@��j����M@��s�?��?��?.7ǽ��g��=>?��?B�?!��>����l޾���
{�$h������>�ӿ>�^׼�B����L ��dm���s����?��?��?%�>Q��=�)�>�4���5�/����Yl�e+���<��\&���ek��ib��h���EǾ����fP�>v��<�ݟ>a?�M�>�˥>�-�>�E�=�g�>��A>���>{&�> �I>NH�=pG=?�z�P�<�KR?����"�'���辽���h3B?�qd?J1�>�i�;��������?���?Ts�?'=v>h��,+�~n?�>�>E��Wq
?GT:=9�;�<V��{��#3��%�-��>E׽� :��M�?nf�vj
?�/?
����̾�;׽`k��V8�=�}\?h:?�}C���K�,b��;��F�$ɯ=#�������ts�W�\�����R���Ď��|B��[�=Q�9?n:�?��辅T����ܾ�y���A�6��>���>��>"��>ܯ�<��>��$���d��"����Q�>�Tp?�o�>q�I?
�;?�FP?��L?d�>$�>ʳ�$��>�u\;���>A��>��8?S%-?�/?Y�?ȃ+?�`>Z|��������־�M?�Y?vS?0�?m ?0���Ztн��¼�Qݻ�q�+ʋ��<R=�)�<ø�3�q��{=��R>um?�~�:�8�����̙j>P7?���>�:�>q��>F���.�<t�>��
?Ύ>�> ��r�J��7��>�҂?g��"=e�)>�5�=K���Y�����=��ļ�R�=>$��\B?���<��=j�=Q�}��n!���R:.�@;N9�<	�?1.?��I>�j�>�BW�	鄾R�����=��=c�>6��>��ݽ��~��M���m�v�?>�=�?R%�?��I>�g>jD�<�)������S�.~(�6OG>�Vl?��?��?v=�?+C-?��A?)�>D|��L~�awd�O��;�I?� ,?ߌ�>���f�ʾ�d�3���?�[?�;a����,<)���¾ս��>�\/��/~�����D�4�����a{�����?��?�A�T�6��w辨����Y����C?�!�>�S�>=�>+�)���g�"$�w:;>��>�R?�6�>]�G?�j?��G?Z�>���N������Sܷ���=qr-?,�l?��?�o�?�/	?��>G=ӽ�����	�����~�ny����;ՅN>�]>���>X�>%7�=���������P����=��p>Q)�>��>��>�z>lD=tI?���>��Ѿ�
�? 侊1����=�h?�O�?6"?�&=3y@�{<N��f�͘�>B�?���?R�4?Ѵ�?�=eo�&��D��hh�>FӤ>A�t>Wz�=ռ��Z<2X�>�}�>>�Z�=��n�ž<��=G��>��?�>��3ÿ��k��������=�E�r�]$ҽ�?#�Cgn=%5#�/k���&X���н_����-��|����M���W��	�?nW>Q�;=A��=&�&�M@�=�v��G?��I��&tI=܋����ڻ��=D��Xj �"�< O@�`�;��t�=�˾�}?�;I?�+?��C?�y>�;>.�3�~��>�����@?�V>+�P�Y�����;�B���u ��"�ؾJx׾��c�lʟ�II>{_I�Z�>�83>�G�=�Q�<f�=s=QÎ=r�Q�\=�#�=�O�=�g�=-��=*�>�U>��v?T��˗��mLP����*�4?�A�>��=a���>?�=>��� �����Oz?x�?��?��?$�d�77�>�%��W���.=y��7�/>�ǹ=��-�x@�>[�8>���˛�VS˽���?W5@ì??� ���ο��>�8�>���=�T�DS�����<h��0��v&?P�)�g�ƾ�Ί>�ӻ���������M�=/L�><�>�r���R��B=����<M4=_,�<�щ>g�4>=�=m�ʽ�Wo<�i'�aW�=W~�>���<$M�;(�k=��9=x��=s�8>���=���>�'?��,?f�h?��>r,A���̾�Fоmh>9�=�K�>$��=�2#>~�>�4?o�B?��M?��>@�Z=���>���>I�*���n��侯�����}<J�?zֆ?{ȸ>+Ù<�=�+���k:��3ս;�?�.?�?dT�>��q �Z�7��7��B����j���=\�ؼ� o>�9�l;��{e>��>q�?{?i��犽t��>e��>$�>��=F
�<�~>
j;�j�=݄=�@������Xֳ<�b�=9c���I;�. >��L=DҞ;U4W���>�Ao��c�="�?��U>E��>Ӳ�={f¾o;>!���rQL�7-��ܾT:F��9g�y/��ur$����&9>ʏ=>#�I��]��d7?���>gٍ>M
�?=5a?ϊ>����&徫 ��]����-���h=���=in���WC��k�!;W��������>��>���>��l>J,��%?�eNw=���^5���>����9��:��2q��@�������i��8�ڟD?$@��ߢ�=} ~?��I?�ݏ?�~�>���7yؾ�D0>N����=���Lq��\����?�'?���>���!�D�ڔ��N�<\ p>���=r){�����6�=��=oR�� a�>.Ҿ�}��!3�^��ʗ�rIA�
� >DCM?���?D�����D��� ��?�b*S�=?�F?���>V��>a�?����������r��1�=�?���?G?�?��=ZX�=#����>��?��?�S�?Ɣp?��f�1��>��o�5>�Vh�H��=)��=�`�=�A�=}�?S?Z?�1���Y��$�)��cN���j< ��=-�>C�>H@a>��=7�r==�y=�A>�> ��>�Yl>�i�>���>́�EC��8�z?��s>N�>�2?�9�>���=؛�����e�l�z��\��ؽ0l��FM+���0�~}��1�� ?�Jʿ��?�>"����W?Om)�N�VT>h>}�Z;�(?���>��>;��>�<�>���>FB�>�k�=YPӾs6>���o!�=RC�k>R�pѾP3z>�t����#�L���X���nG�!���a���i�q[����=��c�<�J�?6����Rk��*)�5� ���?w�>�6?�����o���->@�>���>�j��P��������~�΋?��?��>U��>��f?u[?C�_� 5�c�m��9y���D�k�U�X�X���,�n��AҾ��
=&_?��y?��,?(;ڽe�>��}?��Q��K��ƞ>�T���P��^�X�n>���<�н ���u��j�O==G�>.�?K�{?�6�>V�f���m��'>��:?%�1?�Ot?��1?��;?����$?�n3>�F?�q?�N5?��.?�
?62>Y�=ma��"�'=�3��J�ѽG~ʽ�����3=�]{=�>ڸy�
<��=�<�����ټK�;}<���,�<�:=�=�(�=��>��Z?���>)�>3�F?���tB�]`쾦S?���b��p��h����Ѿ�76>DCi?���?t}C?��>��C�PB�/�>*��>Q�1>��f>1�>fԻ�rFL�%�<s�*>5>��?=�^7��9��]
�_�j�r��= b4>?�>��z=�}5����%������"�վ����:�c|"��֙��0�>�A?B�'?��k>��׾6��s�`��07?;�R?�j?��y?��*>s+7���9��K����-�=B�>���;��4�����`���ս��w>��ɾ~����0b> ���ݾ7�n��J���}*T=N|���W=�*�e־��U�=��>����� ��	��<����~J?R�o=b���7�S�>麾?^>�>��>z�7�j�y�&@�!������=���>��9>�Ɵ�{�PG�x��]>�>[QE?:W_?k�?"��Ns�;�B�o���Vc��!ȼ<�?jx�>(h?�B>@��=U�������d��G���>���>Z��;�G��;��~0��C�$�
��>U9?ϩ>��?N�R?x�
?u�`?�*?LE?@'�>�������B&? ��?��=V�Խ/�T�) 9��F�;��>�)?
�B����>�?ѽ?\�&?e�Q?$�?R�>� �uC@�Ҕ�>?Y�>B�W��b���_>x�J?���>�=Y?�ԃ?��=>Y�5�0颾�۩�7O�=�>_�2?�5#?/�?��>,=�>�����=��>�1c?떃?p�o?)"�=?�?��1>���>$�=�	�>���>��?��N?�hs?�%K?��>�e�<����R��_�v�SL�+Ӎ;�6D< ~=����:|�5��O�<�!�;rݵ�[Bv�8��̦A�8�5+�;c��>�xr>=����2>��þ����+�<>��ż*+��y��o:��=�р>��?.}�>Q: ��Q�=�^�>w��>[g���'?C�?�"?�8(:D&b��wھ�lG�կ�>sA?(�=��k��Ĕ���v���b=��m?�:^?�YW�������b?��]?~m��=���þ��b�'��]�O?5�
?}�G�V�>'?\�q?e{�>�Qf�3Tn�����Gb��ij���=��><���d�O�>�7?�'�>��b>�a�=H۾֫w�j����?��?���?@�?��)>��n�P.�Gx��NC��
�]?M��>�o����"?�Q�p�Ͼ.Z��
�������L
���C������&%��胾�a׽��=3?� s?x?q?��_?� �d�30^�u���XV��&�)��E�<5E���C�M�n�Ph���������H=X�I�`H��O�?g�'?�C����?j�����Uo��[�=����"�-�=3м�>��=t�B��Nƽ4�����%?O�>|�%>:M=?q^7�y;��L�K�b�An��]W>��>�x>��	?�
P>���</ර4����H���C��)v>�}c?��K?>�n?�\��'1�����!��l/�R\����B>�v>6��>��W����:&� \>�-�r����|��p�	���~=�2?g'�>���>:N�?J?lv	�!j���\x�l�1�ك<�4�>�i?�E�>��>
�Ͻ,� �	�>�
h?�l�>z}�>���������v����p�>�>�X?6�>"@�Ԕ^� B��pV���G�q0F=�Ro?����6�[Ώ>e�Q?�c=;͓< H�>�;���|'� �L��s��=�8	?3��=��]>(�˾�s�m�Ut��F)?(=?�ޒ�$�*�T~>�#"?��>;+�>�*�?�5�>lþ��:��?)�^?$:J?UA?�L�>�)=�ı�-.Ƚ��&�'�,=]|�>�[>tm=�N�=o���\�ϕ��pD=|ź=�μ�)���<�޴���K<���<?�3>�.Ϳ�S�.��D����R���s��;=@¨�#�ҼZ5��<����Bٽ߯�&#���������&9|���~�1��?�A�?�lϾCa\�!I��k�n�0j���
�>�9��՟A����Ka��)���f��3��c?���2���N��g*�O�'?�����ǿ𰡿�:ܾ2! ?�A ?9�y?��5�"���8�� >RC�< -����뾮����οC�����^?���>��/��r��>ڥ�>�X>�Hq>����螾V1�<��?6�-?
��>ǎr�0�ɿb����¤<���?/�@o�@?�������/�=�_?<�*?-=>RJ����6�������>'��?�W?1�Ѽ��9�q��<��o?֓6>��c�D�*�G>B
3<I�>� p�rle>bU�>�I�mZ�����ٲ�>i,�> 	�%}'��<�����rp>j�7=��X���?��Z���j��8�.����y�=�{I?&�>�u�=p�?�sC�ʿ9�a���S?V$�?f��?�7?ʎ��	�>�ᾔ�N?ا8?�h�>�����k�^�<ƕ�������� �w�[�O�=A��>p/(>�µ�]�=�B�UL���y�<�����ƿ�J#�hv�B�1<�AZ�Ù��a ���B����	�zaw���I��$��=�>?�=>�lc>%�8>��;>�5h?�Xb?�W�>��/>�'�TUf�Q���Y�-<"����۽ɨ���ِ�������侘Ծ�~��$����ǾM=����=�HR��q���� ���b�ۖF�2�.?$>�ʾ��M���(<�Sʾ�Ī��߈�<���=̾�1���m��֟?WB?9ϧV����I
��S��"�W?N��K������,�=蹼'�=|Ɯ>���=;��3� <S�Yz0?�\?>���!i���*>#� �g.=i�+?��?v�X<�0�>�\%?@�*����o[>�33>���>P��>z	>>'����ڽ�?i�T?\��H����Ő>�i��[�z�Ba=�2>�K5�v���[>���<}���<>[� @���޺<�l?�ǽ=$�7��c/���fʒ��=�?sx@?d��>eb�?�V?=(��pl��χ�6�,���H=Y�&?h3m?�Q=�j^>������&��[<?��??@^.��sC�o}���F��Uھ�F?�c?�.�>���"��?L���aK��=?�mx?�[b���������.�>��>���>�-�A��>?0?��p��l��y���Q	)����?�+@hK�?�Q;!��ڡu=:��>�[�>��%��ʩ�i/���o�=�=�>N]���H]�L	��.�tP??u~�?&?��o�����s��=ڕ��Z�?v�?�����]g<I���l��n��w�<�ͫ= �4E"�P��@�7��ƾm�
�m����㿼��>Z@B[车*�>�B8�>6�1TϿn��K\оsRq���?̀�>�Ƚ噣�m�j�Pu��G���H�礌�ڼ>�Y�=uڽ����@�m�=�4�a�=���>�J��;\>�H����퍽�;Ff���>y$�>Rʱ>z�<�پ1�?��
���¿����.h2�F�?%��?��?(�L?̴h>;���O���e�;=ft-?�D?��N?�d[<	�N���Y=0�j?����=`���4��E�rT>2?���>;�,��Ky=\>ʳ�>y>�E/�T�Ŀ�������w{�?Mz�?���C��>�e�?��+?C��.��������*����A?�2>����3!���<�i葾4Y
?Ċ/?(!�=[��rW?�a���[�s ��&�=F��>ӱ���d���N��N�$IM�#�����ǽ^�?!�@�?i���G�4?��>J�;�~� ���=>�>~>>S��G����1>�$�Vn�M ����?���?<?�Ze��]���@��s�?(��>��?*>�?9R]>mMξ?�C���a>'ڙ> >�=f%?�Y?���>��4�����``�%匿�Tg����
q��>'�{?��[?=�>g\�oѽ<]��s�����;k{����՛=��s=yKk>3��>�zC>%�,��ξ��?+p��ؿVi��v'��34?m��><�?����t����:_?&x�>17��+���%���A����?�F�?��?��׾^T̼P>��>nI�>�Խ������7>B?d#��D����o�#�>N��?�@�ծ? i�n�?�.�A싿f�w�qv$����o?>�
1?Π�KSb>���>eX��v�|�%����i�_R�>���?���? �>}=f?_t��1��
��>ӹb?�?#�3�M��z�>X�>1��ܝ����־cBl?9@�	@��_?����(hֿy����I��Ƙ�����=���=�2>T�ٽxf�=��7=��8��0��I��="�>�d>�q>�'O>�`;>��)>+����!��q�������C����}��Z�t��Rv�:{�12��I���B���5ý�u��4
Q�[3&��2`�̶�=�}Y?\�S?�r?t9?�zn�s�>9����p>=���3��=�@�>�3?6�K?,c'?���=嶡���d�=:��©�D:���[�>�HI>\��>���>i��>`�x:IL>�h;>�>���=5<=�;�;�/= �T>�?�>�m�>�δ>�C<>��>Eϴ��1��r�h��
w��̽0�?����K�J��1���9��Ѧ���h�=>b.?�{>���?п_����2H?���x)�ѹ+�|�>l�0?�cW?,�>����T�;:>4��ަj�`>�+ ��l���)��%Q>tl?��e>�(v>Y�2�G8�vWP�K���:�{>��5?핷��;���v��"I���ݾ�oK>��>`�?�Y��2����D��-k��A}=�:?[�?�Ǵ�
D��
t����VKR>*\>��=��=�pM>��d��Ƚ�oI��%=��=�:`>�]?̯+>"2�=���>�x��yOP�>��B>�,>�@?�%?�$�{E��������-�]Mw>e�>� �>�Q>Y\J��!�=�i�>��a>����ك�K��U�?��aW>*�~���_�~�t��x=����AD�=�G�=Q ��=��q%= S~?q-���׈���辗q��1D?�<?�d�=�o<Z�"�^���8g����?@7Ț?d�{�U���?Ib�?�\���t�=8��>u��>�ϾiL��@?�P��H砾G
�p$�"�?�ݟ?E�I�ރ���@k�Mv>�}$?�־Lh�>cx��Z��|����u�ѵ#=#��>�8H?�V��a�O�u>��v
?�?�^�ݩ����ȿ+|v����>N�?���?[�m��A���@�w��> ��?�gY?Moi>�g۾W`Z�Ë�>��@?�R?��>�9�2�'���?�޶?ͯ�?=I>���?�s?�k�>�/x��Z/��6������q=��[;�d�>�W>C���kgF��ד��h��|�j������a>͗$=)�>�D�K4���9�=���H��պf�B��>�,q><�I>W�>w� ?b�>���>Dy=;n��4ှ������K?���?*���2n�jO�<���=|�^��&?yI4?<o[���Ͼ�ը>׺\?h?�[?,d�>4��M>��E迿.~��.��<��K>4�>�H�>�$���FK>��Ծ�4D�Fp�>�ϗ>[����?ھ*-��E]��5B�>�e!?���>�Ѯ=A� ?��#?�Fj>s,�>�lE�,9����E����>b��>)C?t�~?!�?>ӹ�Z3����꡿Џ[�w N>��x?�W?Uϕ>�����x��)�E���I��
����?Zig?�彔?�)�?�t??��A?�f>^��ؾ����q�>�"?�6�2�A���%�u��B,?�?�#�>�i��1�ڽ�"༃0�����o�?D�\?w�&?�����`�G¾6B�<NE��9�8�;36K��>�>�큽\��=�y>d[�=��i��V:��?<}��=k��>W��=��5��w��q(2?�z�-J���;��)n���L�f}f>�\D>H����=?�v��{�ة�^i��C���Yt�?M�?���?�u
�]jj�m�A?�r�?�?�{?�����������%�������"#�O��=v��>*���ZNܾѡ�Z��z/��6u;�U�I��?i��>�R�>9�>"8>I{�>^��1�au	��h>���v�>�!�*;�Ȕ(�z
����0��`��1�þ�à����>��<}M�>>�'?O
�>ᮝ>;��>��<�R�>�>�a�>��>�,;>j�=���E06���R=JR?����2�'�z������/B?LQd?*��>��i����d���m?+��?�}�?ΐv>�eh��%+�o^?�S�>}���l
?�G:=����<IQ���������t����>]`׽]:�}M���f�`
?�*?�0��܍̾l�׽�q��Y�v=�a|?�w)??U2��OR�a�n�S�J��=Q���缹-u����!���m��7��>���
ӂ�X?*��AI=��0?3��?=��l�ھ(µ���o�pY?���j>5��>Kɋ>U8�>pRB>)"��#1��]���&�
{����>�Xz?�r�>D�I?�<?�oP? gL?
Ǝ>Wu�>/��Eq�>J5�;���>\�>�9?��-?�/0?t?�k+?<"c>v>��
����ؾ��?�?�A?]?��?�煾ȁýY��.�h�}�y��P����=��< �׽l�u�)�T=�T> Y?Q����8�v���Gk>Z�7?��>a��>v��i-����<	�>۵
?{F�>O � ~r�c�dV�>���?����=��)>���=S�����Һ~Y�=����=�;��Xz;�[k<O��=]��=�'t������v�:���;�n�<D�?�?e�Q>�Z5><(��A'���ܾ6)>�E}>�Q�>X�L>��ӾvK��	����j�I �>p�?ڽ�?���=��=3�=�s��G��A�	��;þ���#?��+?��V?��?�C?�|?��>K<&��+���z��hJ��LZ ?�!,?>����ʾ.�N�3���?�[?b:a�`��8:)�2�¾��Խ�>z\/��0~����D��A��=���r�����?ſ�?�A���6�&y辎���j]��-�C?�!�>�V�>��>��)���g�5%�+*;>��>w
R?UG�>��:?'L^?E�`?T�>��&��⳿9�����ƽ��=�3?�_?'}�?!��?B� ?O6_>̜&�U2�q����M���W���Yd�<g�>~!z>/S�>���>�*>Xr���V���n$��7=�"9>���>I>�>��>�*>�ж�VLO?*o�>DоK"��˾򡙾k�=Ōp?+�?5�!?�p�=���oM�v�rY�>�-�?
��?COC?� s��)�=� ߽;K���7�i3>��>��>�W/>9�J>L	�>�"�>��>N���Z�Q�R�5����?t�=?m%K>�ɿWu��{o�h����4<�E��3m��o��J��ª=mn}�U�ѽ����ܻJ�阖��I���n��������w��=?�w=��=���=<��:�*��0t�<��p=͘���6S=�ٜ���<��< �*���҈K��&�;�G�<-�G=���X�{�?�*n?��P?�kI?�X>�8>@��<Mg?�h�=�?ɝ�>y�A>���
h2����d���"�پ3ˏ�"(��b���4>��ҽ\�=�1>7c@>�S~<��=T�<J�0>o�g�,�~=�l>�+6>�_>��>\gO>:h}=�"x?ꁿg,��FWV���!��`/?�Y�>q��=v��_:9?�T->���������	��ny?	;�?��?3�?�e�*j�>I���� o��2�=��;�21>D��=�x2���>�g->���y���<��H5�?��@�aB?�儿��ʿ2I>I�;>s��=�JS�|2�*�a���c�]4W��!?��:�7/̾�#�>��=qZ��~ƾ�T2=��<>r�y=���b�[�7R�=,Mu�J>=�Uf=�Պ>@�C>�D�=k�����=Z�==��=E�Q>J�����*��C���H=:v�=�_a>��#>?Lz�>P��>�PU?�_�>�؋���A���+u<!���«�>9h�: ��=�s�>��X?I�M?��D?�]�>����EX�>U�X>�"�t��!�"�����-�=AA�?}��?��>��X$������X��U5�v��>�^?�j�>>�=�~���ݿ�R ���6��2��Q�q��F L�l
��M���O ���9[AB>�4�> ˽>-\�>l�4>���=�.>�u�>���=���;~�>�UN�0�X;�g����=Y����ݘ=�>�V����0[=V�+��w<�/�<w�:;6C=�޳���O�=�w�>�9>�T�>��=�_ƾ@�>m���S0R��M������)U�Fvh���v�� $�IM �5P{>FP�=?Y��G�� ?̥�>aeP>�#�?g�v?t�D>D���;t����턾�w�-�=��=�-���{E��(d���Q��ί���>E�>�F�>��g>��*���=��7V=S�ܾs1�IB�>Ա���÷���q����#��Ml���$�i�D?����i�=�6~?��J?Qz�?s&�>�ޠ�˄پ��$>�Iv�d=E��L�i��ˊ���?3:&?cc�>���pF�ޛ���i���H�=ܣ#�,�z�����,�Y�>ο��J��>NE���:�o�4��=���Ō�<\U���i���>�kE?���?V���W�d��R����$�n�?^K0?ξ�>��>��
?>�t�~��]��ִ�=4h�?Vl�?2
�?�D�=oO=p�w����>)��>���?�(�?}us?�M�M�> ��<l�&>Z!μ��>(�=�~�=�&�=�T?��?q?��m�����K��O:�I�j��~<��>ٿ>h�m>-�>��=���=v�=��E>!S�> ��>��/>��>��>�-��4���LL?�}Ļ���>дV?�>>�'����<��e��H������Aνb����_"<�W�ѱa�|?#=��?�sĿ)�_?r�>�����|7?����9�
��̂<���=�@�={t?'�>di�>m�>G_�>�>��>Sn->/�̾N4>�r����[�L��S��y׾@�>0�#�wW
����p�G��󶾳<�8q�&�����>��^=O�?�����i� �B�Ǽ�>M9�>D�3?��Ʀ��>�%�>A@c>�����$�������.׾좆?.��?"�c>ၞ>N�W?��?�:0��&1�jZ���u�hLA�C(e�p�`���������i
��k��=�_?��x?>�A?e��<�3z>酀?�/&��.��$z�>�.��;�,�3=�a�>����^��dӾOTþ����G>�ko?i�?s}?o�U�8ܾ�Ԝ>�E]??�?��J?�m?zbl?����)?q�?�>k�?�wY?�?�8�>��=g��`�<�C�>���)�Ͼ�'��|���?-��N�=���=�.n;]׽�*=��=ٟy=,4�.$��`�:�R�<7U�=�6�=/x>�-�>�:Q?^�>+��>0A?rɼ�/�Ӂ׾��?_q��to<�l�n���̾W���Z%>�^e?�ʫ?��n?e��=g�>�kA&���=��>��>�&1>���>Wؽ�(A�Uax=[�N>�!>o�t=h�E��V��]Y���I=_|,>�?���=L��h =�!4��)�\�����*�8Z�3����QH�>=�Y?a�>?�V>�߾4�Ⱦ�[��a$?z�H?K�?�[e?B9O>�xS�"���<��$��`�>�i�=t;����7K���"C��� >Ze�>��aߠ��Cb>ݽ��u޾�n�5J�����FM=��{V=��~�վd.����=*
>������ �}���Ҫ��3J?Evj=tw��ZZU��t����>���>ޮ>��:� �v� �@�
���U#�=��>�;>hq�����:}G��8�c>�>+QE?W_?(k�?�!��s�k�B�l����c���ȼ=�?�w�>�g?BB>���=q�������d�mG���>Р�>����G�];���0��I�$�Ŋ�>b9?/�>��?��R?&�
?p�`?�*?]E?�'�>������B&?��?�=��Խ�T�< 9�OF����>'�)?��B�ӹ�>�?ǽ?�&?�Q?�?��>ϭ �cC@�Ӕ�>_Y�>��W��b����_>J�J?L��>�=Y?�ԃ?)�=>J�5��颾ة�aR�=�>y�2?6#?W�?Y��>���>����jQ�=r��>�c?�/�?��o?>��=)�?�62>@��>N&�=;��>���>l?�RO?W�s?��J?N��>;&�<*v��	T���s���O���;n�G<��y=���t�n_�Q|�<��;T)���v��(�񼽞D��y�����;R��>Fs>�&��g-2>�Pþ����/>=>sż�ӝ��ڋ��8�,I�=L&�>�{?�_�>X	"��h�=3n�>�|�>٦���'?RX?��?��	;�)a��dپuyK�l��>��@?3��=�l�s���1v�j�g=��l?�^?��W����@�b?��]?�a�=�=�þ��b�����O?n�
?��G�[�>�? �q?چ�>if�uGn�����Mb���j�1L�=׍�>�5���d��K�>�|7?z%�>��b>²�=�w۾��w�&j���'?��?���?+�?�)>��n��.�C$���2����S?F��>��@�?���򗿾
Q��WK�n�߾��������2j��2Ė�r�8�Cn��#�R.�=�S? �z?�#m?�f?tx ��ck�{ph��9q���T�����T��SB�N��B�Ccl��������Ӈ����<�.v���@���?�&?'�?�>ߑ������"Ҿҿ/>�k��ɖ��?�=[9��UrO=Itg=��f�Ω$�[��]Y ?2��>)��>%{??�bU�,�;�"-5�9�;�����c>>FL�>�	�>�	�>�W�<~��d���l�¾����e��#5v>�xc?T�K?��n?�B��1�B���؜!�EG0�'j����B>Zt>2��>АW�x��I8&�P>���r�����}��`�	�7E=8�2?�,�>�˜>�K�?�?�}	��h���<x�x�1�偁<U"�>�i?�2�>���>��Ͻ�� ��L�>�j?Բ�>~2|>�؇�Oq ��lj��<��>(��>�b?�U�>����X�������C�?�JaF=��d??���2Ƚ�}�>�BE?:��=�{ �K>՚�L�%�����&/�}�C>μ?>�=��F>6fžB50�	V��d���a)?�?K��E�*���{>��!?��>�5�>Z �?�ԛ>yþ@�#��K?�^??mJ?�A?�^�>��=�屽�ǽ�&�3�,=�\�>-[>��p=R��=����%\��~�QD=���=�żK��Ǹ<"=��)�D<Sa�<�4>9%Կ��L���־�C��R���t�W�o�:�v��ڔ�;��&���󩇾�|4��+�g,z�$!h���t��g��"�g�n��?G{�?�˂��5�)畿�Ђ�������>�~��<+�� ������ε��?��3��e�,���K�NYa���a�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@�d@?!�$���h��=���>��?&� >�Ac���&��ﾾ�p�>�S�?���?�-�=˿K�����%�e?9-|��eN�w���F/�=�b�=�K�=�t���i>�=�>"�*�G	^��'�-�b>�т>b�Žs�#��(L��-�<�7t>1vֽ���J��?��L�ln�	g^����*�=��S?]�>���=��>��=�d�ʿ�
R�Q�L?t��?f,�? ?�����l�>w$����A?[�0?���>Fା[L@���սb]��c�ھVC���>֍	?&�V>�ȽE�e����n��?<>�������4e �C����3<�ŉ=��4<�1���-�+�y="���*mB�~�����<�2$>�6>��I>7(�=wf>Kk?�"]?���>�H>}*�辎���l�<�X��� �Lv�����쬥������Ѿ���r��6��Ӿ��<���=M<R�����	� �F�b��F� �.?)s$>��ʾ��M���$<?�ʾ�ڪ��݈��v����˾�c1�@�m��?ϴA?�����$W��"��)�u!���}W?�d����E�����= ����=��>5�=+��h.3��vS�v0?0^?d����^���$*>�� ���=��+?/�?�UZ<�)�>�P%?��*�eM�hA[>�3>Yˣ>���>,B	>���L1۽F�?a�T?4��B���3֐>d`����z�`�`=�*>P65�����[>���<K���ʰW�[r��?ۻ<e\?u�>}�,������ھ�]S���V>�b}?0�=?�R?��?�aY?�-9����է����ӑ�>u��?B�i?[E�=�(>����,bJ�ĞI?aE?kM��O�Ⱦ��-�Tn���	A?6C?�?	,2�����}��8w<���?��v?)^^�9k�����:�W�3�>��>���>��9����>Ԋ>?P#��?������d4����?��@���?��?<����$�=� ?6%�>G)P��6ƾ�㲽�`���s=�N�>XN��pv�����s,��Q8?��?�o�>(m��������=����7z�?�,�?�����xB<���@j�c �/'�<Tr�=|��\$�@��6�xiɾmz�R��(Ӽ�O�>#O@��佇Q�>�6�zh�R�Ͽ����"Ͼly�-k?X�>(�ܽ󟣾�j�Dqu�]5G�k�G�[芾�K�>�a>�&�h����|���VQ�X��0'�>��@�n>��mV۾ÐԾ�_y�~�>��>7��>��<�����r�?�
�uĿ�����'��L?�"�?]fb?~%?�tF���Ǿ|̎�(��e�'?�Ԁ?�!o?�L�Or�����%�j?�_��tU`��4�yHE��U>�"3?C�>-�-���|=>���>g>�#/�{�Ŀ�ٶ����Y��?݉�?�o�&��>h��?os+?�i�8���[����*�	�+��<A?�2>ˌ��2�!�+0=�RҒ���
?0~0?N{�\.��Y?�vQ�`�O��(���m=��>Ş����پ}��vX���I�����\�5´?v��?5Y�?�����"7/?e�>�Aw��}���w@>���>��{>jɽ�z�`��u�>� ��H��{�9=Bi�?B�@?v�������|����?Q��>{ɔ?d�Z>l7�>#>Wa������>`��>1ü֑?I�?(�?�v�F����k�Bt�^4a������T�H��>3&�?�L4?yӎ>��~='�=���˭��ƽ�r�^�u��˵=<��; }i>9>K�G>��������?Lp�9�ؿ j��#p'��54?.��>�?����t�����;_?Nz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�>:�>�I�>=�Խ����\�����7>0�B?Z��D��u�o�y�>���?
�@�ծ?ji�*�	?z�����,	|�j��4�Q����=�[7?̗���y>>��>E��=��w��\-v�ز>.��?���?`r�>(�l?J�o��C���9�1�>N�i?Ҽ?k^�1�ﾫ�6>-D�>?N��=�����3�e?,A
@L�@bY?����ʿ�֐��ϲ�I��٤1>+N!>�e�>�Ә<�k�=�"=�UȽ7��=�C>eӓ>?�>j�>g�q=���=?m	>��w����-���Ǉ�	e-����ʍ��NQ��Rؾ8Lܽ%{'��߹�����_��]�м�����GW�0&��,ڽ��=#�Z?�W?+gn?:?âb��$>���^I=ѷ�e]=��>��4?I�H?H #?� L=����^�c��E~�_#��Pԇ���>WH>���>շ�>s��>+"S9
T>�|I>$>n>�n�=^].=bUb<�*E=�S\>�3�>��>���>�C<>t�>Dϴ��1����h�8w��̽'�?g���L�J��1���9������h�=Pb.?�|>����>п[����2H?/���n)��+���>��0?�cW?�>����T�:>=��h�j��`>.+ �l���)��%Q>pl?D�f>Du>��3��g8���P��z��ds|>F/6?�綾oT9���u�ԵH�3dݾ�BM>Ǿ>1B��g������
��yi���{=�z:?��?!��װ���u��>��	>R>q)\>l.=�x�=�^M>T<c���ƽhH��.=��=!�^>�X?��+>���=�أ>4g���IP�v��>�B>�-,>�@?:*%?�z�a䗽ቃ���-�(w>6V�>R�>�`>�XJ�=��=�k�>@�a>6D�콃�?����?��pW>_~�
�_��Mu��x=�*����=��=�� �v=�,�%=l8~?`ۦ�OI���m��	��D?.
?)x=���;�"�!F��;W�����?��@�S�?���;V��n?P��?�3�����=���>6�>�fϾ�K�#?0���>����u
�� ��L�?G;�?CV��O���<k�o�>� %?I�׾Qh�>yx��Z�������u�Y�#=O��>�8H?�V����O�a>��v
?�?�^�੤���ȿ2|v����>W�?���?h�m��A���@����>:��?�gY?poi>�g۾=`Z����>ѻ@?�R?�>�9�x�'���?�޶?կ�?I>���?��s?�j�>+x��Z/�6��Օ��Â=��[;gf�>�`>����(gF�!ؓ��h���j�V��^�a>��$=�>
9�U2���>�=�����I����f�u��>8*q>��I>V�>
� ?>b�>���>nx={t���ှ(����K?z��?&���2n��S�<4��=ֳ^�P&?I4?By[��ϾWը>��\?k?�[?d�>��C>��7迿6~�����<D�K>W4�>�H�>X"���FK>��Ծ6D��o�>�З>�����@ھB-���M���A�>�e!?\��>Hή=b� ?i�#?�j>s&�>�^E��F��BF����>>��>I;?N�~?��?N#���Q3�C��M֡�	E[�w�N>6�x?Ec?���>��������aQQ���H�kߑ�j~�?IZg?����?H�?Hh??�A?��e>�����׾#���ˀ>'�"?�d�'B�~�$�	%���?)!?w��>"t��y �f<���!�E��?&�_?�*?R����]���˾��<S��ڤ�87A<�j��$1>L#> B���|�=w>���=S~P�%�*����<��=�k�>�F�=K3�.���G,?u�J����~��=�r�B�D�b[�>�M>Fb����^?d�<�ԧ{�����������U���?���?
��?~볽{uh��=?`�?| ?��>:��A�޾W��~�v���w�-3�86>%��>�&e��%�뢤�����~1��4OŽ���	?�?zA�>��>�j>���> ���w:��h�Q�3��Bf���T['��9���6n˾�~N�*̰��)��h�����>���(��>@Z	?�"�>`u�>ؿ�>]�����>�>��/>�͓> �>�Zf�{T
��-=���HR?a����'��]辭=��-B?�d?�w�>l�k���;���P?��?y}�?��v>�<h��+��A?�d�>����g
?Nu8=/(��7�<�ܶ�����2��N���!�>_ս��9��cM��g�bG
?�?�>��-q̾�*۽4,��n�z=��l?�i@?)���P�M}�\/0���U�_ӗ=5�L��;��1��l^r�W4~����B]��{	?���<�9?�ה?)M��p���(���샿��X�}�s>���>���=���>�M����.����0�f�Q=$��PO���>CCr?S"�>��I?�f<?�`P?�sL?T�>J>�>�ޯ�4��>T��;�\�>Fh�>E�9?e�-?�/?�?�F+?l	c>u_��q���یؾ�?ܖ?�6?C8?�?����9½�\��@ e�}�z��ԁ���=���<"�ֽ�Ss���X=f�S>�X?����8�����k>7�7?��>���>V��	-��b�<��>�
?�F�>~ �=~r�c�PV�>���?�����=�)>>��=⊅��ӺY�=������=�<��xz;��k<���=���=�<t�������:�}�;�i�<�n	?�?�:>�(>�dǾ�
�HM���hU>s��>��>e�T>�C��յ���7����s���>ʄ�?!p�?��=+ �=W>����W%����5ָ���C;�f�>u�!?9jY?�%�?o\?�$?Q�>������4�y��c��&*?e!,?7��>c��ǳʾ�񨿣�3�Ɲ?3[?�<a����;)��¾��Խ��>�[/��.~����(D�&酻���7~��:��?׿�?�A��6��x辬���8\���C?�!�>�X�>T�>.�)���g��%�`0;>���>#R?���>��!?�0V?m|?��>Y|����(q��%�.����=P'?�8+?���?�z�?�>?��m>	�\�S��y�g�/͕�~���ϐ����A->a8>�(�>��>�]�=q��<s���d�,�]=5�>�۠>js>�ֲ>l�s>���M?��>ۄ־D���ھ����)>(��?-=�?`�%?�1c=�.���F�B����>���?02�?��Q?��"��G�=K`ؽpY���񋾰�T=��K>�5�>1�t>s�>���>���>Ƙ�>�nW��(���Z���ٽCG?,�Q?�V>�ƿ�{����*헾���;�8{�a���>C��T���>返�U���Y��%Sb��Pr����Jþ^�b�u��$?~��=�U�=m�=j�;KH*��r�����<x�Ǽj�=���:�<��T����1⼮�V�Ǻ�<�ּ��w���˾ȴ�?)v?�V!?�yD?ي{>S�6>����y�>{Q=���>� �>gl>򞏾x�s�T:;�-���fž�����f�9����J\>+<=���9>a;�>W}�=��e<K�>�v�=v�»DVϽK=�";>�2>]52>�d>¤b>'�>�"u?�l��/���t�t4Ҿ�a�>���>�}�=#Z����?#�=J���aR����	rn?T�?޿�?��>ٮj�
�>"о�꺽dd~;��'�L��>�>���կ�>W��=Pr�S���V�l�e�?7m@�%Z?�ք��亿G��=�^8>�>��R���1��^���b�	�Y��o!?�;��h̾��>�<�=�߾,Vƾ��3= 8>�e=�O��D\���=?{���;=��k=�щ>l�D>�~�=��%*�=�eH=��=�:P>���3s4�և'�6=�*�=�fb>�5&>�R?:<�>��>N`?[?PC�=B�˾���JY���j�~��>��.:�����>�K?4�>?��W?��>6u?��F�>��>�?#��׉�l+�I@�`�>m=�?걧?rO�>(����H��Ѿz�_��ay�9�?^�1?�/.?���>}��Pڿ%�,����������ѼH>������<��=>P�̛�;r�>�a>{p�>PQF>OR<���>x������>(\=Pg�<�=$���B�<�ܼ�I=���b~�=+m�=�^��[�R<ct��!=�<=R���xY��=<���=���>}(>r��>\~�=���56>e����rM�p�d=n���{C� e^���y��T/�o��[28>�F>uɍ�g둿2�?�1�>��M>�?os?Q�C>z���a޾�W���h�(Ct�מ=5��=��\��lD��Sb���F��Ҿ���>`�>��>��l>c,�_"?���w=A�#a5�J�>z��|���&��8q��?������xi��=պh�D?UF����=]"~?��I?��?ȍ�>����ؾJ60>1I����=��M)q�;g����?	'?Ӗ�>����D��[���6<(�o>�z�=�=�C���DY���=����>�Cb��h��R�
�w�Y����F�x���Ϳ>��G?64�?�:�y���q���^V���?�NB?��>MB�>!�?���aQ�v!�YȽ�d~?d��?���?�S.>��=1G��D�>��?u�?v��?�r?G�9��K�>��o;�� >7ф���=�>]�=���=��?�?�)
?`g��<��6���߄\��0=�\�=\�>�w�>��q>�\�=��U=,�=��\>��>X�>.f>�#�>�Ȉ>c���侾bW?	>'=���>E�2?�Ȟ>�uW=CP$��i-�G�Y��ho�mO0����!M�������Խ�ǔ=�ͱ���>3�ʿ͇{?��>ˈþon,?4l�R�"�2�>`�1>'��<ߊ�>&^>��>>��>E��>�Yj>�X�>�>"FӾ�>��� d!�B,C�O�R���Ѿw}z>f���k&�ʠ�\|���BI�yn���g��j�i.��p<=����<H�?m���,�k�G�)�&���Փ?�Y�>*6?�ٌ����(�>P��>�ō>CJ��珕�=ȍ�gg�[�?5��?P��>��s>m�e?��?ҽ ����I��\x�&L���w��]�����]�v�$��|���!P?�]?�JC?U�j��M�>�^?[�T��ؽ땼>C�!�T�ъ5� ��>�"\�@��tֵ���=�w�>
A�?�)�?��? ֪��"�>� {?�10?�r?� 7?��*?�盽�_D?ZA�>*L�>z-?�F?��!?��>��a=���=���=u@$=�LȽ��������ɉ��q�<j�>��~�b��<�Ew� �>o@��iw���I���=�(�=��Y=�D%>�9�=���>��V?X��>��><�<?�Y����9��̾�R?Yz*��:�)j���o���߾Bq$>��e?�ͫ?+N?��>
A�}D9���>C��>�*1>V�f>^��>��潡�C���==m	$>�W">��C=�w���cm��^�K���$��<�>>�'?3�o>��ս�O�<p��x���[�� о�_�!��"n5�'���I�&��>�A?�a7?ׄ�=��������DX��;?A�H?Y?�x?�d�>�}M������q��Z��X:�>�<�d4��N��4Ø�&G�z��=�s�=t��.a����>�f+��T7�vo��-��#�Q�򓍾M3(�4<A>�=��l(�3Z6����>�y��S$��+C�.��GG��x!Z?��=Ѩ����a�����"����>$��>�*>3�
���+��Q|���>�n�>}��=�$�>���Ng=� ?��{t>�I?p�?�:�?)�I�JFm��1���T��fe�T%U?rX�>��?Qk=��9�����1��=���>W�>�?3�O�>�/6��Kx����<�[b>9��>	٨>L�?��X?��>��?�+�>
'
?n�?)f�w[��('?�#y?Ri�=-d*�V�n��,��K����>6t?�zr��7�>�9?*�?�0?�(?k)?°V>w��i1�4�>0�d>8~Q������>> >n?'��>�c\?R�Q?��Q>�jI��������8n>��>�E?��"?¸�>)י>3B>cq��W>�D>m+�?N��?d_v?��v<9?�>AN.>a�=nx�=�4�>2�7?�R?���?+�s?�\)?$�=�l�]'�=ƶ5=Un=�m:<Z��<���怢�rWz=� =k��<��?;(���[��G��֮���A#���S����>B�r>�}��E�9>�[����Hm2>'m3�3Œ�r=���t8���=�X|>�*�>��>��O"�=ps�>�>�)�|&?��?�]?L;�<Sb���ؾ�MM�cյ>�>?0��=^�k�*���ir��}�="�l?��]?��2�67���b? �]?�+�Z"=���þ�~b�t����O?9�
?�H�\?�>�!?a�q?�|�>�Uf���m��眿Sb���j��\�=|R�>%L�e��'�>�7?�k�>�6c>�T�=20۾n�w��c���?;��?��?p��?�3*>�n�5!�@�
�Hj��\?��>@���nJ!?��a��AྎU���o��o���o�Ѿ!ţ�񤮾�g��_���8���V�=��$?�w?�xk?X?:��f�T�%_��bw�Q[]��� �ė� �H�Z#K�O=�Z�m�W?��\ ��G��N6<�^��:8����? �"?�DE�.�>=RI�a�پ�:���2 >��q8���/>m�=.�	=�v�䩆��M��ŭ���?�p�>���>zjB?x�C���:�6PI�"QX�G^��>۸�>���>���>KC�_1Y�u���A���c��䑽z�t>�c?��K?��o?6a����1������� � �9�? ����F>Kx>'R�>�,X������%��>�J2q�L��a܏�����3�=BV1?�L|>g/�>q֗?��?C&	����'�r�J1�3�<��>�@g?��>�h�>N>Խ֌!���>�(k?ɇ�>���>�.���M ���v�c
��P|�>���>���>1`>`[7�0j[���������*;�զ�=�Zf?�JV����>��P?C!�;0_;�J�>�V<%�Z���)���=D?0˺=��5>�
ɾ����Az�����)?1�?���1+��}>�"?c��>�N�>p,�?ԛ>�2þ/� ;}?�#^?q�H?A?+�>?�= 1���ǽ�'��=��>�[>ۊr=���=���O�Y��p ���8=]�=�Dܼw����9<��Ѽ�FJ<�o�<�e4>!eԿ#M�E���6���o���Fξ�@���f�a8������о��վ2��M\��"�V���	<���낾MHO����?��?�����1̾t����^L�}�!�N��>�r����`<�`���V�J��NTW�,���@5�>�o���n�]i~�U�(?N>��ȿ�u���$޾:u?�,!?��z?��
��#�*�7�\�>��<�t���㾚��ο3>��Đ\?���>�Aﾖ��8��>���>�O>��u>|`������P��<�?
:,?� �>�q�\ȿ���{��<q�?�@�B?$"�b�ľ/Sn�߭�>�?}�>P���"1�0d�����>O��?��z?��l=V�U��=��c?w����F���d<���=��f=ڲ��2�۽��>!ܠ>���i�^I��6=��1>�Z'�����MT�_"t=12:>��ؽ��ݽVՄ?${\�]f�ģ/��T��U>�T?C-�>A�=Z�,?�6H�9}Ͽ��\�*a?.1�?=��?��(?pۿ�Eך>��ܾщM?_D6?���>ed&�j�t����=�5����N��I%V�\��=4��>��>��,���D�O��*��n��=U���ҿz �5��ح<�;v<�뛼��	6e�����I٬��s��Wӽpy=��=�^>AD�>��>A�n>�wR?u�r?L�>�M�=j�����S�d�Ѿ;ꖼ�V>�Km ���a�}zǽ������ܾ/�	��%
�+H���ľR�:�P��=�P��ڏ��S&��iZ�vYL��S$?��>�¾��L�����7Ѿ�Ğ��W��m��1SӾn�0�޸n�à?��F?�煿�[��A����z��nR?��I���`����=��<���=QU�>�p�=�{ﾜC4��V��`%?^�?�Ⱦ��-���k>�=�w���_3?��>R���Ey>��$?�W�fǬ���`>U�>���>���>h�c>�,⾆م��]7?/2d?އ=�Ⱦ�TS>�⼾m�
<����U;  `�&��&>��)>%6-��q�=}$L>��>�mW?�ߋ>�P)�?W�A^���n2�V"-=��v?�<?Az�>�Lk?r�B?��<���>~R�[P	�`�W=n�W?K�i?��>3%o���ξ�<���7?��e?K�E>Ԕm���澮�-��7��?}5k?Ig?Ct˼�L|�Q���k����5?��v?s^�vs�����;�V�k=�>�[�>���>��9��k�>�>?�#��G�� ���vY4�$Þ?��@���?I�;<' �R��=�;?m\�>�O��>ƾ�z������l�q=�"�>����ev����R,�e�8?ܠ�?���>���������=}�����?}̅?����Ec����	Hj��,�e�;�K�=i1�V<�Ǿ�E5�F�˾���g{��r��.�>��@��w��>���3xݿ,hҿ�����h޾�?���?���>�ީ�  ��-e��Fg�d[:�F�A�+w����>�>ڌ�L�����y�/�8��CH��n�>Zm3��Dy>�*��C��G���ʙ���>�e�>���>+�^-���o�?�i��/�˿%͞�_��}�]?]��?��?ʨ?h�U<�L��!c�!�ɼ�]I?.�o?�|]?��q�5E�/�j?�_��GU`���4�qHE�FU>�"3?B�>ʓ-�;�|=n>���>�h>�#/�5�Ŀ=ٶ�����C��?Չ�?�o�S��>K��?�s+?�h��7��c\����*�6�*��<A?_2>�����!�E0=��Ғ���
?�}0?F{�.�l�_?)�a�n�p���-�t�ƽ�ۡ>\�0�e\�zI�����yXe���e@y����?V^�?Q�?V��� #�<6%?�>`����8ǾV	�<���>�(�>p*N>2H_���u>h���:��h	>���?�~�?Jj?��������lV>	�}?���>��?JA>�	?��
>�$ξ��<�>��=�2�?��S?�/�>G�=�(�6c)�rC�u`;�}d��u6��>��c?��7?c�>�؞�\�_��
��BڽN�U���<�mD�l��N陽@�>���=���=K_�,a���?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Ua~����7�[��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B�k�1=7M�>Ϝk?�s?�Po���j�B>��?!������L��f?�
@u@_�^?)��s�����V{>�K�	>��:���>�r�IeM<�y�=�n������X�=�U�>*)>���>�&L>��>묆>ڈ{�k)�h�������d�v$�����B�.���� �%.�5[������f'�6�}��&�g�I6ѽ��*����=bPV?`T?rq?ל�>H"��6�$>٨��[=�<9�9�)h�=?ʈ>�e1?��I?�|)? �=ݞ��=a�Li��n��F�����>�g8>x��>���>6ި>͇��^B>�L8>�r�><��=Dma=X!��Y�<hoK>/��>��>��>H��>8Q+=Z*���;�������`�/���#�?*u<�[�V�������߾,0�d�=�c1?�>�䚿v?Ŀ�㬿�H?�о�o�Eoj�A�M>� ?��u?~�>��,���<���>�ܿ���������a�>�d_�F��L��>�&?�f�>�uJ>��=�Uz8�W�Q������a�>�aB?ߖ���R���j�`NK�JW¾�;>t��>07ݼNS"������z��VY���==�:?�k?*y��C���u�E�������$>㵀>׺�=���=�p>�V�QD��T<Z��]�=�!>�%x>	?��;>A��=t<�>B�������h�>�ڃ>.>fk5?��-?�<y>5,����گ�>�g�>��>��>s�x��w
>�e�>��>�=>t�=P{���:�Вu>��?����'D�Ò��������=c��=�7)� &��>�~?���(䈿�� e���lD?U+?v �=��F<��"�D ���H��F�?q�@m�?��	��V�>�?�@�?��F��=}�>
׫>�ξ�L��?��Ž7Ǣ�ǔ	�')#�iS�?��?��/�Yʋ�;l��6>�^%?��ӾPh�>{x��Z�������u�w�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?��C>@�?k|w?"D�>��b���0�ӽ��pM��o�/=�%!��ʝ>��>�U���E����0���#h����n�C>��-=���>��ʽf=ľc��=� g�ƪ��qo���>_�n>2`>T"�>f�?���>�>��= �<�^ �������K?{��?����2n��3�<���=
�^��%?_C4?�0[���Ͼۨ>!�\?���? [?\j�>8���=��翿{�����<A�K>�1�>�E�>���^IK>h�Ծ�2D��n�>Zȗ>na��I?ھ(-���F���?�>d!?ؒ�>~Ѯ=8E ?m�#?!�n>���>~�D�[��LF�/�>��>͐?'D�?�@?�����4����蠿?�Y�-K>�Sw?ƻ?��>P쏿�Ν�W�t��5�����.��?YZf?�۽�"?O��?z�<?$�A?�ib>���~	Ҿz佽���>s�'?���ǔ;�=�0����*�?���>R��>���;�Ž���Y�����	?%�H?S.?��龁�g�+˾M�=8�ӼHm��h=��;<=">A�>`x~���=�6">�=d|����7���3�Ft�=��V>|=�=J�1�����:,?�oF��Ճ���=�r�0{D���>a[L>���_�^?�U=���{�
���x��R�T���?���?�k�?���h��"=?��?�?/�><���{޾���OMw�
�x�w��>���>��l�� �r�������]F����Žf���p��>o�>�h?p�>�j=f�>r�<"%��X�Ƃ�MXf�����h�.��/6���޾�kz�������Պ����>A?߽�v�>�w�>ﱧ>�p�>�I�>�6�D�>�L�=��>���>f�>�p�=��>J��~~/��PR?���8�'����&���Q,B?.ud?gK�>�Lh��l���n?���?l�?B�v>�xh�%2+�bd?�&�>���/j
?Y�:=�S�n-�<Ug������=������>p�ֽ�:�s M�+df��e
?�#?!���k̾��ֽTs����q=�[�?��(? �)���Q�w�o�`�W�S��=��Yf��+����$�"�p�aُ��S���	���s(�&=H�*?o�?=��������y�j��<?��'f>>��>s~�>���>J>��	��1�x�]���&�*��
��>�={?҆>$�K?F�:?�Y?�/L? u^>e�>8Y��`��>�q�'(�>
��>/0?�?v~1?^�?�"?6��>�K�#���ɍǾ�;?�s?�J?�S�>�?������Y�j�-��N��8����=c�=��1��s���-�;W0>�W?s��8�p�����j>z�7?Lr�> ��>?-�����Me�<�
�>J�
?�5�>  ��ar�G�#�>N��?90��>=8�)>+a�=�p��!0ͺ{d�=C���i�=����Ɔ;��<I#�={V�=��k��m����:뇇;�<�t�>b�?"��>E�>�?��m� �G�� f�=Y>S>>�Dپ�}���$����g��]y>rw�?�z�?�f=>�=��=|��NT������������<I�?J#?tWT?%��?��=?�i#?�>�*�xM���^�����<�?ĭE?#��=�]!��_��V����M:�.�(?=�"?��1��'�<̭龇���N�P>
6>+�d`��������N5^;�;��y�g��?�Y�?6=��V�1��E��B����?�v�>�e??��>;B�����ʾp�=��?dYs?%�>[8J?FnW?"�^?�!A>�PN�ޥ��ǜ�_bB=Hx>�AI?�	�?=�?`��?}Y�>.>��2��^���rܻ�	���t��Q�;���=i۾=c��>9n�>�C�#��q�;g�O�TI6��2>P��>�}�>�?�N�>=���G?l��>�ƾ�J3�Qा�;����<�^nu?���?�+?�=G��mAE�F����e�>�s�?:��?*?7�T��R�=�ZӼ,�����p�)�>��>`h�>�A�=�F=+>���>�H�>l������7���H��~?]F?W�=�ƿ�q�]�p��ӗ��wg<�ג�{�d�:����Z�1��=C���Շ��թ�b�[�5���'���Nϵ������{����>���=v��=Ͻ�=, �<Aȼ -�<��J=24�<B=�bp���k<NG9�ɵһ�舽L�.6\<��I=�����0ɾ�/~?wHK?��/?�B?�Of>��>�8D��֐>�C���?�8b>E�W��/���j/��˩�ס����Ҿ��پE�`�S&���Q>'�t��->FT3>f|�=	b<b�=U9R=��=5�1���G=2��=k��=p��=�M�=T	>֣�=�6w?X�������4Q��Z罥�:?�8�>f{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=J����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>zê>�=0>�5�|�K�"�U����=R>\��s%?7�X�2�����0>�G�>�������޽�)�>�aq>�+Ծ��F��5=WM��r�� �U>
�>��t>�f=]f��yB>۹E�s&�+m�<k�u��JG�g�=�b콬G�=�;I>,e>��>�?��(?_?9(�>�s̾3���n��$�&>�L�=O�?�>�6|>�ø>��?�3A?ܸ<?�;�>7^{�m�>9,�>�F�v@]��g꾐���Q3=i�?��U?�Ox>\� =|}^����`��p����)?�g'?�"?3��>�����%�p�,���O<�;��=":q�;�B�9�<��R�Ɍ�O?�=җ�>�ʱ>�٭>Rz>L~>�z�>�>��>{�=�+�sb ����=e�&���p=�>�=���<�͚�k�c=�q<���
5V���O�z�Z=�_=X�7�>��>��i=B��>~�=N����=�_���.��]O>5`������F���{�a4&��B��o%<|S;>99�;!�����?.S>�8r>�>�?�,h?/^�>�^��C����о�{���+L����=�B��d^��A�+mc��3徝��>�t�>���>���>��(��-=���1=�߾��'�C��>���k�������n�飡�B���m��j?9T�D?â���
>t?�8G?�m�?�P�>�u��ɾ�>-O����X����U���`����?��?Р�>�g���B�DF̾	����>�<I�]�O�9�t�0����ͷ�D��>����о�"3�Lh��������B�QIr�0�>ϳO?�?>b�X��JVO�������o?�|g?��>�K?,??����{�p��Vn�=n�n?��?�:�?�>	ƽ��F�
P�>��>�-�?��?��o?X������>��;�ʽ�����|�1�Z�>�>��P;C?>%?	.!?�e��-z��ž(䧾������Ƽ�U>.�>��>Zr^>�=���p<r�Z>l>�,>��=歗>Ɖn>|���
��7~#?u�>��c>1]?:��>��>>��Ӊ�=�j����x�	(߽;��<�������H,/�t^��>M�h��>��[�?��>#M�p�?�+#�*�>�{B=����K�>{��>��>s��> ��>�>m\�>X��=wFӾ�>	���d!��,C�<�R�.�Ѿ�}z>�����&���xy���BI��n���g��j�[.��a<=�F˽<H�?������k���)�Y����?J\�>6? ی�T����>���>yǍ>lJ��I���Oȍ��g�z�?��?�6c>n�>-�W?h�?�R1���2��tZ�6�u�0A��e��`�K֍����
����6�_?�x?�qA?ԕ<��y>$��?N�%�TÏ�89�>�#/��;��k;=x@�>���7*a�e�Ӿl�þu����F>��o?�'�?3o?�U�K%n�p%'>ȯ:?φ1?cPt?��1?�;?K����$?Ga3>�=?�q?�95?��.?��
?Y�1>h_�=S����Q(=�(���ߊ��Qѽ�zʽO��I4=��{=�L��e
<��=�1�<=���ټp;O���ǩ< �8=ۦ�=���=$:^>FL?O�	?sÜ>�@?���u�&�u��" ?#�}�0ˇ�P>�3񐾡c��b�>�|Z?�?�b?�W�>9ٗ�H��D>�E�=�%�>`B}>���>/Р���y�ws�=�7>jd>O6��ڭ=��ս��<�玂�V=��<�+ ?V�i>`a���';>i襾�7��B>>X(b�j����p����=���%��H�Hó>�SF?�'?|�<��׾d����f�1>,?�'4?�EL?���?���=��޵8���A�p�)�'q~>_=P���Ϡ�|M����<�u�ƻ��K>2u��b���"Ѝ>��/�
�Z�t���5�kd�)��<^��\�=��Ҿ�K۾ �I���=^B >:���w�e���U��43I?WK�=��ž��_�|㯾)�>
�~>=6�>��=����f�3�gĹ�嵰=���>�(>�_�=���"27�
�-��>v�=?| i?ڍp?6�����k�� :�����n־�r�=h�0?".�>�w?�^�=Pܼ6���l��7/J���9�Xf�>��?�<��qL��J�����L�#�|i#>E��>���>��$?p�B?H�?��Y?���>�? �>Xd
�U`��aT'?9U�?TR<�w �����T�g�H�KG?-MZ>[e �nB�>Z�-?#?{�>��[?:��>P)	>�!þ�+��إ>v��>�]��������=�;=?�ֳ>�K?-�z?|��>�yN�)ؾ�R׾���=��=�f?�<?�A�>���>���>In��,�Q>K�>��v?䁈?h�S?��-�Y5?��?>!�>���=֢+>�?��>�t>?M�?�dQ?�,�>=��<�ꐽ�b��GE˽\{<���=Q�=���<��Z��K�<꫞<z-O=+��<���l�ۭc�m���BAT��6��P�>�t>�敾m�0>��ľ�<��l�@>�U��?Z������K:���=օ�>��?m��>�y#��ڒ=���>�1�>��9H(?l�?f�?�0!;ĉb�	�ھ��K�!!�>�B?�=��l�Rx����u��h=�m?J�^?F�W�Q8����b?0�]?ud�S=���þK�b�"z龐�O?2�
?�G�O�>��~?�q?��>��e�s7n����'Fb���j�)϶=pj�>rP���d�.9�>�7?IQ�>x�b>�E�=y۾��w��m���?�?��?���?� *>?�n��2࿡S��"Z����]?�D�>�Ħ�̮"?����4tϾ�>��s폾o���ڪ��Z�� F��~���.�#�L���[�սg�=�v?#s?)q?��_?�����c�^�vV��XV���a�_}E��:E�w�C�� n�������ؘ��G=yYD��f/�6v�?�&? %r�,��>���ߣ�Д����=�
��*�0���=�Y��K!>�+X=����vHt�`|վ�+?l��>m<�>o�8?+�O�;�I���9���X��{���>7��>�r�>���>�ٺ<���=e���첾a|2�d锽�w>z�b?II?`�o?G��+�0�
b���S �(14��b��ڑA>� >���>q�`��P� '��>�H$s��?�����Su��?�=��1?�v�>��>���?D�?��	��'����w�712��!�<&��>�Eg?���>�x�>��սF�3��>6�l?�j�>xi�>򏌾mS!�}�{�q�ɽ
��>>���>��o>,�,��3\�J_���~��x9� ��=7qh?����U�`�$��>y�Q?�8�:pN<<��>ar���!�A���(�x>�?!{�=�f;>Q3ži��{��鉾ub$?ܠ?������'�?׌>��!?�j�>���>�9�?�>��о�����?ؖ[?
H?R�<?���>*W=�m��
Bн��=���=Yc�>�f>��2=1G�=g�"��}c��z-�I�C=�$�=��V�f������<���㖧;���<�->G�ſk(O�X��,���m�)6뾑ɭ���$<ֺ���qn�K���y�8����瘄�Q���¡��2�O�?�1Q ��@�?q��?򑱽���F}���X;������>�+��{�>��˼L���	
���ҾT���+��!�wBT���k�k�'?nˑ���ǿ ���qIܾj ?�M ?��y?����"���8��L >���<���o�����H�οZʚ���^?#��>��Tڣ����>�n�>�eX>�Xq>�%��! ���]�<�?}u-?L��>P�r�Đɿ�����<���?��@��@?�$��*&�=4��>`?�J>�Z7�U��$E���)�>�G�?�L�?�[=��V�c����d?��<�H�w&�h��=Co�=Bd=�&��MN>o�>��fD��Y��0>��>�A�Q<���V�9��<�U>3���Ľ�ք?|\��f���/�U��(O>��T?_7�>��=��,?�4H�e~Ͽ��\��.a?#0�?���?��(?뿾D��>	�ܾ��M? E6?f��>�l&���t����=!�ἵ;��ް��+V�@��=��>-l>F�,�����O�����2�=�^����ƿP;����=k� <�������@��������G;�l�ȽZ��=����wn�>�\t>��b>4�>tk_?{�^?���>E�]>�j��⏾�ܺ���<�������>Ũ�8��1ݾ���v�����	�Ih�"(�������/����=��O�DE���+��O�4�V�ii(?='Q>�%Ⱦ�6�����f崾�چ�\;�iq���p۾R�0��Co����?��,?xb����B�2r��v��^���Y?
i��^�#*����=�>���dQ=9!�>@3>[ ���K�o�O��6?ڝ<?Ǌƾ_̖��J6>��;�ɻ�c3?��n>�>C͖>�/?<H��!�U���4>��>MW�>5��>��d>���uӽS[*?��U?[H�;��x����=-L���Q��v[=�!�>��2����=�L�>��=�Z��GY6�폓=�]S=w!W?���>��)�,��Z���_���==�x?�g?��>p�k?�C?��<�X����S���S�w=��W?�i?��>�Q����ϾD`��~�5?��e?�[N>2h����1�.�WU��$?��n?�<?Ӗ���l}�;������t6?��v?gr^�6s�����!�V�1>�>M\�>���>"�9�)k�>�>?�#��G�������Y4��?u�@|��?3�;<�!�8��=N;?w[�>1�O�[>ƾ�x��&����q=L#�>ތ���ev�����P,��8?̠�?��>	������lk>֍��.U�?6j�?�;��I�X�!���Xy�	X��<:�=�����<�d���70����{`�����-���7ކ>��@��e�>q9&���俦�οa8���E�ֽG�?�T�>i��̾��瑃��\a���/�A�1�o�*����>���>.�+��7 �,ⅿ������ ;�>PZ>Š/>>c���$Ѿ&gF�	�(>X�:>(?���=f�F���r{�?��S��Z%_��о��+?]ˉ?���?��/?�y~���Ǿ��3��X@��):?��A?x��?Oޞ��m�����+�j?�_��vU`�Ύ4��HE��U>�"3?�B�>I�-�=�|='>x��>�g>�#/�b�Ŀ�ٶ�����=��?Ή�?�o�=��>i��?�s+?di�8��\����*��*��<A?�2>z���V�!�I0=�9Ғ���
?<~0?�z�_.�i�_?-�a�j�p���-��ƽ�ۡ>j�0�Ie\��O��H��zXe����@y����?J^�?Y�?��#�!6%?�>q����8Ǿ��<T��>�(�>X*N>�I_���u>b���:�jh	>���?�~�??j?�������<V>�}?�-�>B�?}��=@��>���=➰��	8��">���=}�<�W�?`�M?F�>$��=�7��%/��F��Q�k��.�C�~χ>�b?�tL?��c>�B��m�2��� ��aʽ��1�?�c�@�>�*��_ݽNf5>؉<>�>=dD�;OҾ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?!�lP�� a~�J��4�6����=��7?-0�8�z>K��>��=4ov�˻��)�s�ո�>�B�?�{�?���>��l?o�o���B���1=�L�>˜k?t?�o���n�B>��?������iL�f?��
@Ou@��^?�� !ֿ�����̾ѧ˾,��=ZC>�PX>�+��)>�6>�|��E���(>��>�>�w>��P>\��>bB�>B���@]��򘿙��VK�i�"�A
��<������1zo��"�l��=�k�sV<���sv����J�lŽ�����x�=� U?!R?��o?T�>�,z�P�%>����j
=�q'�H3�=M��>5�1?�<K?��+?�"�=6;����d�C���������8�>��G>���>�?�>)q�>:b��6�G>�&=>���>��>8�/=���yo=�O>���>�;�>�l�> ��>�I�;�?п�����b�(3�<©����?����ϋ�Y�[����������>��C?�7?��:_�@¾�ƺJ?�B�Ga��Ty �aD>��>�m�?Ɗ6>��#�?�>Uֽ=�쟾ehz�oO>���=Z@��ȿ��(!>l
�>�M�>0"\>68����hJ�$�=��>�y7?�}��+����i�2H�v��Vj�=n�?b%<��1�Q��a_����E������O?Sf�>_9�Ib��$GR������+>�,%>9��=y��=&�>ǣ=�Os>;������C�$>7�=�?��x>��=)��>V��|5��oA�>1�>�ɼ�)?�)G?�~�=E�3=rpN���h����>�G�>�k�>B�;@�X����=t)�>�lt>w�=�c=��\��:U��8)>i/�� ~�..�s�j=!�
��.>t�'<���٭����J>�~?���)䈿��$e���lD?U+?x �=��F<��"�D ���H��E�?r�@m�?��	��V�;�?�@�?��C��=}�>׫>�ξ�L��?��Ž;Ǣ�Ô	�<)#�gS�?��?��/�Yʋ�@l�6>�^%?��ӾPh�>{x��Z�������u�x�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?raB>��?�]t?���>o���*�Cϳ�=���{�K=f<�k�>�%>L����iD�]6�������f��;��FR>l�5=dp�>ۥ�IHǾ@`�=nw�S����ʁ�k��>N4q>�V>2�>9�?�b�>cb�>D2N=�䏽�i|�㺟�g�K?h��?���W2n�zH�<���=?�^��&?tI4?Յ[�z�Ͼ�Ԩ>��\??[?�c�>t��O>��2迿�}��Х�<��K>�3�>�G�>�%��LFK>��Ծ$5D�.p�>З>j���?ھ�,��=D��MB�>Me!?�>�Ю=<� ?�#?��j>�0�>�`E�=:����E�r��>��>J?%�~?��?�ȹ� Z3����䡿��[��1N>��x?�T?DΕ>/���Á��^QE��uI�����?wog?(%��?�2�?�??K�A?(f>`{���׾������>��"?4��JF@�l�$����	?B'?w'�>���:u˽�W&����e�����?d[?($?#� �.a_�𲾾5��<o3M�������}�k�!>G">ol����=E�>��=�;g�Y>�Ǆ.<[|�=r��>���=^2�O����<,?ȤG�uڃ���=��r��wD�|�>JL>�����^?Fl=��{����ax��|	U�� �?Ơ�?Kk�?6	���h�"$=?��?Y	?�"�>�J���~޾֔�QPw�?}x�#w�y�>��>��l�C�����ҙ��lF����Ž�%r��_�>��>BD/?�ο>&{�=x�?��#�hs⾟���Xd�� �S�F�� ����x�Ӿ;���k`�]����y�A��>����׏>>��>|��>��>���>S�2Y>�U�=��>4��>�
�>�d�>ڏ�=Oj��"w��KR?�����'��辘���<3B? rd?z1�>�i�2������;�?~��?"s�?O=v>�~h��,+�(n?6>�>�� q
? Y:=D��5�<�U����A4����>�D׽� :�]M��mf��j
?�/?����̾�<׽�[��pq=P[�?�)?*�,cR�^o�!�X��S�f���e�A;��S�#��rp�x�����;1���(���%=9*?��?'m�$�NP��zk�ix?���b>���> ߗ>�5�>�M>�����0�ץ^��&�^���S��>�B{?W��>�_X?�O?�U?xD?�t`>7>�6��b[�>8�=x��>�Q�>��?n�5?�:/?�|�>wY?'��>�b�<o��>l��2,??į>?3� ?g�>��f��-�=���}"Q��Vn��φ;;̈́=n;=��m����<�=���>B0?�>�~a8�����\"j>��6?j�>5��>A9����v��y<���>��?�>/u����m�6����>]�?m���=}U'>01�=Ǵ��KFq;���=?��b�=U�l��!�14]<n��=��=0P/�P�<;6��;��;�6�<T^�>/�?�>��>���Ԁ �Ē�T��=�rY>�S>*f>�xپ����!���g��My>Vy�?'{�?�xh=-��=��=Fk���Z��'���潾m��<�?�`#?�`T?R��?��=?\#?��>���;���X��W��K�?�L?4��<g�:����ҽ���[D�t/?j��>��g���=�#=�x2��,D=��=V౾Z,|� j����j��Ra�.A��Y��8��?���?�q��a�~�Ԭ'�2����|�6�q?l>�"?S�?�m���`�L�3�	�k�� ?�Џ?���>S�B?GDh?��|?���=�=c�ʇw�:6�������"8>Vbv?\��?|�?��*?\��=AM�>�ٽ�?y�����D��{���Ǿ��뽢�Y>{��>V�>D^�>�x�� ��������a��=��!>���> GW>QJ ?�Y�>N����H?��>�¾V���M���|�GD2���x?ˋ?�E+?��m<�B���G�B���d��>�K�?z\�?ё%?�F���=��Լ
ɵ���y�AC�>ҵ�>{"�>Ά=V�=_�>/@�>>��>, $����:�-f��?2�A?HF�=�ƿ��q��q��З��co<.���H�d����Z���=h����a�2k���bZ� p���!��x����=��d�z�2��>��=��=\m�=��<Egʼ(�<�yI=��<�!=�q�@cl<b�;����ѥ����"\O<��H=&��ɾ�t}?�1I?��,?��C?aYv>��>�A+�%X�>d���?��]>ʮ(�e��E!8�,H��9�����վ$�׾W�a������d>�@T��>�U4>3�=<'7�=��z=9�=Z���=r;�=��=5ݦ=X��=Gx>�O>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>
�|>��j>;JO�SB/�h>�3.��1�O�5?V8�:ܚ�-j>
t>�� ������;=L@>>��'>��k�<���=��b��T�<9%V<4�s>��h>�
>�ڽLJ�=��{=uZ�=��N>;n�Rh��6���#�=�d1>~ER>�@>>��>(?��3?�_? �>9�L�S�ʾ�}���Lp>>��=>+�>�ȶ=�<>%��>�/?��.?�VJ?.+�>��=��>�<�>-4���s���ھ�����b=`Q�?���?|ޥ>�!D��~Y��3(��6I�z5���?~�6?0?���>D
���G-�4�7�a�<�(�=;ʟ��ӕ��5>lB�Eb2���ȼ�B>�?q@>͡>�x�>���>�B�>@��>���=7�=|\>c��=�K��:���>��ؽ��	�P��<���=x|����� X�!=T���^��Ln���=Ԟ�>P>��>=�w=n�����/>�����H����=�آ���>�Wh��.���*��5U��#>�<>���������@?�0X>�E>���?k�y?aYO>H;��_�Pѝ��[X��t��Z�=��>�P�Qc2� W�M���ž���>[�+>ғ=���>��D�M�|�������� �p*#?���6��=w0#�U���%Vf��i���N���K4��/�>�タ�i�>��G?�v_?���?�@#?��d=�si��O>�SȾ1�T>���2��64�{��>�� ?S?��þ�PE�dG̾� ����>ZI��P�����_�0����sӷ����>�᪾��о3�8d����1�B�+(r���>%�O?A�?J�a��H��rO���%����_?0dg?��>�W?+S?�c���I�b�����=��n?��?�+�?
�
>�L��Q�<~�?NE�>롦?zu�?��@?��^��j'?�-�����๾� ˾`eA>*av����γ<?��;?�uC?㱽�uӾG����齾�,���Y*�=�z>	}�>�#>[�,<�c���Ƽ>E3>�
<>���>Ʀ'>�C>
j8>=��1
�@(?i�=g��>��-?���>Vzf=<"��jSD=d��!�����b��������e�<��a����=g�ٚ�>Tſ��?��i>�*��\?�E�a��;47>\$>�c�����>�G[>��>U��>���>>B��>d�>�FӾX>����d!��,C�X�R�~�Ѿz}z>�����	&����w���BI��n��ng��j�P.��]<=�ʽ<$H�?����
�k��)�����X�?�[�>�6?�ڌ������>���>�Ǎ>�J��g���Oȍ��gᾙ�?<��?��b>n��>��W?>b?>^/��J1�$Z�Ru���@�+�d�_�`����������
�S���_?�y?�A?�[�<�ky>�[�?c@&��ݐ��>�u.��w:�� ?=gb�>�0��zc�HLԾ��ľ�H���D>q�o?e"�?(�?`�U�n�*8'>!;?!H1?��t?��1?[5;?�A��Q%? �3>?) ?A_4?�K/?��
?�&1>Vf�=���� /=o���fC��4�ν��ʽ;$���w.=�ey=�=\:�.)<@n=�Ӡ<-��߼$�$;�����<��<=q��=���=��>"�S?f��>��4>x�D?V��O�'���I?t>zU��7��w�/ھ�n�=�BQ?I��?��`?7*�>�1N��v����(>��>\�A>�) >�=y>���-�=��=F�>ߺ>y��=�94={���]�DN��գD�G��=���>�z>�Qu��,>l��[z���p> �Q�t���zz\���F�S�1� �q��>
�M?�/?�ރ=ղ�!}���Qd��n(?l�<?3_M?�#}?�j�=c�ݾ��<��=L�H��2�>m�<�c�����.���w9�C0i9z�w>�ܝ�����*n>-@�4�־t.k�1�J�M��x��=��/�T=��}KԾo|r���=Oc>QG��2>#��ϕ�Q����DF?S�z=F�����V�"赾�>m��>oh�>0JS���R���@������Ȫ=��>��&>d��_�GHI��?�@��>{�G?�u_?���?P@2�'p��]Ry�c����v��>)?�>�!#?��=K9��ﾡ�<�)JP��K�{��>u�>G.L��<R�⮆�@\�;����;>!�>��<�D8?�S?t�> �#?5��>�%?#y>D�d=YG��j�/?���?�n�=U� �0�J���3��O�a7?ml
?s� �QX�>��!?�g7?��>�S?��?N5�=�C �&KL�b��>�|t>��S�&+��;�.>-G?���>�yH?��\?<�g>?2�ӝ��lE�AS6>dAW>�U.?o?��?�8�>>�>�����$>,��>l{q?n~?F�^?F�G=�`?�+>���>��?<�q�=�d?3
?�c%?Zo]?^�C?�}?��l<���ꈑ�G������<�<|=�����.=ߌ�=�C~�G%����;D�T�
�=�#����.�P�:���G<���>>������:>���k��2y>ʤ��U.���(��Σ�#�>�3]>= ?Sð>�?(�:9�=�>��>3b"��� ?�v?ju?��=�P��]־��ӽx8�>
�,? ��< �n��~����|���H=u�b?�}T?|���ɾOUe?�\?�Q߾�3�L������3�G?�)�>��)�7��>U��?�"|?޾�>x�C�]�[�V*��>Q[�%v��w�=�r�>�~���p�+Z�>8v4?��>`r>' �<��ž�Gh�k����1?N7�?�Ȳ?���?\�4>md��7ۿ{���5.��ӣ^?���>)q���=#?����2̾�0������y�XȪ��)���ϕ��U���K)�񭁾)7ݽo$�=S?h1r?ؕr?Q]_?�D���d�QV]���V���o��lgE���B��D�>xm��o�����f��yD=5�2���B�>ٸ?�4?��e�L��>����<B��J殾_+>����B%���</��5�
>n�u����V������4="?i��>�?��<?�8w�`yj�Sn+�M�e���E�_>P�>�+^>�g?)���(L"�����c�V��Zy��0�>�#_?�MG?z�i?Cs#�2	>����R'$��нU���Yu>t>K��>\,���Խ�%(�E_C�� p��������͝�-k=�$ ?g>2J�>��?E�?UH���ɾI�<��%��tļ��>�q?l��>к�>>z���"�ʰ�>��l?,��>���>߅���O!�h�{���ʽ-�>�ŭ>��>��o>��,��\�e��
���c9����=Ţh?����C�`�r˅>�R?&�:�H<]��>�[v��!����#�'�9�>z?۪=w�;>/�ž�5���{�XM��md?�?*al�!��>Ñ?&��>%�>�k�?ޞ�>k{վ�q@����>�od?�-O?H�5?VR�>�b=�G���ý@�1��=�<,8�>xQ_>�j�=v��=����gC�4�&�8Sk=J��=���v�1E�<{Q�T)`<�'��:>);ȿ��G��O����*��ѾMA����<�'��������^L���v7��iF�y#�㐈�.̊���W�/m�?�	@Fu��M5�}���نq���+�!��>�v�;���SE��G�R��Е��侬�;����n�0�x�q9v�V�'?�����ǿ󰡿�:ܾ/! ?�A ?B�y?��;�"���8�� >8D�<�-����뾛����οk�����^?���>��/�����>ۥ�>��X>�Hq>����螾U5�<��?#�-?"��>��r�0�ɿ`����¤<���?-�@#A?�y&�Q�D�C=���>Y�	?�aA>D	3�R:����?j�>X��?�j�?��_=�V�V
�-mf?�X�;�F�..�(1�=�ߥ=��=��	��I>��>���6�g߽��2>.��>�|�4���9]�-�<Wc>�tӽ�8��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=u6�󉤻{���&V�}��=[��>c�>,������O��I��U��=����
Ϳ�
(�M_�v�T��FO=ꔑ=�Q׽Iq�u�n<D=���f�����]2=v�=6<�>Kқ>���><�>$v]?΋w?���>��A=�2���o�aԾQ�=�pI���E���h��� ��Ũ�6\�w!վڑ	�ě2�6���y�����.�_>sp��8��/�B���<�>�Q�M3?���>�j��VB���$.����þѣG��`>����<%��U�l�?u�W?��R��)�L#�=�Y��56G?a�~�!����j�"�ȼ�ut�!�u>��~>W���q������44?o-?�!�� 	���M�=¢8<$R�=��?v��>}�.����>zEP?Mu��c��<�JC>��>�7�>2�>|��<Z�ƾ�����	?��A?rZ�w���?k>�ɾR�H<�B���=E�#,m��.O><�U��d0B>���g>�&W?��>��)����]������n==]�x?�?F)�>Jyk?��B?Ő�< f��W�S�*�͂w=��W?�&i?��>r���V
о[����5?V�e?��N>�`h���龦�.��S�9$?-�n?t`?�>��Ov}����!��Pj6?��v?s^�xs�����K�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?��;<��P��=�;?k\�>�O��>ƾ�z������2�q=�"�>���~ev����R,�e�8?ݠ�?���>��������8>씊��!�?F�?�mپzl[��_�ҡs��v�`B>R���˽�#">�v�����������)ܾ˯����>yO@��K��\�>�7�|.��$�� n���.���2���"?���>��=�5޽3^��Ѓ����n�:�/�ag����>C:>�{�����i�{��<;�����i�>��>��>d�R��������d�4<F(�>ޮ�>���>}����|��
��?���nοI���D����X?�,�?�l�?g�?�c
<n�t��z�����F?S�s?�2Z? !%��`^���F�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�[�_?)�a�K�p���-�{�ƽ�ۡ> �0��e\��M�����Xe����@y����?M^�?h�?ѵ�� #�h6%?�>d����8Ǿ��<���>�(�>�)N>hH_���u>����:�	i	>���?�~�?Qj?���������U>	�}?P��>�?��>x�?i�=-%�ѽ���>����L�?�?? p�>�ֈ=7:�<*D,�%II��#2��N���C�s	�>�kl?�>?U�>d鼣�����@�U��1��ߓ����J>�<V�|�{u�=��=��=����U1����?Up�7�ؿ�i��p'��54?3��>�?��o�t����;_?\z�>�6��+���%��|B�a��?�G�?>�?��׾wR̼
>#�>�I�>��Խ����[�����7>(�B?Z��D��p�o�o�>���?�@�ծ?^i��	?���P��Ja~����7����=��7?�0�*�z>���>9�=�nv�໪�`�s����>�B�?�{�?��>�l?��o�O�B�&�1=LM�>Ҝk?�s?_Ho���g�B>��?������L��f?�
@~u@b�^?$>ٿ� ��/�;�Ҽ��G>^�=�,>���q>%O)>n��ّ�;0�'>���><�X>�|j<�݃>E�>�_�>ο���^�F!��L��&*�ZG!�Bb�D��9��@^�p�쾤�������载>�O����MD���H�*{�Z�>SHT?[�T?o[j?�W�>
��$7�=��ؾ{a����/�*�=0(�>Q�,?��A?p�3?F@)=S$����[��o��3����j����>��?>���>���>Xd�>f%�<
k*>��>��g>�>�K�<�}���
��e\>�>�*�>�>�r�>ԅ>Eʿ-㹿����
D=�����?4lj��U��5�l�4j¾  e����P�>R�?�}��m�ݿ\.���~J?��׾n޺�������=a�>�dX?Ufg>X�y��&pO>ȳн����S�=I3A=h�"�����w�	�>Ɍn>B{u>��4�w�9�ES��v��?"z>��8?�>���M@��Fs�n#I��!پ(G>���>�tJ;����헿5$���td��z`=��;?і?�᯽��~�k�=p����L>��o> K =���=��T>�H���ؽ�M�5=ӫ�=Rc>�?��K>��q=�ؐ>۝�/0��n�>+$>w]>�i5?��(?��=��$w[��>!��,d>ب�>ίj>�b�=d_��I�=6��>D�m>�H�;;4��?� �СG����>d���Sd����3e�=[���G�=gG=�H����7�n�t=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾOh�>x�yZ��k����u�ܷ#=���>�8H?�V��%�O��>�dv
?�?J_�������ȿ'|v����>4�?}��?%�m��A���@�I��>E��?�gY?�pi>�g۾@`Z�ǋ�>��@?lR?��>�9�W�'���?߶?Ư�?1�N>�Q�?�v?�'�>�5�r61�l���������-޻*��>�->��؂H�L���`z���6j��`���,>�uH=o�>��y=���I�=b�>�O������zk�>�\>P+_>��>Y�>��>t�e>��=�9X�b�v�S@����P?YQ�?1Z	�>lm�t��:L�=��}��`?�?�&<%ʭ�휶>�`?�qr?��W?�>�=�NA��o]��_���N�<ţ1>Y��>x��>jL���n>baɾ,�d��Ai>0��>2�6���� 2�^�/���>}y#?�f�>J��=�� ?�%#?sOp>w�>#E�c����	G�+'�>��>$�?��|?V-?����AT1�U��'����\��;F>4
w?_O?���>�L���(������O[�i����<�?|�e?�འ�?�&�?�>?�WC?�F`>`��9�ؾe��jw~>,$?9����P>�z�'�c���O?Z� ?���>ŽŽwhĽ�6���'���뾥�?�Z?8'?ea���^��(˾�~�<����!���;`��]V(>	-(>�y��:��=}>�=,(d���O��=u�=駌>"�=�"0��Hx�=,?\�G��ڃ���=>�r�PxD���>~JL>����^?�j=���{�����x��gU�� �?���?Ak�?C��5�h��$=?�?C	?�"�>�J���}޾e�ྰOw��|x��w�9�>���>��l���6���Ù���F����Ž�Fս�[?��{>�?�
?��>��?6Q��������H�D�|���/�x`�ʏ[���2@��i�I� ��`Ǿ�_�H+C>~�ѽͳ�>��?�G>��F> �>��P=��?�H�>Z��>���>�^�>|3T>߲]>���<zI�~KR?,����'�b��>���0B?hnd?l,�>+2i�鉅�#��J�?`��?�r�?
Dv>:}h�)+��l?\7�>{���o
?��:=��+ǉ<S��.����X��ģ�>�O׽`!:�M�ixf�ni
?�.?E퍼x�̾�׽fŝ�Ķz=�q�?Av*?tS)�(�S��3p�3�X��R��X���h�៾��!� o��⏿����nY���+)���=�`*?ǰ�?�F�Sv���ڎj�>�@���_>��>$��>���>�N>�.	�~�.�cx^�B�&�pY��ps�>9z?���>BfK?��-?�n;?��@?�Y�>��>����G?��սZ�>��?�J?a4,?�i"?�|�>��K?�TY>*���c����վ��*?z^!?��9? ��>��>M�B�������.yپW�O��ڟ��p���'�> ��o>�Z�>��?S�ݮ7�hw���5m>�7?���>�k�>�4������M6�<]N�>�	?���>����`7r�C
��Y�>S(�?	�o7�<ag)>�
�=� ��2�Ѻ Y�=ͽ��b �=?f��UB�,Q�;Rռ=�Ó=��V����M�P�~��;�P�<��>CF?m�>�j>�e����K"	��5=I�3><u>%�>$�ľň�w��I�a��Lv>�%�?.b�?���=��=��=�A���\ξ\V	�&��mj@=��>�R(?��W?�(�?��;?��!?h�'>P#�K����"��"q��C?H�G?�Hr>N)�Zϡ��)����7����>���>t~P�C�6��$羞@��}>���=R�P�g�	��|���2���N�ss������?�*�?!��=�f^�@ӗ��,���ff�Al{?��O>��=�}�>�V��v�.R��:�<�� ?�`o?��>�SG?�i?��M?�p�=��U��Ƨ�<甿�N.�S(>�_?��y?���?:��?.u�>�>�=�W��O��K�����~����bU��ֻrP>7S�>��>�X�>d���兾,",=u�������u�=@$
?��>8��>T��>�h:���G?&
�>?d���m�ﰤ��]��%H7���u?�r�?Bq+?�=��F�Q���I~�>�J�?0�?*?A�S�Vj�=׹Լ�ٶ�!r�2��>�>�7�>m�=~�F=	>�Y�>���>�Y�Q��O8��YL��/?�F?���=��ſӹr��t���>d<?ő�ta��z���9Y�H�=�������!����[��(���C��!Ѳ�=���/v����>�Ҁ=� �=&{�=q#�<�k�����<�R=�I�<='=�v��@l< �7��R׻7���'S:�m<�Q=5���]��s?��>?��?�D?Ȇ�>_�?>Z(]�^��>C^߽ȴ�>?�r>��ǽK����)������v���ݮ��þ�2d�`���!� >�|e<.�>
>͡>i��=E�H>Ӱ=��<y�����;Uz=We�=P��=� �=ƎS>��9>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�K�>}��>;�3��9��D���㭽�VF�Ge?�c[�xr���>朞>ܝ��喆�?��=}�>�o�=�:���c��u�;	]���w��i�:=:6>��>Ns>VT�ԏ�=���k�=�F�>7���ȋ�=��Ͻ<k��O�>�T>�rs>o��>z?�I0?0d?��>�<n�&RϾi����l�>@�=�ӱ>_�=�@>w�>��7?-D?�K?���>h�=fʹ>���>Dt+�U�l�)㾔'��WB�<Ӕ�?cX�?_�>�9<��C��[���>���ŽE|?q1?v	?�Q�>�������5������=#ߙ�X�g=0����=7�c>R_=#bl���>eB�>���>�A�>�n�>�	?iR�>�d�>T[=�e�b
>��v�B�=?��=ΐ�=>����<a�q���t<���<��Ľ��Լ/8>Nl=�7p=�ۧ=���=���>��>L'�>��=܃��H�<>^;��8�L��g�=Ẫ���E��7e�?.�<0��@9�o�:>|V>ǆ��	��bB?�WW>�m4>_��?d�v?�A)>����Ҿ؈��$�e�s�Q��W�=c��=��?��9��zZ���I��ϾӜ�>�m�>7�D>p��>19.���>�Z~>��̾q�!�?G?.��=/��P���r��~���?��Mz��A#��?�P����d>7oR?l�?�٫?�? ��>Г ��G>B^��w۽��+����������>3�>v�&?�s�t_�*̾VR����>��H�1�O�����E>0��~��ŷ�X��>����ԴѾaJ3�Lv�� ����B�E�r�%Ⱥ>��O?�Į?��a�S��-rO��]������?��g?& �>�.?@?�㡽����р���=0�n?=��?�=�?�>	�3=�����>Y�>Ũ�?��?�Y?�}I��X?~�����
��殽]!���>��=����4�>?��?�'�����a!��it���1��xϼז=��}>M��>�p�>���<��۽�}�<pҸ>�+�>v�u>��><=K>OG�>q�v��q�'��>!a�> ��>�r,?]_�>�9D>cn+�kt8>��2>�i��p��*Ƽ�Y������s�=\�p<(���]�>	gƿ��?�Xr>�G5����>��վ�t���yZ>p��=z���t?"">m��>ͯ?xy�=�Y[>��>��=FӾC�>���7d!��,C�/�R�<�Ѿ�~z>����&�L��~��8CI�^o���g�`j�G.��?<=�%Ľ<�G�?�����k�A�)�������?f\�>6?=ڌ���%�>���>�ƍ>sK��`���ȍ�pfᾞ�?���?�4c>�f�>X�W?m�?�L0��2��MZ�`Ku�P�@�;1e���`�[��������n
����E�_?�?y?|�A?F��<^y>�m�?wA%��q��O͋>��.���:��>='��>����n?a��uԾޓþ���@E>�o?��?W�?=\S����N>n= �5?��?Y߀?Y�(?��?]�x��D]?T_	�� Y>2��>-<�>�V?	j?JE��}��=|0>פ�>��;���}��^��#�<3vH=�l�=��=��͸L�ȱֹ{8�=j&�=|ς;��};�B��������v��!>#�=IӉ>4�T?�?��C>f:E?�K̻�, ����hP�>-��2���oD��[�,��?D=�NM?��?��d?+��>��c��'W����=!Q4=��>M->���>��H�x���p�=*4%>=>K��=�-ܽ9�F�#��1ž)-<f�t=2��>�S�>�f��.>{�����t��eW>��G��_���9h��XC�<?,�@��B0�>�J?ք?�0�=��߾ ��"f��f%?"�@?�L?��?�2�=3ھ2�K���'��6�>{_,�1����0w���~4����;辆>,������_>m:���߾A�o�2�H����jg=)��5P=g	�ά־?���Y�=H�>����ʈ�XQ��&����_I?`�M=�����N��<����>v��>m�>�^�AU�Yy>�;��)0�=H[�>zb:>2V���h�ȶH��O�g�>3�0?��b?Q��?���t�d�I�Q���j�dm���4??�k�>#u*?�Y>���vB¾}���[C���R��G�>��>�$�uf�������Dc@����>��?!�>��"?_?���>d7�?�u>?1{�>��>%k��wL���/?�+p?�ށ=�,<�ҼK�`����V� f?��?��9�wԼ>�/9?�x:?��?u.P?a 4?���=Ne�=�0�7�>KS:>�mo�.���V�l=�Q?��>��Y?�7z?�:�>��G�w1b�jy`��9>!/�>t�R?'?b��>֛�>��>����	�=���>�:f?��?��m?��=�+?�G)>4��>)��=�O�>��> �?�3M?�p?�kK?�a�>ݬ5<HȽ��½}�p����//<<���;ԵL=��2l�,E�n!7=��;Ӱ��R����ݼ�j�#���U.<�K�>�t>8G��,2>�-ľG�����?>#h���;��KR��n�7�{�=�>E�?p�>�4$��׏=Hj�>���>U���'?�?�C?��;�sa��ھ8CJ����>��@?��=��l��+��d�u��^= <m?<6^?R^X�����H�b?�]?�5�d=���þ�1b������O?<�
?8�G��$�>�?�r?���>��e���m�����4b�p�j��o�=s0�>�{��e�u̝>�7?;L�>{6c>���=4۾��w��1���?��?�?��?Q%*>��n��	�#����f���6^?Խ�>l���hp!?5W�:�ҾrJ���a�����윪��p���b�������#��z����۽���=yh?��q?M�q?�_?u����b��]�Cz����W�Y��ʜ�fuD��B�K�C�f�l�{��|r���+���67=��C�7=M�S>�?�E/?fc��v�>Xj���)�7?��i�>>��bE�f�|>�O�4옼��=�I���X�`���?n'�>���>��J?�<h���>��.�׫J���4�B�b>�>�>VC�>��>�m���P½�i{��~�����sM�Nl>a?UwM?�u?悮�\O,�Ch�����Z���{*þ�;s>�$>I�>_CN�N�#���#�V�;��n�)
�2��ρ��<E=*`+?7߀>���>
@�?f�?P��F����6���{6�"�<���>��L?��>Ɖ�>v����,�ީ�>J�l?���>�@�>i���T!�d�{�nGʽ���>���>���>!p>L�,��\�X_��b��9�F(�=G�h?ّ���`��Ѕ>|R?�|�:YM<�o�>��u���!�S����'���>?s?�Q�=��:>)Fž�
�ʪ{��j��Xy4?�?�Ư�h8�b�5>048?i3�>��?C�j?�щ>�����>x!?�^R?KTK?Tƀ?���>h���'�Ͻ�)���ý9/�fB]>�~Q>"�=�B>����G��H��y�����=�i=�� c�-Q��,/��H�=fȺ�fM(>J�ڿG�K�]��(����=��O���n���>��24���\��̥��AH�Sچ�����ڻ׾�ƌ��&꼅��}�?��@Y�M�	�ž�Ʃ�ULT����M��>�6����4�_n���ʽ5������U���vLL��-e�R�Y�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >_C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾o1�<��?7�-?��>Ǝr�1�ɿc���|¤<���?0�@�/D?(�"��	��ý<O�>*�	?�9<>�m��k��I���j�>���?Յ�?�k=��]����>i?�{���dH�'"<W\�=0��=��~=�5	���>_��>�����[H۽�v>�W>��d����H���#<�j8>W'��5�ʽ5Մ?,{\��f���/��T��U>��T?+�>C:�=��,?V7H�a}Ͽ�\��*a?�0�?���?%�(?;ۿ��ؚ>��ܾ��M?bD6?���>�d&��t���=�6�n���v���&V�f��=_��>g�>��,�ߋ���O�/J��U��=I��Aؿ��'��$�۪]=B�����(���	��p=�
/<B�R��i��g	�O��\��=�/�=��s>���>���>�0c?��v?%v�>�:>G�w�EK�����{�%�N���A�PɎ�k���w��������@��%4� ��򉳾��+�C�>ĵR�!��z�L���,���l��?>��>}�ǽ�A�aȽ�~���Z���X�=���V羥�Ӿ@��F�?��)?���c�B�w���MG<F�M�U�`?�9��
���.徏��=&�v�o�8>�S�=2�>�3��$9�y�q���4?Q�.?���`ʾ��="̜=I1�=�n'?���>�j=?�=>W�L?w���E�<�N�>�>n��>h>Q�=H羳9��JH-?X�A?u���誾Xө>�E�!i��ZQ�
==ؾ�Q���>�=����V�<�Dἅ�>>)W?��>��)���m�����Q==B�x?+�?:$�>Jyk?��B?M�<l^��&�S�X�ٲw=��W?�i?��>w���?�Ͼ8s��v�5? �e?��N>Xh������.�~H��?��n?�Y?�d���r}�'�����0h6?N�v?p^��u�����N�V��=�>Q[�>G��>�9��b�>��>?!#� H�������[4����?Z�@���?|�:<
��y�=	??�]�>ϩO��IƾpP�����9q=�$�>1���hv�����J,��8?���?O��>�������y�=���b��?���?\����ґ�����-���.��7�=1]K=�1�^w�=�����1��վ"l�����e�X=�>p@�����>59G��5���ҿw�{�0n�>Q���+;?:T�>Xc����Y�.�[�sg��<7�E:?�P�z���>��E>L�'�m��������F+�`�ϽE��>%�}=�X�>U���C*���ד���=�y>Ο�>�|�>����0t��)��?]�-jҿH2��� �p=O?p3�?�@�?[�?��6�F���@���$���@?�G?��\?&�=G:���7��l�j?�_���V`�4�$IE��U>�"3?bD�>��-��|=�!>��>ba>�"/�I�Ŀyض�J���O��?O��?wn꾿��>ǁ�?�s+?_i��8���X��2�*�O%2�X=A?)2>���~�!��.=�1ђ�׻
?�|0?~��).�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>hH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?s�>`s?��k>�l?g�C>Ιо�⯽�E>\N��;�� ?��Y?4��>d�=�O���r7���M���*�Ϛž|C�m)�>��I?zOO?n`�>;�>�ih�r�?��:I��!V��^�@|ս�V��>��:B>�lq>["��E�¾��?�p�*�ؿ�i��Hp'�b54?!��>��?���-�t�R���;_?$y�>�6��+���%��A�L��?|G�?�?��׾JU̼8>=�>�I�>��Խ��������7>i�B?��D��[�o�H�>���?�@�ծ?Xi��	?���P��Za~�E��7�g��=��7?0���z>}��>��=�nv�����q�s�߹�>�B�?q{�?���>"�l?��o�S�B���1=M�>��k?�s?@o���[�B>��?�������K�f?��
@iu@�^?�qֿ� ��3T��襺��=��=Ñ2>�!ڽ:�=��7=]7�v�hP�=Rۗ>;�d>��p>92O>��;>
�)>S����!�:m��랒�^�C����{�@�Z�����Iv��n�,������tu���$ýc8��,�P��	&�3�`����=��U?�R?�p?%� ?EPy��n>G]��	��<�%��T�=;c�>y2?n7L?8J*?�ג=晝���d�� ������D�� Q�>U'I>0q�>f��>���>.�:��J>4�<>�a>���=�2*=��g���=��O>[s�>��>�`�>�S<>Ι>�Ѵ�q1��z�h���v��<̽���?1l��S�J�0���8��䥷�=��=�S.?�>���8п{��5H?=���-�$�+���>��0?�eW?#�>���e5U�'J>%��Q�j�$a>�N ��pl�P�)�qQ>yd?a*�>{�F>�BA���3�!&Z�k����ʎ>l-9?@oо�2,���V�I�L�h7�G^>�(�>t�b<�m�MW��B׀�;�a��;D�M?�?��ݽ�Z߾BrX�K���k>��>}0�<a�ϼ���>o��꙽m�H���G�(<�R>E%?�'&>���=u��>�����RX���>l�B>�+>_�<?ŗ?��k��8nm���"���l>���>�6r>zd�='O��=���>�Ac>����4���/��A?��+\>����-=m�5j�g�=�������=U��=d���?���6=�~?���(䈿��e���lD?S+?[ �=�F<��"�E ���H��G�?r�@m�?��	��V�?�?�@�?��L��=}�>	׫>�ξ�L��?��Ž5Ǣ�ɔ	�0)#�jS�?��?��/�Zʋ�=l�~6>�^%?��Ӿ^h�>�w��Z�������u�4�#=���>�8H?�U��l�O��>��v
?�?j^�ة��f�ȿ�{v����>�?���?��m��A��R@�J��>��?�gY?�oi>�g۾VaZ����>ջ@?�R?��>:� �'���?�޶?���?�H>l�?&�s?���>s�f�~�.�����t���io=44���>/>������E�U̓�~���+�i����^>;�"=��>��彉ܼ���=iޅ����\�\�*9�>3<n>M�G>���>� ?z#�>aE�>��"=�����	��0_���~L?��?m���pn����<���=�;b�QD?%�2?�#=��KϾ>�Z\?�D�?ǒZ?��>i����K��c�����<��B>^�>_@�> ���f�Q>�`վɫD��$�>[�>	����M߾������FD�>��!?N��>���=ޙ ?�#?�j>�$�>+WE�*4��$�E����>Β�>�>?��~?]?x���TW3�W���ߡ���[�G-N>��x?LZ?y��>f������HH�p�H�
��q��?�rg?*��# ?H2�?��??��A?�Zf>�a��ؾ򾭽���>��"?Y~���B���&������	?�?|~�>�y��WH׽��¼�\���0�?d�Z?��)?�[�}`�Zþr��<w�+�� ��Y
<��;��>Y!>���yѦ=~Y>�ī=J�n��<�m��<^�=��>�~�=39�`鏽,�,?��g����=�Ts���C�C*�>,�P>��¾I?]?{6�C�{��묿:�����Y���?A,�?�S�?3!���bg���:?͢�?]? ��>�~��z۾#>���|���p�[���=���>4-7��z�񣿮D��<���Ƚ��C��f�>�j�>m�?�*?r�>�?�y���Y�ң��9 �
^�{�<���-�zK�̿��6����=<���=���GVL���j>F�T�gM�>��>���>���>���>E�>��>��N�֠�>�c�>��
>�iu><�A>�m���ND�5LR?�����'����+���]-B?End?L5�>�ei���������}?'��?�p�?�4v>#yh��(+�El?�1�>d��k
?ѯ:=;3��Z�<�X�����H*��yu�ѧ�>�%׽k":��M��nf��g
?�*?�[����̾b2׽�3��~�m=�Y�?�<)?��)��R�4Xo�X�c[S������g�^J���2$���p��Џ�G]��������(��Q!=�f*?�?K�������k���?�>f>�~�>fǖ>�S�>p�I>�	�]�0���]��'�=w��2��>+A{?<j�>��H?w�6?T7>?�@? ��>Nd�>����f� ?��ɼ�aX>4�>�� ?�@ ?t\=?T�?|�)?r�,>04,��J���Ҿ�#?[?-�!?�P?�0�> �Z�l�z˽M�~����Z���l�p);�F��~�Ȼ }�=�d�>fX?-���8�����k>?�7?���>���>���#-���<�>ҵ
?xF�>�  �x}r�c�\W�>y��? �؁=S�)>���=Y����<Ӻ�W�=����?�=/-���y;��w<E��=e��=2It�4쁹���:Wz�;�`�<Dp�>�?6��>A�>:��J� �`��k�=" Y>(S>/>wJپ.~���#����g��_y>3w�?�y�?��f=��=B��=�x���Z����3���v#�<��?�I#?WYT??s�=?�k#?��>�#��K��-_�����~�?]>?w�=u��ic��@^��L�J��q?���>md��%�S��.���|�=��>&�4�U=<�C���y��d%����{zܽ&v�?�^�?w����A��%�����z<ɽ��.?��>8*�>�V?����	�C�k.0���>E�Q?��>�})?J3l? �U?�K+>]����͟��9u�)��>M?e?U#v?���?�I�?��?�`�Ǣʾ�8�����������"���sy��2x>a�>�K�>��?�b	�eY̾DR�x�Ҽ.x:������?���>d�K>j��>�-P>C0I?���>��������龍H&�-˽=�s?hϐ?�N?�bw�����*9�0��2d>���?3�?2�?4H|�a�P>�]
�)پJ���L=�> ȵ>���>��=�4ɽf�?_?���>�Xc����1�5�x��~�?U�'?dE�<��ο탿�F~�����j�<�v����M��G���a��	�=z���V� ��	&u��坾E-��֨��x����D��.�>O[`=�)�=e:�=�Z)=�󑻵��<� =�U+<F�#=pJ�2��<�KL�Rp	���x�h�<��_=���=�.���!���z?�5I?2�2?$�J?��g>ɦ�=2�=([>���0�?<>;�ټ�-˾�����L�������1ɾ�⾢;�y���Ye�=�o�LZ>��W>g=��<)_>lZD=o�=��6=��=оg<�J�]�>x�>�0!>�+�<�,x?�S��?��Y�O�� 
���6?]Ŗ>��=�W;m�;?�BS>7����Ը�{���u?��?|�?�?2{��X�>d������]�=~���
>N��=Ml5�g��>��_>�������$M��dD�?�o@�;?d-����ϿXt&>�bl>`��=��j�ld1�#�����3��F�='?K?1���Ծp��>BF�=����_}5�#�P>X�=�Q�wN]���=��ܽ{�=�=�$�>���=�u!>��������G5=��^>���=D�	��q@�҃q��԰<l�5=��2>�G�=�v�>�?3h0?uLd?eb�>��m��wϾj��n�>��=��>���=�C>>�>��7?�uD?�iK?��>F��=�ݺ>Ǧ>!�,�a�m�^\�ꦾu�<���?Y��?g��>�G<fA��E�='>��}Ž�?=/1?|?�e�>����eW)�$5�y;�}�<(d�=�����&�kQ�<k'���SȽA��=���>�/�>��g>��>$��>cip>v�>��>1�.=��=�m���mo;�����g�=�z�:��	=��\��.���*[��Pq������b-���<�g�=��=�H�>ܐ>��>��=����0>��nUL�/7�=����9�?�́d���}���,���<��P:>:�X>j}�
F��.$?�'X>�@>Zi�?Wrv?D+>Mg�9@վ)Ɲ��Fb��GX�I�=��>�B���:�7�\�D�J��о�!�>��x>�ȗ>
7�>�$��"7�:��=|� �x)��)�>y��]?�|	R���h�� ���ڞ��v�s�ʼ�z0?|ٌ�.	>��m?w�>?�ߖ?�?��=;Ϥ���>�����m�<�g�7����׽�C?�8?S?)����5�K̾S侽`ѷ>W_I�iP�x���}�0�5g�e���*��>�����оX!3�me�����e�B� Yr���>v�O?��?|b�ZU���WO�t���
���l?�yg?��>L?m;?4"���x�d��vu�=��n?:��?�6�?+�
>�sǽ?a�p��>3�>Ɋ�?�?߽z?����44�>} �SW;�翾7ܽ�q�e��=x�=�Z�>�m!?�#?�l�b��&Jþ� �B�'����"x�;V;c>ů�>��>O$�=)N#>Õ>�R�>	 �>�Z�>��>�/�=3L��K���� ��?��>�+�>��?�%�>�zE<���=��>Ż,��e��>ӽ���ZO�A\=)Q�=�Q���㽍.�>[)��~S�?�>�����>�꾔�8�8�/>E>��a�� ?z1�>a�=<ѝ>�'�>�>�_>�<a=u@Ӿ>x>���^!��+C���R�̽Ѿ6bz>V����	&�h���r��
II�,m���d�Fj��/���;=����<C�?������k�W�)�P�����?7k�>�6?�ڌ��"����>U��>���>�O��ٍ���ȍ��^ᾫ�?���?��b>��>��W?��?!�0�j2�gDZ���u�)A��e�V�`��፿�����
�a���;�_?	y?ŋA?C=�<�y>���?x�%��
�>j/��;�"j<=��>�����`���Ӿ�þq���KF>^}o?/	�?TX?�]V� Ҝ��$>g9?�((?�sw?��1?�:?S@�S�%?m�%>�� ??5?�t/?$?l�?�4>s�=��<�nt=�0��a�����~���¤�	mY=�1=���Kx\<��!=zҔ<�l�:5W��zI���k$�<�}b=�3�=��='�s>�O?��?�ޔ>#�M?� <s��ӳ��H?>�������)��P���0�q�m:�R?��?Gh?Jw�>����I�����=fy�>|��>kOY>5`�>.{X�|vƾ<�&��5;>��������_��oLϾ	���懾�19>��}>�O�>N`>�Ҋ<��>0����nL��z�=`����Y�R����f�G�j{�>)
=?�4�>�	ϼb�����<��~��?
?b'1?GM?Ψ�?��>j�_�"�/���$���V|>�'�=��,�F���<���:��1=7J?漧��͑�%fr>��`��}qt��B��3�a�=o/�f��=����ھ�S~����=���=�ش��!������驿�rI?'=Zu��[7����I�=#�>'X�>g����쟽K�6�vj��v?�=���>=#>.Z���z���G��D�A�>�;?_�j?�}�?��Q�fsr��SB�;��A �{�?��;?���>IT.?�U_>;��k���w��yT���:��H�>\��>�<��M�娼���ɾ��+���?>��?z>U�?%hp?���>�]?0?F�>�¨>ok�����2�.?���?�]�=��e��鐾}��4P��5?��?�VB����> '.?�x1?��?��&?��'?̓>�W �T}:�oŹ>}�C>+#r�兯�k�=��8?0��>��h?��y?6@�>�kF��/���B�5�v>��>A�9?�,?���>b��>�\�>�H�� 0�=��>��d?�?3Ao?֕�=H�?�o">�^�>1�V=��>q#�>P@?:qF?K:o?JJ?���>�X�<|鷽u���/9�+��:�(�<qBU<Q�J=��A�D@���μ�RB=�Ŭ<�0��aJ������3����}%ټ���>��t>V���в1>� ¾հ��L>>gz���D��T,����8����=|D}>}� ?Ó�>�$'�	ś=�c�>���> ���'?�?ۂ?�&<"�`�� پ�#J��.�>��??z��=vJn�R����$u�c-\=�l?T]?[:S������b?��]?��;;=�h>ľ�sa�e	꾧0P?\�
?2oG�O�>9?�r?�e�>��e��Qm�+̜�D$b�]�k����=�>����e��՝>�w7?/�>�yd>��=BFھ%�w��V��
�?��?L�?��?M�)>[�n���߿�D��j����]?�E�>���; "?9J�:�Z̾�*��i���F����R���=���2�&����$[ͽ`�=�.?r?��r?�w_?�'���c�w^�xC��/0W�y�����[F��hA���B�^�m�L6�Q���	0��:�7=��Z���c�OB�?f�?twn���>90 ��F��K��� ��>�'ݾ�����&�=�P�x�>!�6;[���������ʾ��?V�>\�?�MK?��U��mX�U�L�W�C��3��>R>~��>�7>B�-?t��=_��!�1�s�$�~�ܾ�jӽ�Ku>Ooa?�K?�n?<����)1�8"���[ �Tf�9@����J>�B>D}�>gMS�l��%��K?�Jp��w�@���l�[�=/f0?K5>�[�>�;�?��?h'�c�������^N2�b�;C��>Vbe?̤�>�-�>i-̽������>��l?��>f�>_���(L!���{���ʽ��>]˭>@��>��o>&�,�l!\�Ih��ہ��h9�'u�=��h?i�����`��܅>*	R??�:&�G<@v�>_�v�'�!����)�'�m�>#r?f{�=Z{;>
mž���{����W@?8�?ɥ��Z8��\M>�{'?x{�>Ɍ�>�e?!	�>A�޾d�^>��?g�A?X�5? �`?��>}���1�+���{�z[(����y�>��>��=��>W:�$�H�_E;���=��V>B�����T�Ņ��Yo=`O��>�޿D_�\���Fk�;���x��vq���}��Γ��4�������V���ɯ�Գ�4����Y���_�I|�?9�@�悾"׶��Vh��YD��n>�Z�;�>N���y|D�1�!�(���󥊽�-��T��+D�Eـ�Q�'?�����ǿ򰡿�:ܾ3! ?�A ?8�y?��7�"���8�� >#C�<�,����뾫����οC�����^?���>��/��u��>ܥ�>��X>�Hq>����螾x1�<��?4�-?��>��r�0�ɿb���.¤<���?/�@�}A?1�'��쾎�U=L�>ʝ	?M�=>�1�{�1������>&�?9O�?�D=E%W�b �1�e?O��;R�E���)�6�=|�=�I=��	�s�L>T�>
���<��gؽ0�4>��>�"�����{\�⎀<�M^>�eĽ�<{�5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=g����Ͽ�$�d�Î=.F=�{,�~w̽��̽Лƽ%r��� m����f�<"hs=�m>6�n>%`x>�d>�b?�dn?y޴>�`>	zT�U���>�����潁����н���;OD��#����	��,;M?�m ��B���达�3�yď>�SQ�i����J��#�p����;?P�>uuB=\�C�� ⽒�D�;���n>'�W�������|6n���?g-S?A炿��v��3ɾ���zI�d0r?�~O����������=򡌽�Ǻ=<�r>a'u>Q|���eG���E�YS>?̯?h|��ᵋ���>#��=b��)?�'�>���Ph>3�X?�{x��,G�\�=�<u>T?���=���=�"ʾ���g� ?��<?+wּ��-�"�b>v5þ�����<�d>��侔��.c�=�,�<v���[�>�"F>]�>@"W?Ҡ�>o�)�w���K����* ==p�x?��?��>!sk?��B?�4�<uj��?�S�k$�a�x=W�W?0+i?r�>�e��*�Ͼ o��,�5?_�e?=�N>`Sh�Ԭ龈�.�@[���?d�n?�V?�	���l}�&�������6?��v?s^�xs�����L�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?z�;<��T��=�;?l\�> �O��>ƾ�z������4�q=�"�>���ev����R,�f�8?ݠ�?���>��������>=������?~u�?G����x?����j`T�ʉ��D>�ّ=Έ�xq+>�.���a)� $���#.�:Ч�ε���p�>U�@<<��#�?6q~�S��ɿӿ�����o�+���A?3t�>\�	=#��&o�bb���2�s�M�NF��4�>'>� ��ji����{��:��\��Z��>Ł��É>�T���������ȗ<;ђ>�<�>m��>����Q]�� ��?G���$ο�_��I'�>&X?!_�?j�?J'?�<��v���z��.�s�F?�{r?�7Z?�e���^�h@6�%�j?�_��wU`��4�tHE��U>�"3?�B�>S�-�_�|=�>���>g>�#/�y�Ŀ�ٶ�=���Y��?��?�o���>r��?ts+?�i�8���[����*�\�+��<A?�2>���I�!�C0=�UҒ���
?U~0?{�c.�3�_?�a�#�p���-��ƽ�ۡ>��0��e\�,I�����Xe����@y����?M^�?g�?V��� #��6%?�>`����8Ǿq�<���>�(�>�)N>H_��u>}���:��h	>���?�~�?Pj?�������U>��}?���>���?���=h��>k��=츰�o�1��	#>�=�^A�Ӣ?	�M?���>���=X�8��/�dCF��
R��
�P�C��*�>q�a?�2L?�b>����/��� �S�̽;�1�2)！�@��R/��a�κ3>��=>>��D�R�Ҿ��?Mp�9�ؿ�i��p'��54?0��>�?����t�����;_?Nz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>A�Խ����\�����7>1�B?Y��D��t�o�y�>���?
�@�ծ?ji��	?���P��Ba~����7����=��7?�0�#�z>���>��=�nv�ܻ��Y�s����>�B�?�{�?��>�l?��o�L�B�F�1=9M�>Ϝk?�s?[Io��󾀲B>��?�������K��f?�
@|u@e�^?%,��3��C�ľ"0���?�=b��=o�6>|���U�B>A��=���̖���&->�ԟ>�a>��R>6�Z>'n�>=�>��JI"��-��Y$��u(9�9O!�E���W4��*վ~*������ғ��7Bؽ�k�󄕽Mn�������m��=_�P?�ZQ?6p?n��>G����>���}7�8�-�cʟ=4I�>�u-?�6H?�#*?�b=�)��a ^� U~�XA�����o��>;>H��>�G�>�R�>��};��K>u�1>'~\>ҍ�=��	<�^��Q��;Q2F>�4�>�>1�>!��>�"~>xa��/9��뾁�h�A�)�D�ܰ�?�D��t������_�������"�41�>/��>��q�"ž�L-���hJ?0�⾩��H=I��h��>v��?�O�=-\����z�>�	ٽ"���zՖ>��ѾJ>>�v��K�l=S�>�^�>�[>��A��`:��\��Q����>Z�6?.���WU�۴`���H��a�bj>\[�>���<J� ��ʔ����4�S����<|�7?�?zH���Ӿ1�a�O֡��>H�]>�8�=v|@=� b>�h�<z�����`�t╼�;�=C4>�?��3>8��=P�>�L���&�m��>8�8>�e1>"-6?��"?3x��6⣽�͇�j�-���H>z�>ǻz>n�>t_���=��>�wb>~�c<�v-�Q+��W6�	�|>������{�<���T�<WԨ��W�=_=����Y����>�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾLh�>vx��Z�������u�1�#=X��>�8H?�V����O�l>��v
?�?�^�ީ����ȿ3|v����>T�?���?d�m��A���@����><��?�gY?�oi>�g۾8`Z����>ϻ@?�R?�>�9�v�'���? ߶?կ�?�BC>�0�?�*q?L��>�(�����X�������<ݼz��o��>�|5>����[�F�ʔ�����;PZ�	��-�:>�*`=��>��	�>_ľyb�=DƗ�󰾢�7���>�GD>�\>�ө>0*?��>��|>�#�= ��:��^����M?���?����o�s�<��=K�e���?��1?MV0���о:m�>[}[?��~?�Y?�Ğ>���[⚿+d��j����<g�9>��>���>�Rz�@%O>�Ӿ�@��h�>w��>
�ͻ�fݾ����޺�\P�>z�?���>��=�� ?��#?��j>:(�>�`E�Z9��g�E�7��>,��>�G?D�~?]�?Dҹ�~Z3����?桿Ց[��9N>��x?V?�ɕ>T���
���ڡE�V>I�&���i��?�tg?4L�t?�1�?��??S�A?�+f>����ؾ������>×#?ԉ���A��V'������?v?�D�>󱑽�Խ,F��!�[h��ǯ?��Y?��(?�|���a���ľ�"�<�?G�Y/��BR<O�ͻr1>�>}����s�=-�>)��=��c��&=�ү<<�2�=*>�>y��=��:��-��'=,?m�G�pۃ���={�r�3xD���>�IL>�����^?yl=��{�����x���U�� �?���?Xk�?	��9�h��$=?�?P	?l"�>�J���}޾/�྘Pw�~x��w��>���>Z�l���H���ۙ���F���Ž��-��.�>���>]�?=A?�/>/�>�E0����rྱDҾfP@�a�2�23��&� 0)������,ݽfn��¾\l\�09>k0��Dh�>`t0?Wr�> ��>��>k�<��>�99>,H�=M�B>�)�=�G>=b�>���=����YJR?�����'���&���S3B?�md?0.�>�h��������~?%��?�p�?75v>�~h�8'+� m?�A�>F���p
?�g:=g����<�R����01��������>la׽�$:��M�Inf��g
?�-?�-����̾��ֽR_��1�h=C��?�P)?Z*�(OR�9Wo�'X��S�"C�J3f������$$���o�I���G�����$$)���%=e�)?��?��r��֫�R�j���>���e>�,�>M��>+��>D�I>��	��2��t]���'�� ���p�>Y{?���>�/G?Y9?hM?x�I?r��>���>t��P��><��:>
��>ǭ4?ݧ'?ِ,?BL?�.?4�_>P�ڽ1 �uѾ2F?Iq?��?��?# ?Z6������%�μ��n'�������a=�?x<[���\�9ݛ=�>X?���w�8�����k>�7?;r�>���>e���3��3��<��>��
?�9�>R  ��qr��\�XB�>J��?H���=�)>���=Pi����˺h�=� ¼G��=����2l;�!�<�d�=�Ȕ=$~�(x��~�:Wi�;�s�<�t�>9�?���>�C�>q@��� �`���e�=�Y>�S>}>�Eپ�}���$��r�g��]y>�w�?�z�?��f=��=��=�|���U�����:������<�?CJ#?XT?P��?X�=?Lj#?ŵ>+�ZM���^�����Į?�+I?�zF=> 0�k?�lᵿ��`�{�?ퟅ>]�]��j	��ڛ�P����i �>YR��xK��ר�6>c���s�e�X��d�?^p�?�;�<G�D��IѾ���ٖ�39??�t�>�Ӝ>�X?���	<��W:��>�F�>�X?e�>w�&?��w?��j?[~M>��f��ҥ��8������Id>Dه?��?�?��?���>��.�[>���ĺ�t����sս�Aľ�|�3�}>}>?w��>3"�>�SG=�+��_�2�/��� �������>؏�>,5�>��>x��<�G?���>�������jV��b�����=���u?��?�[+?
=�J���E�;l��$��>i�?#ӫ?�)?CT����=��ܼn�����p�Ա�>�>Q��>7��=� C=�>�K�>s�>������8���K���?��E?��=}�ſEq��Eo������o<{v��
�d��{��h \����=�3�����r驾�[�s���֓��ൾAK��4{��p�>�B�=���=�#�=�<7���	�<�K=0��<�?=�p�1do<��8�.P����������s<�^E=�����'��͢o?԰M?	�,?��8?��>�u�=��Y�1��=��d�?3��>�4���kȾ�2|�O?��0i��p�ɾ��ƾJ;��xV�H��=v���d�>�JT>ҙ�=[==/-�=�ֻ��=�=X��=��<`Jg�p�	>�qB>4�g=�\�=�6w?V�������4Q��Z罠�:?�8�>}{�=��ƾj@?��>>�2������tb��-?���?�T�?8�?Sti��d�>S��~㎽�q�=Q����=2>y��=y�2�B��>��J>���K��1����4�?��@��??�ዿ̢Ͽ#a/>���>f�->F�R�9|2�i�E�� �$7l�_�,?/�+��Ǿj#>�>�Cܾ4���dT<<��>��=�u����W�^��=*i��W�D=��=&d�>�o>���==�����=�����=�p\>�,����}�G̬��F<Lf>�w3>S�#>���>I�?0?�c?���>�Tj�?wϾ>ݿ�^!�>T�=A��>.؊=�@>�}�>�6?��B?HK?O)�>W�=t��>5�>z�+���l��?㾙¤�j��<"�?��?���>�B�;��H��K�@�=���ȽX?��0?�
?`��>�U����%Y&���.�����`e0�G+=�mr��PU�����=m�@�㽖�=�p�>���>��>JTy>�9>�N>t�>��>T6�<�p�={݌����<� ��p��=;�����<�vż���tj&��+�V�����;Ǵ�;,�]<���;ǒ�=w��>�>���>=�=;���sU/>3��*L�d��=�B��D�A�^4d�F�}�R�.��z8�a#C>^�W>�_�������?^�X>-?>���?%8u?�s!>��
���Ӿ�2��6�f�U�U�׉�=�$>�=���:��_���L�0�оm��>Az_>@�s>��> 10�E&`��K>��|����>��v�Jm��e���J��I��Hi���_��}&�F�?�����J>�<L?�p$?�Q�?�Y
?B�>�ü{��>�r���̽����xen��?%��>�?������˾����kʶ>v�E�Y-O�ƕ�@K/������;�>U��\Ѿ��3��(�������=C��s���>�N?/�?a��u����N��D�<<s�<? �h?���>.	?f�?d��H�(����}�=�qn?��?�_�?ni>�3!�<=c��>}�>l��?�tz?�j?�&��� ?+Q<�}롽������J�a�>>2>�,?�SK?v
J?ʦ罦}	��䏾cn���)���K=�G�="�X>5=�
>���=��Y>-�h>��=Q�^>�@�>dI�>*Zp>m�=\��^u%�7?�0>��>x�?7R�>1��>q4%<z>���;�k]���������w	�]v�ÿc=��/>�毽Ъ�>�Vÿ�ڪ?�=�� ��>Y׾ւm�i�=��>9��4Ҧ>v��>엄>�>���>p��<Y�>���<�-Ӿ�f>3��TJ!�O-C�R�v�Ѿv*z>י����%�������9I�ya��o��j��+��!B=���<�8�?�d��^�k�6�)�m���D�?�m�>�!6?������9�>���>��>�^��M���ō�QF��? ��?��b>k�>��W?e?�/���1��.Z��wu���@�� e���`��э�q����
�/u��J�_?�y?��A?��<�Hy>�z�?��%�����T�>�/���:�6f:= �>ϐ��A�a���Ӿn�þ����3F>t�o?1�?�A?o�T����ا=�f>?v*?�܀?�a??�!??׎g�Š)?�γ=���>^��>�(%??�?5��>~�>P=0>>��<��>7����u���+���W���<��=pH�=r�8��l�=�/=R��<���<V�e�1Y����<�<�=�G�=���=�m�=ig9?�U?��=hp>?d�;=ԕƾ�F���Y?��o�%��˅Ҿ���~�����>#�Z?��?i?V�5?�GQ��5�6c8>u�>���=D��=n@�>za�y����<>��>D�d:V�y1>�u���m�~��Щ=��>���>g�{>8'��Z,(>�K��$z��{d>IR�PȺ��S��G�N�1�؂v�jM�>��K?�?��=�.龸����-f��)?H<?L#M?Ⱦ?X&�=2x۾8�9�ҙJ��s�b��>���<Z		�Һ��N���:����:fts>S➾*���G�>8G8�����u��C�I]�u�~�(�(�%�;>7ۉ�띾�膾�m>1�>����HA�_윿������q?���Xl���W=���f�=��>�T�>�A
�*	>���S5�`L�=��>l�/>�νUw��@J��>¾�ٝ>��!?G�<?�R?	���:d���j������S��_�����>�۠>��>��y>i��=�૾��(�1���
"A�b�>�ٰ>��Y��-�ӏþ+^���%���=T�>?@?^>�̪>�p?_�D?�-�?ciW?�{&?�e)>rP�;W"��A&?)��?:�=��Խ\�T�� 9�OF�"��>b�)?��B����>;�?ݽ?�&?�Q?��?��> � ��C@����>zY�>��W�mb��V�_>�J?욳>9=Y?�ԃ?T�=>C�5�	ꢾ_ש��T�=:>^�2?�5#?@�?���>$w�>�j��z�=���>�!c?k0�?0�o?���=z�?�"2>���>>��=㬟>Dt�>�
?�YO?��s?��J?��>里<�k��5��ojt��xN�2��;7�H<#�y=�(�7t��3�H��<*I�;�������Y<�_E�����h��;�c�>�s>����0>��ľ
X����@>ǝ��4���Ȋ�=Y:��7�=�t�>9�?w��>�~#��=Z��>fH�>���u2(?��??��*;B�b���ھ߃K�$�>��A?���=��l����[�u�M�g=#�m?S�^?��W����m�b?��]?���G�<��xľ��c���7NO?/�
?��G����>Ó~? kq?���>e[e���m�D����b���k�
�=&&�>����d��_�>)�5?Cu�>�a>El�=�ھ2�w��ើ�? 0�?Q�?:!�?�c)>+8n��H�?���E2���_?���>Z��W�#?����;0M������f⾔���dh�������3���$�����޽���=\�?�Ur?'�p?��_?����b�v7^��:��*�U�>����QzE��D�4B�7�m�Z������-"��

L= cC���H���?M�'?�����?3���Ƶ���޾	�8>x����n����<bѽ��<WD<=�*i�����i���?ka�>\X�>��??�(_���.��\9�CE��wᾒ#>�3�>�oz>���>�S=���*�Q��	ƾ��¾�6���+v>�{c?߀K?!�n?.��"1�����Q�!��0�q���B>�<>���>�W�Π��,&��U>���r����)u����	�^�~=��2?K�>���>5I�?`�?7t	��[����x�{1����<��>i?%+�>�φ>�Ͻy� ��7�>fyl?��>F��>����� ��{���Ž���>v�>i��>n�m>%$.��\�hc�� B��7t8�E�=��h?Tl��i�^���>�Q?4w;K�i<_��>P�|���!� B��)�U�>�4?�2�=68>�VžKt���{�i���P)?D?t蒾Ü*��0~>�"?�q�>\0�>3�?�5�>�VþeN���?a�^?CJ?KA?E�>��=4�=KȽL�&��-=i��>� [>�Am=H��=<��b\��y�3�D=e�=D?μ�_���<����ZzL<��<|�3>��Կ��zm�.D�����MǾ䥾Ų�
w����� ������R*{��(��9!�୧�^nY�\�i�)�����?Ir�?�پ�>��!����Ά�]#��\�=B;��BWe��
�Qt=�>�������4��$�+�7j:��~������+-?�����gɿOឿM���#?��(?T$`?N'�<���%�+�W��=w�y=K}M��$�������ɿA����g?:��>�n��������>��>�lS>|�>>���ģW����@|�>��?���>�ʪ��Sƿ>����p%=e�?��@S�A?�)�'Z��D=<��>�%?r{E>��,�=���߬���>�I�?��?-�K=n^V�-8���c?���<?`E������h�=Г�="��<Cj��5C>��>�X��:�FZ̽rd=>G�>�i<��9�%�_����<�e>�7׽���5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=CK�h����m.�4�E�ʊ=��=,�r��9:��Ӝ�$��<[����~��᧜��c>�N>���>�-�>���>ĢT>��g?�?���>9��=�T\�h�\�Yh龿6½���|�=�
 ��?p��}����׫۾�j���*�`(���Ǿ5<�ڳ�=�#Z�Ua����!��A\�x�I�_?߉�=�8��=���&��$Ͼ|���#����㓽������3�H�r�C �?c�=?���R�>�b��>�������)H?�|+����/P��'=>�����=���>��$=~0��>�4W���1?��?^�����u�<�>�gY�K��=�K?Z�2?ǥ=K1�>�6@?�b������BU>��л�=?'��>�:�> �����;/(?'�S?5�ʽ�Z�7`>��4C��&�P{<��z��>"��=k8���uŽ*���6A,<#_��W?�_w>F�)�pY��V��!���!��=�u?Q8
?�~�>ɼr?�G?6K����UZM��x���=Y�V?/�e?�>D�e��rɾ����3? �a?��6>&_\�/ؾ��(�VS���?�q]?8�?��\���t��������|7?��u?��c����� ��"c���>���>2,�>6�4��~�>)�0?@�yb��1��$�5��D�?	�@�X�?��=� ���=9�?�N�>c��}����q^��w��w���>/�̾��r�0����򽉺/?mq�?��?+l>��9�>=^����?Y�?�뫾��>�u��cN����4�j�\A>�Kֽ^�y���-���EX�!⾴��=��z>r�@����"�>pD��װܿ��п�䈿 ���I���]H ?�6�>T��@eo��TT��7u�v\G�MO�쭾���>+�
>%ǰ�LW���lu���9���ZJ�>佾�K��>]$����;����;�̏>g_�>�t>�g������?�?�
���ʿ���UM�C?B?���?�؇?��#?�U=ԁ+�tt@�f<ijF?��g?yg@?%�r�97�U�I;u�l?$�ξ,lh���4���L��=>��+?C^�>������= 	�=T�>�>��8�������X��;��?SP�?�"ݾ8y�>wr�?P&(?�5	��o��r/Ӿ�.��U�<T�?�7>�b��M)2��)A��C��˹?4w9?Q�U�N�_?�a�2�p�Z�-���ƽ�ڡ>e�0�#f\�MD��Σ�xXe�����?y����?D^�?V�?���#� 6%?�>�����8Ǿ��<���>H(�>)N>H_���u>q���:�Ij	>���?�~�?�j?̕�������V>��}?�!�>�?�o�=�d�>L��=�밾��,��h#>
�=2?�m�?�M?4D�>+F�={�8� /�wXF��DR��#��C���>��a?SL?�Hb>g���32��	!�ԉͽ�g1�H��/a@��,�G�߽�5>��=>h	>��D�gӾ��+?�
7�x�ѿw����z���&?��v>���>�2���x�O�f��u>?��c>��-�A���a��j��d��?Dn�?� �>� ƾ=8�=��:>��>$�>/��̀=�6h�����p�5?���lf���Bm�c�|>/Ϳ?l:@6��?��d�@d?������"mu�j��}�j��B�=]w=?�Yվ�Y>���>�=9b������8�s��Z�> �?LS�??��>6�V?j\�Ae�J K=k��>�0b?@?=�W<n� Nu=U2�>�L�����O���xY?+		@�Z@�Qe?}d���׿�n��~[��{�¾�.�=�р=F�C>a����=s
�=e�<�\��m#>}K�>	�v>~�>�H�>s�F>�| >^i��Sy!��5��K���Z�z�!���G!��m��XEH�Z#�J��J�����Q�Խ`�ҽ��a�#'+������=kb[?R3Q?!Rt?�?-4�J�2>V�����<��-��"�=�j>��.?m4G?�C%?�ɭ="����8_�����槾�b���>��F>5�>D��>A��>�y�Q2K>%YW>=]�>>��=Ħv<�Ҽ�~/=Z]>��>B�>.�>D<>:�>Lϴ��1����h�w�9̽� �?ʁ����J��1��R9�������i�=)b.?�{>���?пS����2H?����;)���+���>s�0?dW?��>u��4�T�<9>����j��_>%, �1�l���)��%Q>�l?��f>�*u>��3�_8� �P��y���a|>o06?���K9���u�E�H��fݾ�;M>0��>S�C�ql�m����� qi�V{{=w:?�?aK��Cܰ��u��G���PR>�?\>0=�o�=�JM>��c�׼ƽgH��=.=P��=��^>�?��k=���E�=>ý��j����>L�>뮴>l@?ҿJ?PJ>b7��F�L�:���c��?�΢>qwx>��E��b>��>��V>�j�=O�"=�[[�qH�Q\p>E�轏���]ꀽ���� ��e>y��= W�$T�1�>�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ���> ��m.��K؆���v��8'=f)�>��D?�#񾞵�2@�j�?�?�C���B��&ɿ5�u����>B,�?��?,�l�����u�=����>Fr�?��R?0�x>��о�*d����>��=?�N?�Ѫ>�Q���&�	?-��?i��?��H>/��?��s?`�>�w��M/��-��d����}=	I;�1�>3>1���LnF��ړ��b���j�\����a>�$=|��>�Q佒K��K�=F����:��=�f���>Dq>��I>�g�>�� ?�F�>鱙>s4=����'瀾-���^�K?���?��n�{��<���=��^��?�S4?H�W���Ͼ��>+�\?jɀ?[?Ĝ�>a���7��y鿿ٌ����<J�K>B=�>X�>f���;dK>��Ծ�qD��;�>�ܗ>����eھ!M������K�>|!?�s�>��=$#?�7?y-1>'��>:%@������%�K��>��>h�?G�?��?�r����#�?ჿ�ڠ�M�Z^�>��[?1'?��=����t=���@O��/�\N=c�?�Cj?��ǻѓ+?R��?��,?%�=?$�1>'߈�n=��pe�N�>��!?3����A�R-&����^?�H?���>�*��:�ս5-Ӽ���F���+�?/
\?�$&?���ya��þ���<�o"��mP����;:�D���>	�>��@��=}>WG�=mHm���6��_<��=MZ�>���=p$7�ꍽ�g,?}
�;�D� �B<�`[�43 �Wxk>�Y>֍�P�?h]���(i�,o��`������A��?���?�l�?��=��
l�|K?#�?M3�>�a�>�.P�q^˾\�ݾ��ƾ蚾�*���ڻk�>Sc>t&�[A��{����r}�|#��s&�~�+?�\�>��>FB?m��>hv�>��4=#�O���X��F���j���辿|G�bi\��" �P���IP�U!l=��<罬�>�$�)-�>���>�4�>?�>k�r>RW>�>��>-�>Ro�>m�>�v">@��=����j^�CLR?R�����'�7�� ���&B?�qd?/0�>I�h��������2�?��?�n�?f1v>�h��'+��q?�<�>����f
?��9=|���:�<�Y��<���憽<�����>�׽�:��M�8ff�`d
?�&?����̾��ֽW㞾�j=�W�?О(?h�)�DP��p�O�V�:�R�jM���c������p%�G�o�@l���h��H�����)�E�3=;�)?{�?Lm�K�������5l���?�ݗ`>2L�>�1�>׸�>�RM>%��L�/�}�\��&�ވ��MD�>�x?4�6>~�e?)T?z�p?>1c?�ٮ>g�>��f� ��>\L�<E�>���>K�A?#?r� ?L?8S3?>�E>�3����B�ʾx� ?�R??4?8��>Hף>	ƌ�KӺ0>o'>�"�?��U�<yD>�K�=����c=��s>`�?�c8��;�5����9'>z�$?���>l�>зg�<MB��t�=��>�H�>M�>5���z�x� ��D�>�i�?�Ｔ��<am>�z�=b�ػi�;�e�=���;�=u�@��L��p�<�Z =7��=͡/��Y�:-�]=�\	�C��=�<�>X�?m
�>d`�>���)% �l�=��=t�W>� R>S�>�ؾ9&������k�f��%w>���?D��?9�Z=��= :�=����^d¾�s	��翾zX=O ?��#?�GT?���?[V>?�#?�!>�g�g���E���P���L?�!,?��>�����ʾ���3�2�?�Z?Z;a����;)�K�¾2�Խ��>O\/�0~�h��+D�f䄻"���������?j��?dA���6��z辝���:Y����C?��>�X�>��>��)���g��$��3;>���>�R?)�>°�>�z?2�Q?w_�<����`Ž��J}�@�>���>��>y�?rү?� �?@z?�\?s�.���߾:X���=╽*��8�T>U�>���>���>pU<>�pD=��=���<�Խ\�T>��W>'��>Yp�>v�>Y}�>�����G?S��>�^��M��f�:̃���<���u?N��?�+?Ż=$z���E�!E���E�>�i�?���?6*?�S�#��=Z�ּ�޶�o�q���>�׹>r2�>]ړ=luF=�_>i�>���>E/�^�yo8�cPM���?F?e��=� ƿ�q���p��ۗ��6h<�ܒ��d������[����=��������ʩ���[�����j��M뵾ᘜ�ؽ{����>O��=:��=s�=���<��Ǽ4м<n/J=X*�<�,=�Bp��k<k+9��Hϻ-p���#�3,]</�I=x��}�ľ�}�?(B?�u3??�Q?$��>��>y���p>���?�>�﻽/ƾn�/�z���?��_�Ӿ!��6`K�d;���/>nk߽\��=�A>�r�=�h4�a�	>f�=�1=��=�(<>6�<�_�==�a=���=:�5>��(>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>|6>dx>��Q��-��HN�C�b�%NW� ?,�:�:d̾ٹ�>bK�=�@�r�ž�J=C,5>��T=�t�ϗ\����=��x��%F=o(L=K��>j�G>6�=桹�w�=�5Q=���=|�J>kԛ�ns�8$:���=��=_a>W.(>���>�?
�.?�0c?�˹>��l�AE;6þM��>Gg�=+��>G
�=y>>�>W�6?H�B?�I?~9�>��w=ͽ>l�>4-���o��|쾉Q�����<���?u�?/��>"c�<�4��0��:�R½=e?�1?��	?翡>X��m�{�'�y�f�X�񽇱�@�=��¾cf�<.�>����)-����M>ci�>0��>��>ɰ>�0�>x�>��>�F;>�	���QO�=%$>C�佋�0=Ǧ���=�c5������M�A}0�%�x�'=!�d=b��=P.=��>V��>:gR>I=�>�/�=�`>���	>��"���J�a�b�<�쾹71�)S��g���@��At��L->;�>J_�=Đ��:5?�(�>���>�?��b?�S�lǅ��:���	�����4jþ��=��=�m���X/������r��b�����>��><�>��l>��+�P?�E{w=����g5���>D���2��W��2q��@��b�i��E��?�D?F��8��=�~?V�I?�܏?7�>�qsؾq0>�K����=��xq�*�����?S�&?�R�>�H�.�D�iʾ�z��
��>�I�ӡO�6���ت/�E�%��w��X��>"Ԩ���ξ��2�G���w����B�iyr���>��N?v��?��f��\���P����?��Y�?��g?~`�>��?�3?&ϙ�Zk���}�|��=P�l?�b�?8��?>T#;�~�<��?Dn?�ן?���?7ց?)�νY�>!酽�M >����Wk5>��=��=�k/>��>�*?�C?P�߽����t	�8��������<�,>�^�>?[{>�%�=F����zx=;��=�e>�I�>٨7>z[Z>ڣ>�m�>�@}����<�'?���=�r�>J8?p�>��<>�`�H��Ӕ�v�V�o�����z�,]?��7�<���Nv�; ��<]?��¿wG�?��>�=��~?������/4�>�>�>]�=]K�>p��>Q)�>��?�W�>��j>�ɢ>�..>��e�P�=��0�ӣ� d�{�9��d���d<פ��4`>_#��������$����x#��r`�'}��U�����o�?�&����D�Yu%�{��<�?Y��>��_?y�+�����or�eD�>��>��
�`!����@[侭�?|��?�:c>��>d�W?f�?j�1��3�'uZ���u�$(A�be���`�፿���9�
����\�_?��x?xA?E-�<*<z>��?�%��Տ�x%�>l/��%;��6<=�,�>v'��u�`�-�Ӿ\�þW6��IF><�o?�$�?�Y?PPV�&�U�z��>��f?=�H?
��?�J?/gZ?[o�;��?s	�=T��>$&�>Vj5?; ?#�?��>���=A1�=R��=��A'���hQ��9��o�e�ѩ=]>���<��u==���0����M=��3����*���Y��&�F���	>6+(>}>�>��]?�v�>i��>�N8?�{��8��[���Q.?bk2=
I���ы��@����!�>(�j?��?�Y?@a>FB�KlB�S�>@K�>I%>��\>�q�>���RF�@#�=/>�>a7�=��]�m'����	�2���9�<�;>v��>]8�>�խ�6�>m����蜾���=gY{��ۅ�M.�ǒ�/g��Z�v# ?�bO?χ???ae=����!?���Uh��#E?�?�%?�ӄ?oh>�"\��	��v�F)��7�>󄢾�R\����ZѺ�T�3��=a�>�Q��Z��8�>�8=�tC�?P����/�T�۾�2�F��k��>�Q���ؾj ��g5>�(>s[����9�T%��K^��d}?W�K�N��^\N�t�����=HT�>��>u��=?z�ٝ3��=����=e�>�6�=L���2�t$f��X��ߤ>�??�z`?��o?')���W��<p�er㾕՘�WRܻ�-�>D��>o9�>���>���=��=l������L���>��> 8���P���3�{�@�M��+�Y>��1?��=��?�?�?O�L?��?� J?��Z?`҄>�:��ǻ��?&?*��?�;�=cԽ��T���8��#F����>�)?Z�B����>ʄ?R�?��&?]xQ?�?��>3� �vC@���>uM�>��W�#d����_>6�J?ǹ�>�>Y?�҃?5>>��5��颾�h����=>R�2?�.#?$�?ﶸ>g�>��@�=���>/$c?4<�?Ep?��=L�?#z2>|��>�o�=���>���>�?�DO?��s?��J?�k�>�ڋ<?Ӭ������t���I�j+�;-uG<6}y=�����p�����<��;0m��O�|�G���D�{܋�h��;���>��r>����0> %ž����wIA>Ӯ���ڛ�։����9�̸=+�>E�?ѿ�>y$�O��=9��>H��>����'?�?y)?_�#;�}b�C�ھ\SK����>ͪA?\��=%�l��z��x�u��h=��m?ܸ^?��V�������b?�]?ig�=�O�þy�b�I��}�O?v�
?�G���>&�~?��q?���>��e�':n�F���Cb�9�j��ж=wq�>�W���d��>�>��7?�M�>>�b>�'�=rt۾��w�Bq��p?��?��?���?�**>��n�D4��]㍿=na?��>�,���T%?���\�˾����Uy����׾����԰��ȝ��詾�:"��1�����NG�=�?��o?��i?�Z?���T:Y��r]��{��(S�<������E�~�J��_F�Zzp�g��zT�G(��"gg=V:�)�:�\ʲ?�#3?����� ?𛟾^쭾z��(X>
���*�]�5q�=H����i�[
�=��냌��8��l�?pQ�>��>�P?�Ol��/�"4E��69��o��=%S>�U�>�]]>���>��:���)���U� Q��Ș��3�ؼ�w>>c?�{L?�o?aY �=�,��&���<!���*�Щ����F>�>�!�>��_�f��ڰ%���=�S\q�EW�8]��ef�KP\=��.?��x>���>���?��?>�������w�g�1��S!<N��>m�d?���>�̆>��ʽ���ư�>�6m?r��>��>�胾��Qv�Km��$�>Aؠ>���>RAk>2.���\��D��cr��*|:��� >yog?*u����^�%�>�:P?/֨���<5��>�ᚽ�� �����&���>'u?��=��7>E þ�����{������O)?�L?{咾�*�F8~>4%"?.��>l,�>�0�?�+�>!oþ��H�N�?=�^?�AJ?�SA?IK�>��=���?Ƚ��&�k�,=���>��Z>� m=�}�=
���o\��r���D=�p�=R�μsN��[�<>j��]K<V��<��3>�ǿT���n��@�l������u��4��!⠾	�=h�U޾x�f��N��-;</���|�)�e���4�o]�?dD�?���������qDw�k���>n���F�F���������]�k=ž��ǾL#%�	j�ձF�<�c�e
0?9뭾�ȿ4ӣ�ͽ	��2?��?L�p?�<���8�1��=�m�<:e��l�����pϿ���q�^?�1�>���6�?=���>�P�>��>>/P>�ڈ<�MI�,�[�>߼9?�N�>��������I���#�=;g�?��	@yA?��(��쾾BW=#��>�	?��?>�71��8�T���a�>�3�?c�?HL=��W��K
��ae?�<��F��໅*�=��=o�=����J>�D�>�f��zA���ܽŻ4>˵�>E�$���#�^���<��]>ȇս���5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=����������%�zG+�׍>�:�=P�h=��Y�꽭i�=�L��' ��=�ܽ��=�:>]6�>@�>�� >[Ob>�[a?�~v?u�>�i1�=�6���q�����~�Ц��N�v��+��=��������ž��������*�:#��{8��B>�)U�u�� f��Y���B���?B�=j����6;��)��tG���p����h�����</Ծ��-���i�K�?��>?OɈ�UC��]���_�l�ʽ��M?���P}��������>ޡ�;Ó�=���>��D=�m�Y�7��>a�po1?V+?�л�U��a�	>�+��e�=��/?$$?��=��>Z�!?��S�?l	�6>��>s^�>���>��0>�l���v��	#?�CW??ʽ���ڂ>P{��E����4=p�=<�-�������X>�)�<)��O��A��X�u<Q	W?�|�>7�(�_������1Q�i�p=��w?��?7��>��m?��B?�S`<���~�R����[Y=�#Y?8j?�>����о�[��ƨ3?�c??iN>S�e��i羾�,��I ���?S'i?�z?-N��Y�{��ِ�,��Q�5?
�v?(h^�5^�����b>W�B��>+M�>9��>��9�%B�>+�>?��"�O��㴿�l4����?�@Fz�?7sD<�F �/�=lH?[�>�O��ƾuz��4�����n=g��>0֧�Mcv�����X,�fz8??���>�l�������>���Gح? ��?�̾�M�=�;���U�Qj��4=�j�=�4Ľ]�ýǤ��Lz<��4Ѿ����0Ǿ�������>H�@Ceɽ\��>��?��׿�ο䉿����=sl���?�è>	�%�e����Q�1��p%P��H�sш�=z�>��>tf���V��g�{�"�:�������>ܵ����>��R��赾B���)<Xp�>��>��>6��&��ֳ�?����z οP�������W?觟?�n�?j`?Ƀ[<e$v�Õz�̭ٻ�]G?s?ԧY?n(�L�[���0���n?n־�Q��:3��zD��A�<�?),?D�ھǯ=H$=9E�>��#<(I�����t��A��o�?/��? T߾���>	-�?DK?^�־Xߜ�����{b�^�����>�v�>�����7�h�(�J�dK?��\?�>��]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?' �>{�?z��=�W�>Q��=�Ӱ�ŧ*�ʑ#>[�=�]@�?.�M?�;�>���=�$9��$/�ZcF��:R����C�S�>n�a?\�L?�b>G��s2�H!�"eͽ�L1� �輐W@�l�,�IN߽(5>�>>E'>�*E��(Ӿf?]��`ؿ�W��
)��3?��>�k?}!���r�;����^?�>d����M��	��D�?�-�?�?�f׾����z>)]�>�5�>u�ս=�4톾/�5>6XB?.���;����o�&��>���?��@�®?�`h��	?��P��`~����
7����=��7?�,�0�z>��>��=�ov�����R�s���>�A�?�z�?���>ɬl?;o���B��1=�L�>o�k?�r?-p�W�q�B>��?�������K��f?9�
@u@��^?9�I�ӿ�����@!��L�8>�P�=$�>�%O��Ȋ=-F������$K��vB�>v�>'{�>�\�>~�>V1>��5>D=����֘��q����������Y��?��;?۾`���
���ľG���ӭ6��N�e��;1ۙ��42��cۼ{f�=�T_?�-W?�]t?ɋ?7C ��g_>(��=1`���B��q=a�e>��/?M?�G$?%I=�탾�g]�O~��|��T}l�H߻>y�G>�b�>�9�>a��>_��t�y>\�>$˃>x�=��o=l��=%��=���>���>2� ?��>�x<>ъ>;ִ�-��5�h��	w���˽��?[z���J�� ��O��u���r�=hP.?�(>���n@п�����;H?�J������+��>P�0?�\W?k">F̰��iU���>N����j��� >�� ���l���)�k�P>��?
�f>�qv>�3�?8�H�O�g���A�|>��6?�C���N<��tv��DH��ݾ�L>�Ƽ>(�b������F�~���h�#�p=��:?"?�ͷ�~1����v����9�R>n�]>Z=���=�=M>�9Z�{ý�HE�	?2=>�=?;[>�?6�=QpZ���i>�*�p����?�&�>Hd�>�K?x�_?Z��<�B侊���`I���	νCz?�?��>�o�EhC>�?�Ω>36>b8�=)�I�V������=$�!����ͯ�O�=�ˈ�ɷ�=��>*=�m<����~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ��>?��{���F����v��t%=Ő�>�9H?���]<��?���?�?&��z��7�ȿ�Aw����>U��?~I�?�Jm�բ����>�!��>�f�?�+X?��v>N�׾_\�1�>��A?��P?U��>D���""�ޮ?f��?~P�?-�c>��?�0|?�?�u��Ԃ��oᶿ����<=�W�{�>��=�W��^wM�1Ԋ�ǈ���`��!�w�>F�M=`��>eG��-��#+=?�߽nn��q먽��>��6>���=&��>h2�>��>+��>4X6��I ��+p�~Q��m�K?S��?����1n�ZK�<B��=��^�A&?J4?�V[�Q�Ͼ�ר>h�\?�?3[?�e�>>��C>��<迿�}��7��<#�K>`4�>bH�>#���FK>��Ծr5D��o�>gЗ>\����?ھL-���Z��8B�>�e!?ѓ�>�Ү=�%?�?��|>�s�>�#E��?���I��>s��>u ?��z?1�?+|����y���K��>D]���>=[?��?�%=\����բ��F �5e׾l��>d�x?4(??.f>��1?��{?w`-?�=?r>��T�1�վ��=>�? ?��!?�(��A��G&�0N��^?^?S��>�ǒ��&սm�м���L�����?Q\?x&?]��/a���¾�1�<,R#���]�ٱ�;�=E�C�>�}>���8��=S�>à�=<ym���6�d<�g�=�~�>>��=|'7�7���B-?�Rü��}�J�=s���H�e9{>r�c>Y��C^W?�6�|st�kŭ��t���[m���?�X�?�#�?)r��H�g�=?���?��?��>bߤ���ھ�]⾏%��A�������=�0�>����jXھ�Z��*ڦ�)р�������Լ��>?�c�>^��>Od+?���>�=?>��<��n��o�r��',������T�T)D��,>�:����<ʽ�3I=��ɾH�B��>FI4=T�=Q��>Cʞ>�����>۫�=��o>a��=�S�>ܥ?M�G>��{>d� >�����ER?����Q�'����[���|*B?�od?ME�>��i�b������5{?+�??j�?��u>�h�D9+��h?�8�>���=_
?��:=t^�=��<�K�����銇�Ӷ�_��>\׽q:��M��Bf��j
?�/?{���I�̾�׽8r��g��=��?�1?�#���?���u�AKT�)8L�[���1�F�?Օ��\)��q����iҀ��Ɂ��v%��Q�<�X"?�Z�?�	�����-��دX��~:�~�`>�0�>�&j>(��>3�#><����7��qc��93��w�xz�>z�t?9��>�Q?�'@?�S?��N?Z��>��>�ٴ��d�>�˪:R�>�n�>��7?�0?�(-?�M?�,?�e>א��~���Z�˾�,?�u?�D?Ⱥ?9�>�<����y�$}=C�1;�r��nHx����=��:=����������=��a>&�?p5��2�J��Ղ�=K?� ?~�>I@N�?���X�e>>��>�5�>��f>(S����{�=��� ?�Ȇ?WP�֩���=��f=��4�8�<'=�=Й�.��=�Ƽ�J���J�Ţ��2<��<��O��=��<�<�<�7�>w?%��>���>ä���������٩=�7Z>�YE>�>��־�Њ�h$���f��Hp>���?���?��I=���=��=�棾D�ž����{���6=��?�s#?2	T?�?�Q;?��$?�E>>���z��Z*��l���`�?"�,?�K�>a���ξI���N�1�G�?ov?�^����~M*�������ѽ��>�0���}�����ͼC����;���۫��c��?�ʝ?w��57�c(��_�������@?�r�>
J�>-Z�>��)��Cf�`N���G>M��>��Q?E��>�|
?	�J?�x?Z�=�����������?��>;�5?�N�?�?c�?��s?f�?V���.���]��T*��� �T�����>���>��>�!�>��C>)��=%�B=���0����=L�<��?}is>}{>�5�>[gͼ��G?\��>�]��ɒ����X샾�+<���u?i��?��+?�n= p���E��Z��d�>%\�?���?�5*?RS�T��=B�ռr���^�q��'�>Nù>� �>6��=z�E=�*>���>˅�>GE�jY��g8��L�&?�F?��=�ƿ5�q���p��Η�Guf< 𒾸e��ꔽW[�6��=麘���X�����[������s��u䵾������{����>=��=��=���=k8�<�Gɼ�T�<S�J=��<n-=�p��Xl<�9�&�ϻ������SH\<a�I=����O˾��}?�YI?R�+?��C?d�z>�8>�\5�w�>����A?��U>��R��b���Z;�J���A֔��gؾBu׾i�c�x���L�>� L�K�>63>۔�=+׉<���=�et=���=��l�_.=[��=��=7�=���=jO>�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�8>\�>��R�w|1���\�v c���Y�p�!?�,;��-̾�U�>�e�=#i߾��ƾd,=�6>մb=;���\��e�=fSz�X�<=�Rl=�ŉ>��C>Y�=н��8>�=Z�H=S�=F]O>䇠���7�k',��4=���=��b>��%>;r�>��?L�1?��e?�~�>uT\��Oվ	O���>���=�r�>8H�=��2>�[�>�5?�JA?�vH??b�>L�n=�ع>JJ�>�P-���n����@b����=�?]s�?�2�>}W+<�hF�-��~�<�{�ѽ@�?+�/?7�?n#�>(#��Ϳ{|1�B�M���><s,>���b�%7��1ؽ!bs�񔘾j��>5�??vb?f�1?��?��>�a'>��>�܊=#>�$��;S/=co|>��>�&E�6=�=���<��'���
6d���e�~���Q�=�a�<蓔<��s>���>���>踰>6م>*�F�ebb>B�1>.�K��T\�ٛ�R��d��R����/�]��O`>rq�>F�>[���i� ?���=�/�=��?:��?z]->��j���J�Jԧ����>W��g�Y>��c����6.��l�.;W�����l��>mt�>���>��g>��*�@�=��̀=�Wܾ��5�5�>t�����!�� �p��@������ �i�"�"���C?����`�=�~?�BJ?Sǎ?[��>�,���پ.0>ǲ����=0���o�
��b�?�g'?��>���(E�I�Ⱦ�:ǽ:�>��N��EP���&�/�T �|����>���0Nо�#2�t���᏿�}B�v�ǋ�>��P?b��?.@a�#I���L��e��V���f?�ei?u��>!E?_>?�Í����l����ѵ=�;o?���?�.�?i^>��=@�l=N?I�?�p�?�^�?q.�?�ac�!�>���;5�$>	V��>��Q>3��=3��=�N?��?�X�>{ӽ���A�׾�Z�4�9�_=�=|�|>8ť>�>l�>�Aa<�ь=%B~>��>')�>�pN>kU�>�n�>+#~�5��Q�)?x6>�Ê>��6?>�p>�u5>M7������D֖��W�cb���ؽ�_�	�d< ?���ڽA1����>�sǿ�d�?,�>\�2�h?�|��@���>�[�>��=���>OM>{�$>AW�>���>�^�>�R�=Sg >HLo���=��>�jE1�Y�p���9��ި��>����Ѽ-2վj�;pD��褾�`�y,p��p��,]�w���3o�?�3��!�@�a�1�ո~�& ?�>W	j?O��sϽ�|��>��>��e>�x���������WѾŤ~?�@�Dc>#"�>��W?6�?ć1��2��~Z�G�u�zA�{e�L�`��؍�ܝ��ڞ
��$����_?X�x?XmA?�0�<%z>R��?�%�Z⏾��>0
/�\;��g<==�>dC����`�κӾ��þn�_�E>�to?� �?�R?�:V���j�W`>� A?��4?�Mx?t�8?�\B?� �
?�M?>YN?��>�&1?�02?�	?�T6>L>���</� =�Q�������?��2|ڽ�9��H=��h=�k�{�<�=P�=��������;�)�t}D=5O=b�=Xa�=�Ц>2�]?��>��>��7?R����8��Ѯ���.?��2=�ځ���������Ţ�$>0kj?R��?Z?��b>��A��5B�b�>�Z�>2%>�M]>�0�>��F����=ڂ>g�>h�=��S������9
�*���)�<KD>���>u��>z��=ʱ>G|��1P���(=�8p�a5e���T� ��n�0a ��>ѡO?��'?d�c���ݾ�3�G�\�]O)?1?��/?(J^?���>־ݾ�#��v� _���ۭ>��M�4�N��i���0��`:f�S�%=��h>)4�8s��g�>��S���G2h�x���۬�&���B�2��>�ʭ����ؽ���>9�M>g�*�́���wr���� �v?� n��4��:����V�=��>��>��">�Cؽ|?�<�v�#��>�
?
�Q�L�5!����;���	�C�>8�?�c?��m?�3ܾJzu�Ŋj��������@k��N�	?�A�>�<$?�T�>t��=�����o���0��߲>�1�>��F�]g�p����N�4v ����<��9?�@ܻ�?
��?	��>^�M?�H?%�3?O4�:z.��,��A&?���?��=��Խ_�T�� 9��F����>9�)?��B�l��>R�?�?�&?��Q?4�?��>"� �D@�+��>�Y�>��W�:b���_>��J?���>�<Y?�Ӄ?��=>f�5�뢾ة��Q�=`>=�2?6#?�?��>��>�����=��>��e?>ā?�4n?A>�>�P>l��>�=h%�>��>\?��K?_�o?�M?��>��;,����ΐ�;bǼ�.:25�0̊<,s�=��>k�-c�����<��#;�+��0��;ݢ
�Φ!��D�f3Y80��>(�q>��z�0> �ž�s����B>�t���)���l����4�0��=�`>)�?���>],%�K�=�R�>>�>���<�'?�8?�;?��;��a��۾�EL����>1hB?u��=��l�������u��Kh=j�m?�R^?��W�Y���
�b?�]?�d��=���þ��b����Y�O?��
?p�G���>��~?��q?3��>m�e�O3n�����Eb���j��Ͷ=l�>\�M�d�/=�>��7?�K�>j�b>�3�=y۾D�w��d���?\�?�?���?$*>��n��3࿞6��<��8 ^?���>�ߦ�A�"?����	оC�������c��Ԉ���O��ݸ$��򃾽P׽��=M�?��r?@:q?~{_?�� ���c��^����@}V�c�����E�� E�0�C�s�n����������XH=1IR�s>��F�?9�7?AƁ�&�?����Ȝ��W:��>' ��
n(�Qa>M�q	���P�=i���az�{�����?v�>�$�><�(?=s���Q��Y��E.�O2���?�>��>�g�>��>l��=�|ĽTs?�B ���������"v>�~c?��K?U�n?�� ���0�����2�!��0������A>�>��>nvX����&��J>���r�����w����	���~=�42?;�>���>$�?=�?E�	��%��[Ax���1��`�<���>A�h?�h�>��>j�ͽa� ����>��l?M��>��>a��0I!�T�{���ʽk��>��>��>�o>��,��%\�v_�����m9����=�h?Z����`���>&R?�h�:��J<�n�>�hw��!�����'�-�>0e?.l�=]�;>ۈž��/�{�z+���P)?I=?�ʒ���*�"a~>�"?]j�>R'�>(�?L�>�VþP@���?�^?r8J?�HA??*�>��=���eVȽ�&�W�-=��>�[>+m=���=���b\�R�<{E=4r�=�ͼ&B���,<-�����O<^��<�3>��ܿ�	1���۾����8�wL���m��3!�,�j�ýy���hB��p�������������1�l�r��e���?��? ����.��'ŗ��fv����3Ӎ>H�`�n��Ƈ��HϽ���b;Ӽ����\-U�"�l���j��3?%Mؾ�#ȿ�ɠ��@���?�G"?�ch?adо�
���8���%>�NR>�������$����?ȿ���vn?HG�>$������=�s�>Ș>_��==�o=r����V̾�Ks����>��-?	,�>�����K��U���G6Y����?E
@�I?+85��%�j���&>��>���>4 <�L�ʾ�e�:9�>�:�?-Ǖ?~`>�T�}E����Y?F(���P�u�<d_���>�~a�-h��!8>��>~S&=��
��g���=3"�>do��aN���վ߽<Y2=ǚ��
�>5Մ?,{\��f���/��T��U>��T?�*�>T:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=j6�։��{���&V�~��=[��>b�>Â,������O��I��W��=���HE���-��zL��>ym�=�yüSI��M7C��?�=�܅��W���I$�.��=��Z>"��>� ?�>T�> �v?��?�>�>� �������վ��&���>����i�
�1;���ݾ&���_��D���7��b�!Ѿ�B�P��=s/Q��7���3�n�Z�C=���?c�>Ĺ�.)C����?�̾[��Q�лq���:��*-��dk�]��?��>?���R�Au��������G?C��{o�Κ��l>Ә�/e=wɞ>^y�=�쾬5�b�V���0?�?��e�Nm�U��>��^��Z�=s�*?���>�HX>�u�>�7?ڷ���j��9O>��>��>��?���>�ʼ�V_u���?Yxj?!��E7���>Z�������.���h7_>�b'�U����S>��>���A�;�G�����~S?|/>G�"� ��䋾��d�>Ħl?"��>к�>C��?f�)?%�Ƚm���~I�QX���=�8r?�j?���=�jA<������W`]?�	x?��=�U����	���޾(�'��b�>/�Q?���>J� =M2D��T��5�	��?��v?�r^�sq�����?�V��0�> ^�>1��>�9�Bo�>.�>?P#�\G������[Y4�3��?�@��?�=<z$�Y��=9?lH�>+�O�4/ƾ���� @q=�+�>�����gv�6���g,��8?)��?B��>.���������=�J���W�?�D�?{�����<6���Zi��- ����<K��=?���L	��B�7�<ƾ�e	��<���j��Lۆ>��@��ݽG��>Yv<�VZ��Ͽ�΅�s"ʾ�pn���?�B�>�H˽t5����h���t���G�pDH�b⋾n>s>�3[> B����}p��z �oZs�&\>8X�&Y�>��׽i��3�'�==Y�>+?��y>��޽�{a�?A��hѿ<���7���E?�g�?�s?L?�?�=��q���Y��ˉ=ԆP?�)^?l=1?J>���;Z�؆��{.i?�����M�SP.���B��������>�s?���rU�<�I�=��>���=�R�Kÿ擰��d�1�?=q�?/(�s[�>�s�?^~?<dӾM����վ��n���>�B'>��Ҿ�AY�L��b�Z�h�>P�N?�%x>RZ�6�_?�a�v�p���-���ƽsۡ>J�0�Jg\�SL�����IXe�����@y����?4^�?V�?1��� #��5%?��>ƞ��H9Ǿc
�<L��>�(�>�)N>�E_�3�u>~��:��h	>���?�~�?-j?�������1V>��}?
(�>��?N%�=Yi�>���=�ϰ�Ѱ)�L~#>�M�==���?9�M?L�>Ka�=��8��/��DF�vR�|����C���>��a?��L?�Eb>�ĸ��{2�!�/νM�1�����@�K/��߽w;5>�U=>��>��D���ҾR�?���m�ؿ3`���'��	4?+��>0?F��4�t�����2_?�]�>	=�n*��!(��wi�藫?�@�?[�?E�׾A+ʼ��>��>R'�>�5սT柽�����7>��B?JL��K����o��
�>o��?�@�ծ?��h��	?�!�iO���_~����7�]��= �7?U/���z>%��>�=�ov�^���T�s�K��>�@�?{�?��>��l?�|o��B�j�1=,P�>%�k?4q?�Vp�󾂧B>��?ô������J�kf?��
@�t@�^?9��ٿ�����^�����h�==��=��J>���ٚ�=�{�;�^ػ+��>��>��p>�!�>�y>.�]>�8>�˄�C#�Z���c�����D������ �ɣf�;� �k���~_	��g��(ž����v���-����V9�N��U��r�k=4%i?��`?�Ԁ?��?~<%=�؍>����5={=k�R�3�'�W�%>�%?�:J?{L4?6A�=~��o�\�I~�񾲾�k�=V�>�>�I�>�!�>���>�M=�ef>^M�>.ف><��=���=�m�<8?>��>�>���>X��>=>:B>ᴿ�,����h�P�v�iKʽTҢ?Aǜ��gJ�%��*3��֔��m��=��-?sn>�䑿@п�᭿6H?�S����v-,���>D�0?DIW?�>���gX��>����Qj���=����l���)���O>�?��f>.�t>��3�6g8���P�Gq���f|>�"6?$Ͷ��9���u��H�z4ݾ��M>뱾>^vD��]�K������Oi�E�z=~q:?~x?�=��ް�su�!���}R>V�[>/�=m��=�vM>$�c�
|ǽH���.=D�=��^>��?���=�U=۰y>m
�Wp�=��>a˄>��#>��C?^_C?85��W�2͕�l�O�>�ͻ>��>��>zE�F��=m�>|; >zp�=s=�w7�&Id��h�=W��<�ℾI8���B�;D��4`>���=O�ý��P��=�~?��刿��0t���kD?�*?;��=�F<΀"�|���bI��!�?I�@�k�?��	���V���?;>�?�����=�|�>�ԫ>%ξ=�L���?��Ž�¢���	�t,#��R�?Y�?� 0�ˋ��l��6>[%?�Ӿby�>����I��f
����u��B"=���>�5H?W;��(�O��X=��z
??cL򾝟���ȿjxv��*�>���?C�?��m�~=��	�?��)�>�w�?LwY?P(j>\۾�WZ��>ҽ@?��Q?i=�>9�/�'���?:۶?կ�?��D>F��?�q?�t�>ćA��s&��&�������sW=VN<Z��>�=�ʾ��G������S���nh����xBL>»,=�B�>�"��о�,�=�㎽�_��,����>�i>O>��>�S ?�>�>���>�G<0塽��V�D�����K?r�?r����m�-K�<2	�=K�_���?ǈ4?�[��yϾz��>#�\?���?|4[?'ߔ>8��>.���ۿ��w�����<"pL>{��>���>������L>��Ծ�F�	Y�>C��>A����ھ꜂��껮
�>�v!?I[�>�C�=6� ?�
?U�U>[~�>A�@���������>�>���>	�>�?��?�C���%�����k���!]�b�>I�o?��?w�q=�ԋ����s�I��c��1�R>+ƕ?8Hd?+�\>L?���?��3?_eJ?6��=^�:�����n>=�> �!?�Y�~�A��Q&��Z��p?�K?���>�[���Uս�0׼5���$�� ?3\?y6&?>���/a��0þ�/�<�(�Q�M����;��D���>b�>�����ϴ=+�>E��=;m�66���^<�)�=�x�>���=��7�f쌽=,?�J��Ѓ�9��=$�r��vD���>cqL>���%�^?�h=�&�{���jx���;U�d�?��?j�?������h��'=?J�?p�?�8�>"!��az޾=���w���x������>���>��l�����������I��]9ƽ=g��X5?	G?b�?5&1?���>�F�>��.�D@�
�<�����T�ՅT�K�=����1M�N��lZ�gȈ�ؐɾ�Y��ѸN>W*>r�I>��?���>B�=�w�>�9d��Hʽ�fM>���>���>3�X>�V�>�ں>���������GR?���U�'���x����A?`{d?m�>`�f�zn���E�O�?�k�?_]�?D~u>Dh�f+�@�?=d�>���3
?��7=���|�<�O��t���J��=�zَ>��ս�:�TM�of��=
?[?|�� b̾�Yֽ7|��D�~=���?D�(?˶(�`;P��o���W�Z~R�9���i�x>���!%���p�Hj���
���ჿ3�'�� =*?c�?J���`�]���I�j��<��Mj>
��>V/�>W�>
-J>I[���0�4�]��Z'�^�����>�H{?x�>��Q?�_C?i�W?�O?a��>���>L)�����>(6�ޏ>�,�>ȵ1?�*?��2?dY?��4?��Q>��_E ���˾�q?k�?(�?��> �?�Jr�4��P;<��&�"bz��-A����={��=�c�y~���o=ۙX>N�?
6�@#�A*��
"Y>�`?�~�>�Q�>�҂�M!�L�>���>��>0�F>����c���*?��?�Y���<��?>$ >��*=zV	=���=�=8l�=�%�<FiV��	=Qf�='`�=i��<6�=��=.iJ�b�B=m��>2?7�>�P�>�؄��<��;��gb�=��U>�S>c�>�vؾ����՗��f��t>*�?���?��\=x
�=��=&��/nž6������G�%=r[?�"?��R?Ē?r�=?�?$?��>V����+���?����?4L,?�ӏ>�B�A˾٨�x43�z?�q?��`��x�hE)�����ѵϽL>&�/��~�����\D�덄� ��������?謝?>@<�87��龟.��	��*C?}�>c~�>�}�>C*�ܳg��e��9>��>�=R?k��>���>��?�~N?�7E��ˍ�����A�x�a= ?p���-A	?Rf�?���?�Ƈ?ϪH?�>��	�����6�Ur��P���ʤ���=��j>�>���>��=/��=���=�2��7�t��<��=�A�>\$�=�_�>0��>��<��G?���>�_�����(���,؃��]<�֝u?}��?��+?�=�v���E��;���3�>Lc�?M��?�?*?ÊS����=�ּ>㶾�r��:�>:�>��>po�=�,F=O�>��>�>�D�2g�3g8���L�w�?^F?S��=mƿKq�q��
����f< ͒���d�ݺ��w[��6�=�������쩾��[��������3����v���{���>9��=���=��=:��<iɼ�V�<�SG=�.�<�7=�>m�<�s<�8���ǻㆈ�j�u-Q<��F=dz�.�ƾ�l}?�1H?�,?~)B?��>�� >�d��>��>��o�y�?�WL>�����¾��;�M���×��>׾=پ�a_����� >��Xp>0>�W�=.��<��=ڷo=<M�=����m*=��=��=���=Q��=�6'>ċ>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>G�7>y	>��R�u�1�֋\�v�b�ULZ�;�!?b9;��'̾�U�>c�=L/߾��ƾU�-=�H6>�a=����2\�ƙ=��z�X�;=��k=z�>�D>�:�=P8��Y��=�#J=�\�=��O>7��� 8�R,�4=U�=g�b>�&>�t�>?�L0?C,d?��>�:m��CϾ+z����>/P�=�װ>�a�=P�A>��>�7?�SD?�xK?Ym�>ڽ�=�$�>T�>	�,�#n�%�往-��jɾ<���?��?�|�>��j<h{@���h
>��Cƽ�'?��0?D�?�m�>H���+�t(�L�6�U�h�V�<�>�=m���߄�������p���a3>�v�>)3�>+�>�s�>mV>��^>� �>��>�E:�ĉ=gH��ϣ=&����=8�'���=�y�e���3w��C���|H޼�;��=��;E.j<�4>⽣>��>�Ӏ>��Y>�����0�=����ch��I��<�����E�ʸ{�:��-�2��Ծ��>FHs>��=�Ԓ�t-?=�J>&�,>ΐ�?+�n?��=5儾nA�-p������`�Ӿ�^��<��=Ñ3�G�7���9�6m��f׾y�>��>��>��g>��+��z?��tk=��ܾ�L5����>�C����!�Yc�~�q�|B��k����\g��;)E?� ��Xh�=�Q~?]HG?a��?��>�8��^�׾Y�$>ׂ����<���u�l����?UD&?��>+��`�D��˾�Ž�P��>9I��O��v��)0�(�������>�ީ���Ͼ"�2��<���Ǐ���B���s�Y��>�|O?���?�d��L���yO��E��=��\^?�#h?�^�>,�?�&?�󜽱�뾂~�d{�=�m?�?�?SH�?g�>d�=�ro=�;
?�F?���? ג?�?V�.���>9���u�=2�����=�\0>�6>;�>DT)?���>��>c�޽�Z����ξkF����Q!=�>�q�>ȕ�>eq�>�>���=g��=n�S>(�>=h�>��l>(�>X��>�2��v���
�? ID>�ݨ>0YD?���>�c>1^���!�2�{�8vZ�kr��ݛʽ3BG����=��;���<��x����>g�ĿZ��?�4�>�QG��1?����l<p�>�X�>Rٳ=\��>s�>" �>���>�c�>�>o�'>�K>�ϼ�؝3>�'����Ճ6���?�λӾ�yB>����Z%����N��[ET�?������(d���~�n\-�a{<nK�?{5�j�|�@�B><��{�>���>�RE?���􊟽�
a>t� ?S!�>��ݾ�ː�Ʊ�������?���?6c>�!�>)�W?H�?̃1�"3��sZ�X�u�?%A�fe�.�`�%ߍ�I�����
�W����_?��x?�rA?��<-z>���?]�%��ڏ�m$�>�/�W!;��K<=� �>'���`��Ӿk�þ�6��/F>��o?�"�?nY?�QV�]G���x>f�H?>9?wI{?��9?�IM?�5�_E!?��*>���>���>W�0?"(.?|w?USL>BV>�,;t��<^6��<τ�u���0?
��m����F=1�= `={��(��=��?=��C���l7B�Gy9�v�	=$�=�:�=+�=�ȥ>��]?:��>É�>x�7?����8�����d�,?4K=M̓��f��󥥾x���j�>t�g?���?~�W?�^>�D��i>���>��>)�'>I�]>8�>+f��O�j�=	�>��>�f�=�Fi�a����8��Ґ�rA=ٺ>���>�U�>��F��>A┾6!��z�=K���Ԍ-��1��0-��g/B����>S�M?�&?ђ�����w�;��\�Ȃ;?�KI?I+3?��}?W�>����+B-�~�y�����S�3>U!����+��������C��[l=}>	8$��A�o�.>�>��A��z��S�J��M��w��E�e>�I�����\�����>ߗ]>c;�������Dn���vi?T�j�vj���w�v��='��>4��>14>���K�4��)��c��>d��>����!�������Y�W�{�c>KD?�tY?�pK?�0k�Q�a�ta�x%�'���;=A>v<�>���>�g!?�N�>BP1<�N�q�1�m�*���j���>�}�>k-E�y�L�WXʾ>:
��?۾��N<��?�[>�F�>F`?Vt?��C?��O?��B?��> J����� �%?1h�?H��=�ֽ]pU��w9�bnF��*�>Od)? 8@���>�?J??��&?�uQ?x�?{]>|N�L~@�g�>eϊ>%�W�Iү���^>�xI?��>�X?S�?��:>_
5��k��=������=��#>F	3?�"?0p?�s�>���>�ß�6x�=jx�>�U`?m��?�jl?xx�=�?H<>D��> >��>�=�>�?��J?�@l?VfF?���>�"<�I����ao����[��9���W�V��=�$6�ҟ��B���=�
M<E] �@�a��]��o���*�kL�<�S�>�Xn>] ���0>ԛǾ�ʌ�ۣD>�ㄼ�{��o�����,���=�s|>f\?�6�>�j%�䛎=�"�>��>���&?�?��?p^;��a�Wؾ��H�Uv�>�AB?@i�=K�l�K<����t�x=�?m?�t^?	�U��m����b?��]?g��=�#�þ�b���M�O?��
?^�G��>��~?��q?t��>��e��7n�P��WDb���j��Ѷ=�q�>�X��d��>�>�7?(N�>��b>-1�=nv۾A�w��o���?��?b�?���?�)*>;�n��3࿟�ܾO����QG?ȣ�>m�����;?Y!��ʤ����5�ξVR	���ʾP]��.&��̽ʾ�s۽������'���>��?g�Y?��}?��_?��ξL�m��V_��V���S?�凢�(i�t1�)lD�#E'�f�k��K쾩"����H>V ~�j�>�*F�?QX*?�2�-.�>7����xо{�+>`y���N!��@�=֒��L�=A�w=0n�EO3��6���? A�>	��>�c:?`\���<��%/��k7�=��u_;>â>m�>�~�>-�o;v�0�5>޽�`˾'�~�k���=8b>4�e?��K?ߘs?�ӷ���)�
��#�0�z��v/>tY�=��v>WS��.	��*� d<��u���������߼�=P:?'�|>6s�>։�?� ?e����]C~��65����n�>��Y?� �>��>àĽ.����>��l?p��>d�>�e���F!���{�"�ʽY�>}ϭ>���>�o>��,��(\��a���}���9���=ëh?�����`��؅>�R?Lv�:%K<eq�>Zw�)�!�6���'��>Vx?�ު=�p;>�jž���{�l<��£)?�{?M����u*���~>�?"?7h�>?1�>�?���>�¾���;�t?��\?�`I?Ŷ@?��>,!=tF��Řɽ1�%�K�.=���>4'[>�Tf=�r�=K���]��H!���5=�	�=o�Ƽ-+����<�x����<I=߅4>��࿱W)��7Ѿ��1��ƾ<nҾ�ء�S-U�����U��A���f�Ծ�����l���"=�/ֽ[&�˯��H�����?b��?��Ⱦ���M���`�V0��R&>��I�P]Y=�?_�6��i���u���p�*�-���~���P�3�d��6?�V���ֿ����հ�@�?_�?u�p?3`���Z���5��k>>�(�>�m�	���u������Tؾ��Q?��>j�����=`^?aJ�>G�=4lU>v��=�b��R� ����>�Fo?$ӯ>�����=��S฿��9Z�?Tn@FVB?'!+�<i���y�<���>�?<�?>gF4�+<��l��f��>s�?��?^��=%X��a%�_c?sߔ� G�'1`���=L�=R�=����>>X�>�o��4�A�,���.>�ً>�弈-.��xu��`�< �U>(�н�R.�5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=r6�񉤻{���&V�}��=[��>c�>,������O��I��U��=��
���ƿU'��v3�� �=r�Y=��;g����TܽR����.��	���W�=)J2>n.�>4�>y�6>|s>k�h?u2�?i2�>�廼(ν�'E��)	�]��o����!ｳR��2F���ʾiU��վm�����,���;i?��>W�U�3ᖿ���k�H�"zR��
?�^ >�Ι��=�Lh����о�o�Z�=W%���)���(�b�p�G6�?��2?�T��c*F�[�"ռ͊��w??�21��߾�����q�=�9=�L8>F�>s�C�{�`e,�#?W���6?���>땗�ƨ���sf>�>"����=78?��?�z>��>�n/?�(���$���M>[\G=�r�>�S?��>a0����ݽ��>�%?�i��ϼﾼa�>�j���I�>>�U`>ӶҾ��ü}e:>��=�@оV��=ϥ<P��z^?t (>�l�5�Ӈ�PL�D�I>$�b?��/?/��>���?֐O?%.ӽ���2�=���!1
>u�R?A�q?:��=X�ѻqa�ȾD�E?$gu?�62=�gv�����z�+�[<��W??�N?���>�A�ݯS�����kI7?��v?�u^��g�����#gW�j��>�7�>���>��9�H�>�>?��"�mN�������h4��?��@���?��C<m ���=�N?^��>{�N�Q�žR������Em=���>�֧��rv����p
,�2l8?���?"��>Ր��(�����=�j��u��?�ք?!:��~�<_�/=^��	���0���=�d��EE�����lF�¾��*�XՖ��G<G}g>]�@۲�<	��>�|̽��޿jsп4ׁ�=Ǿ`=�VK?��>��彝��=�f��6t��#I�(�+�����(7�>AS�=���d���L���52���ʼ���>�B<�C�>:�$���Л|���=��>��>�'�>��s̾ ��?zr�*˿â���"
�M�H?&��?¿�?Qe?�� �H`�-�h�,{-=cs4?��X?��O?r���ees��љ��dk?2���`�����V�����E?�[$?��;��9��/>�-?'>ڟG�	��`x�����쥛?(��?fXھ��>=��?�W?��������kɵ�u�M���.?Ǯ�>�龭�{�L�?8�k�?n�"?�Z�=����_?��a���p���-�
�ƽ�ۡ>
�0�;h\��H��ԡ�.Xe����?y����?#^�?�?F��� #��5%?{�>����9Ǿ�<D�>�(�>+N>IF_���u>z���:��h	>���?�~�?�i?䕏������S>c�}?ߩ�>s�?g��=Z��>�7�= ���"��	">���=�LA�<�?�M?��>y��=�$8���.�O�E�)oR����C��z�>$<a?c�L?��a>'J���0�!5!��w̽�96�џ �+�@�&�(��ڽ��2>��>>o�>cG���Ҿh�?����ؿ5O��U(���3?���>>?�����t�6��
C_?N�>�G�W&��x'��k����?�;�?�?�y׾z}ȼ=�>�ѭ>3�>�Zս�m��������7>��B?��_X����o�<��>���?֪@�Ǯ?��h�	?4,��I���C~������7�v��=V�7?��?�z>���>�c�=�~v�>�����s����>�0�?�t�?w��>�l?,Yo���B��0=�t�>�k?!T?��{�U�LB>�?��[���N3��f?��
@�n@�^?n墿��ٿ���-�������Ͽ=��=�MB>�Tܽ2/�=��=Ԯ7=9��@!�=Fq�>w?�>5׬>��>��s>n">�����B"�����z���fB�s=����HC�����f���ov���Uľ��ʽ�������@f�/��
ꁽ��(���l?FS?�݃?�	?5��=w��>n��Hbw���V��ɱ�3� >�x?�&Y?e8,?��]>Q)�#�\�]�o��î��"����>f�>�b�>")�>�N�>rޅ=�Y�=șv>�tF>���=M��<?u�=l�=���>��>|�>iOi>�a?>4y>mO���>���i�q�t�c+˽��?X���~I��ҕ��i�����Ls�=��,?2�>�6��huп�񭿋�G?�1������+�7�>Y�/?WX?�e%>�°�QMi��*>����d����=@����l�J�(��N>��?�f>��t>ՙ3�t]8���P��m��pE|>2)6?�޶��T9�n�u�$�H��NݾUJM>^��>[�B��m�k����	�9li��f{="w:?H�?�"���氾�u��?��BBR>�D\>yd=pT�=�=M>�}c�tǽ[H�)�-=��=��^>ʛ?-D*�b%�<��H>7���龹\�>~q�>��>��Y?��?K�>�*��/3���=A�*=��>��?ض�>_�E�=M�=$j�>D��=�:!>���=q���l�5>�'��"G��D)��o�;x��T�=�1>vһ=�M��w�<�~?�v��
����뾼���5ND?P ?��=�W<�1"��ߦ�~ݹ�3�?��@#�?�o	��:V�3?H�?~��s-�=��>\��> ξw�L�-?{���X�����	��h#�";�?�	�?�8��=�k��>�
%?�iҾrn�>����[������u�ب#=���>�;H?%K��]�O�>��{
?�?]`�)�����ȿ�yv���>@�?��?��m�]:��B@����>k��?daY?�i>�d۾�cZ�4��>��@??�Q?�
�><5��'���?�?���?��
>�=�?�Њ?�}�>{��<��񽿣�z�����}hT�E?4>��%=�G���2�����YK}�����ϾVN�=�|=+_�>��Ƚ��ݾN��=`��Kq���)��Z�>��>� ?>L��>�j?�
�>7��>i!��3�2=�	�b	�k]I?�X�?�&��f�s�i<,��<z��O�>�Z9?R�ֻL�̾��>�][?�?xea?���>���Xy����������b �<�-V>x��>0�>y�A��M>`Ⱦ/�H��U�>��>?��ྣ�z�|]�I�>�� ?�>���=��!?�&?�ZN>9��>��T�怍�Ӿ!�+V�>]'�>=��>
��?wY2?������%�������J�u�>9�k?��?���=X9�����ã�
�z�MM<Xч?�^k?|�< �P?G�?v�4?��;?n�>by������="��>g�!?�����A��+&�����-?�m?R��>2���KJԽE�ż���]����?�1\?%&?n����`�a�¾��<X�&���b����; ~>�E�>��>G5��P�=��>�=G�m�v6��bb<�W�=���>�y�=G7�BI��A,?�c^�۷��Ǘ=o�r�L�D��>��M>���K^?�<�s�{��!���]���V�?�c�?Vo�?�ʱ��h�=?$�?ca?{o�>�ڭ�}�޾3ླ{�[�y���dw>��>�=j����X`���9���1���{ǽhgS���?��>-�? �5?CI�>�W�>�p�"�E�%v3����ЁG�*~�'�?�դ.�w�͔*���l�ٌ:2Dž$&��#>��=oB�=5X?�\�>d5>�2�>������<��9>���>���>� >e�k>> \>�	�=���JR?jB����'��J�5����VA?|d?�T�>W]c��A�����/�?�K�?�>�?<�v>�lh�+�k�?8��>�����	?M8=Ĭ�u`�<է�������m��[�>>mнY�9���L�EAf��
?�?����˾ �Խ�*��}Ua=S�?�)?�%�p�M�;�q�`T��eT���`�F�o�*ࡾRC$��"n��=���p���Ӆ�XJ%���F=��%?�Љ?,�h�龸W���wl�`�C�Z>���>,��>s?�>��L>I2�}g-���[��(�Jچ���>�p?��@>�a^?��G?fn[?}8X?���>��>lH���5�>��F<���>	�>�1?��:?��7?��.?Z>?��->������� p���7?�F?Ni?��>���>��m�������s=m�i=z��Iu��d]�;:$ =�j��I��<�\I=Rk>1�?~
���/�Ѱ��Fqp>zG7?��>?��>�R���i��=���>p� ?`np>n��P1i�N	�!�>�?G�#��o=I&(><��=V��$l���Б=�3;}�A=>���v�����;[h�=�[=�*�:i^L��ߴ��O�<_z�<s �>��?�ދ>(�>��辀��Y�R=�VJ>�%->�>���OF������\�^{>�F�?�ĭ?A�+=`�.>M�@=L���J� �Z��'�㾅�8�i?�+?2�K?a��?J�T?�K'?wF&>?��-���(��0�I���"?(D,?���>�\���ʾ�稿�S3���?ڳ?l�`�R���>)�.��M�ͽp>ޣ/��c~�oگ���C�_��ì�l���P��?+۝?�;���6���辁=��z.��D'C?2�>Х�>���>�*��eg�5[��?:>ݧ�>aMR?y�>�JH?�`>?�w,?t)�= p��[���7��W�R>�jJ>!�?��?P�?Mh?uI?\E�>ݾE!���e��������?�S>>>TT>���>J�>0�>&�5�C?���� �;Y���'b>�~?64>�*�>Ц9>c�f=��H?i��>�ۿ�V\����� ��l	���5t?g�?S�.?�=G��%F�֩����>���?���?;".?�f?��C�=���%����x�NQ�>�g�>[�>`�=�~=�>��>�/�>?�������9�]C��"?0x>?�M�=��ſ�q���p�r����ac<�ڒ�� e�֔��[��.�=�Ș�¾��ͩ���[������w��q���ϫ����{�/��>�I�=?��=�'�=�B�<>#ʼM��<cJ=ٍ<2&=��o���l<�,9��ϻ�҈��f���Z<A�I=�F�a~˾�}?�<I?h
,?��C?�{>��>V69�Bޕ>�a����?T>°V�n��c�:��󧾀�k�پ9�־�d������>�]>��>6�4>�j�=/��<�1�=�g=-��=�3���J=c�="�=�g�=��=��>/e>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>v�7>��>ӮR��u1�n�\�x�b��3Z��!?�2;�W\̾�n�>|p�=CT߾��ƾ�>,=ѝ5>�Ab=�C��\��j�=�]{��8<=��j=�>q<D>W]�=�K��G��=�MH=3�=�FO>a���7�6_+��L5=�*�=��b>�s%>7&�>�}?�/??Ku?(á>`�4�j����ξu>���=���>�=� >e��>��0?��E?D?�$�>�=,�>��>��/���x���コ�~��;Hڇ?9��?���>�:d=���	=��K-�+����>�A,?��?`��>��� ����|1���?�F�+<Tկ=2�d�/�)�*o�
�$�K��>�^�>��>eĬ>�V�>	�2>n^5>���>��">��;;};�;��!=n14�9�y=M��.�=U�<�#���b�������4ӻ��=���<v6�<a>�	�>�\>0,j>��n>Y����0�=�a���h�F�پ��`�.�=�|���~���'�s���"T>��u>
Q>������?`�d>qK>PS�?o8�?���V��г������޾�:���B>8��=���� ��b2���X��Ͼ]��>Ӓ�>~��>�k>�,���?���s=��ݾ�4��K�>:�����p���q�����l��~�g�T��;>�D?yۇ���=�@~?�QG?hߏ?؟�>����K�ؾ��$>5҃��5�<1���v�#ˎ�7�?]�&?fa�>�u뾼�D�8̾��Bٷ>X I���O� ����0�2���ŷ����>Y~�оG)3�Ee�������B��?r�L��>�O?��?�@b�@S���\O�����E���g?Lwg?��>xB?t>?��u�a��sY�=��n?��?;�?y>P�=N������>;J?�?E	�?��s?�&I���>~5�=�>�o��m9�=$�>���=j�>��?��?�?������n���y�1�n����<�d�=�Q�>��>%i>���=�1v=�p�=,Z>(<�>�L�>Fo>�u�>�>@������S?T��=��>_�O?��3>��;>�Z��.��ی\��P�.���B.*��e^�V>����:�=�ν4<�>�u˿�J�?��>9�>���?�8��}b�c#�>Oa�>0l�t�>]ub>�d�>d?�>���>�h�<�J>β{>�y���=�f(��t-�r�R���B������=U>fy�=��5���5�U�z��0������Da��o�B-N�_H�����?�<��	i�8!�\E����>�"�>��K?���:��5�=��?���>�;��֙�K��I�����?� �?�b>pj�>a�W?}<?��1���1�`�Y�u�u��A�9�d�}�`��Ս����D�
�hO����_?-�x?�A?0$�<F5{>2N�?`�%�YS�����>��.�1�:�D?=�*�>GI���_��Ҿ�FþӬ�DOE>Q�n?��?z�?5U��&$�uP�>�WR?��@?�W�?!�9?�U?Շ��>X�K>�?�>��>|1?'d??�?	�>U˥>��6���Z<�F�dA����T�_~��2�<�O=r_�=J&U�t&X;�Pg=U�=�Eɽ<(<=d4<��k^<�pv=�Ԃ=���=ks�>��]?��>���>�7?,��	8����[�.?I':=쉂����Ǣ�u��aP>G�j?��?� Z?$�d>�B��B�h>�l�>�.&>�\>�i�>�1�p�E��Ԇ=��>��>p��=��M�qɁ���	�-�����<+>}��>6��>T��R_u>��~�ՠ����=8'���w����R�;��d��j���>ATX?l�?*E��L��K��	i���"?��O?6*`?�u�?��>O�b��W��b��
��s>,�����w���_���|.�N>c�4>Rs�-.���d�>�$�Z��!r���6�o羸��y	��B'>�T��ྡྷ#��zy>�t>�Ŧ�G0��^��L&��{$d?�����Q¾p��y�оJ�">2f�>(�>/�=ʢ���6�����+��=���>!�>'펼k<���r=�[D	��x�>ھ>?gS?��E?����i���P�S���v�o�a�(��>G��>�P�>(�Q>0r�=����,3��n��K���>�l�>�d'�;0�Nܡ�����޾�d->+3?!Ϊ<A��>�S?s�>mO?�CO?:�>���>S���7Eվ9;&?��?TE�=FTս"�T�59�5!F����>Ճ)?P�B���>��?��?��&?N�Q?�?�>y� �S@��|�>��>6�W��A���}_>hJ?ؔ�>%Y?{у?{}=>[b5�p����	�����=N�>��2?�2#?��?w�>�K�>.���ك=��>[Ac?~�?	p?���=�?�p2>>��>��=��>�e�>�"?�kO?��s?z�J?�U�>܂�<Jc��~ ��J�s��H����;��D<��y=	�\+r�߱�4��<�Q�;Ƈ��IL��	���E�����Z��;�s�>1�S>�~��7(P>I�Ͼ=���Dm>�=��s�$[m�P6a��'>��>p�?"��>��,��?=n��>���>�`��?k��>�?nA��`$`�Tm;��=�`��>O*>?�.>��[�4o��;!\�s�=�Il?�a?(�H�߶󾈱b?��]?A��?=��þ�b����vO?��
?BG����>o�~?)�q?a��>�f�N�m�G#���Eb��ok��=�Q�>�x�%�d�4��>�7?L��>�a>I�=r�۾�w�,���d�?�݌?��?YՊ?�B*>F�n��࿩(���1^?^l�>>���uP#?����}̾?ߋ����i⾜%��䊫��ȕ��%��~9 �����m�ܽ1��=\1?�r?oq?~"_?)� ��b��^�^�~�+�U�\5�i����D��oE��~B�/Wn�:/��7���Y��z2W=?%O��W9�8�?$�0?ɾH���?�E��0ɯ�����W>9$��j���L^="�����i8�=�7��&c�tZ���?��>�8�>S�,?�P��p(�`?���-�]�Ӿ��p>���>���>���>�`=u�L���\,ؾ�7��쁅��|>�I]?dmK?_�f?߂�8��R�� �$���D��;�b>M�>R��=�3D���ɽo�(���@��bn�������e��̗���:?$6�>h1�>�f�?���>0��𡵾��`��D#�Z[��U�>��Q?�A�>v��>���|�1P�>��l?�^�>�>	a��!� ��{���Ž��>Ђ�>��>7�o>�.�$�[�hE������A9�!��=�1h?1���d�`���>K�Q?oߣ9��E<�O�>>z�!���X�'��>w�?��=[�9>+�ľ����({�o���E)?r8?=���?�*�`2}>4�!?���>���>T.�?��>u/þ=�:��?��^?[]J?AA?ٌ�>Th=]7���Ƚ��&��3.=���>ݝZ>��n=���=S6�C{\�2�N�F=�>�="�ϼ3���	<Im���@<v��<�!4>{�ٿ�\'�y־�=�p橾_�ξ����jS�7�x��8�=�_���s�=���!� �G<Q�6^q���k�'_����?�� @<贾6��&|���t|�Ķ	�L�G>�얾I}$���|��j�ֲ|���墾����f��pl��j`�/�'?5鑾S�ǿ;����Cܾ. ?K, ?9�y?����"�ڐ8�7� >��<�Z��X�������ο_Κ���^?n��>(��r����>̗�>�6X>�q>�܇�����#��<��?��-?qK�>s�َɿ"���ܧ�<���?�@�rN?3}I��1(����'y>�6�>���=&�ɽ&����ѽ�:�>�}{?��?���=-�A����=H<k? ͵�}�&�>�;ɍ�����>�Q�=�����O��9��=�f>�����־@-�=�?�_�}w �LnȾE��=�A<'�� �>2Մ?.{\��f���/��T��aU>��T?k*�>�=�=ײ,?+7H�T}ϿT�\�<+a?�0�?ɦ�?c�(?�ۿ��ך>��ܾ�M?lD6?���>d&���t����=&�R������&V�1��=X��>�>��,����ȆO��X�����=R�ƿ���@�&���;>�д=��-��2�˸ɽjQ�=�~���+i�V9��h�w=V�=>ٟ>��>gS�>�E>�!e?��s? ɂ>ݣ%��r�iM@�F��y�d��o���҄��sh���y��h� ������1*���6�,���7���A�],O>	�S�N��~��GX�׆D�L�?�ݎ=!���D�3�]� ��X�� ����� =�^R���Ⱦ�F5���j����?�F?o��MPE�����D�^����1?�t8�%����'��$�U>	�F=s�>և�> �>{�ľM.��V��N.?:�?\5Ҿ |O�">�&��v��=��0?�\�>�<%ҫ>j[?ʰ�
��gO>���=�d�>9Z?C$T>�ξ��6�V�?�9T?=�нa�~��`�>
�پ�������<�o>z�v�^����K�>\��=7Yw���=\���Wϼ@�T?v�5=d�-��"	�YMվ�Q���O>��=?�g ?�m?�r?
�I?�H3�sg���:�DZ���|=B9L?Уl?��>��i<�o��Q��B?���?|�.>g��q��A��KJ|�pi>�"h?�8)>0*��H7���*��?WG���??��t?.Jb��7���^���C���8_>�!�>U��>XI7�F�>��9?^���!B������5�>�&L�?l�@���?N��<:B����=��?��>�Qݽ_^��;��]c��%Pk���>�����{�O$�90�R8?��?�}?�k� ��x�>b-��?���?�5�����=��<iO�����]=y�=oT׽S���n⾼D�~�����	��(�����<�Nr>�<@���[��>���׿_4ؿ��/���j�e��{?���>�*�5B����a���s�J�U�JA�fS�� ;�>�_>D'׾&X��'������*����= ּ��?�;�@Ѿ@9G�Br�>��?5��>T^u>N̽6��(�?� F�Ѹ��@K� K���:?�+�?�vu?O�Q?� >��o�pƍ�ٕ�=,�H?U*?�C/?Ԛ)>]�_�� �O�i?������S������X����	?�{?�ؾv����>��?�<>T�ޟ��ڝ��ϒؾo��?	8�?0������>GR�?�n?[��x��:gY����6Ɲ�h��>��|>��dYM�v9(�0;��-��>q�/?� >$9&�\�_?%�a�[�p���-��ƽ�ۡ>��0�0f\��L������Xe����@y����?H^�?a�?���� #�D6%?6�>�����8Ǿ��<���>�(�>*N>LG_���u>����:�i	>���?�~�?1j?񕏿�����U>�}?���>E~�?Lx�=+
?h4>�����aI=_>V��=C ���?m�=?���>�Z�=@	 �w�;�]75���6��cݾ�MP�a�>��j?(]K?	��>�DV�r�r��m/��5��k�jnQ�d�a��PŽ����%>�B>�v$>� ����þ~�?n���ؿra���'�p)4?���>m?���e�t�V��=_?/|�>�<��(���$���N�a��?FD�?��?7�׾��˼E>g�>D�>��Խlݟ�������7>&�B?�C�6@��Y�o���>���?Գ@�Ԯ?'i�=
?�P�{h���#z���	��CX�2Z�=�e9?�F��]>|��>5~�=��z��a����v����>��?Q��?x��>�d?��g�uL<��=���>;�h?�A
?˼n�����45>q�?V9�5#��1� ���c?�/	@f1@��\?���hֿ����^N��Q�����=���=ֆ2>�ٽ-_�=��7=��8�?=�����=u�>��d>,q>E(O>�a;>�)>���P�!�r��\���R�C�������Z�C��Xv�Wz��3�������?���3ýy���Q�2&�?`�f��=��Q?ON?�U?_t�>��<���+>?���=�߃�}:�<���>*/6?�B?[8?y&�=Zx���P�
鄿���6�l�_}�>v+>�x�>���>M_>cr�=�f1>���>�>��w=>~=!�;=��=P�>yD�>�h ?��>�C<>_�>Kϴ��1��v�h��
w��̽�?�����J��1���9��/����j�=<b.?I|>���?пe����2H?|���Y)�v�+���>V�0?�cW?�>���@�T��9>]��l�j�P_>D, ��~l���)��$Q>�l?GCg>]Nu>I%3��I8��P�Q����>z>�5?յ�Ԋ9�jWu�b�G���ܾ�N>�f�>��>���G얿�-��oi��x=�*:?7s?�߳�.����v�Y���kR>h�[>p�=�!�=�M>v<b��Ž�IG��g.=�G�=�g^>�(?璜=�y�=쳽>F�Ǿ������>s��>�M�>5�=?5�\?�A>꽐�罚3Խkg>�9�>%��>�!F>&�Q���<�ȿ>�*>�z������M)��w]��0Q> ��5��j��o�r,���=X��=�۫��wW�k�<�~?���*䈿��De���lD?Q+?? �=��F<��"�B ���H��G�?r�@m�?��	�֢V�8�?�@�?�
����=}�>
׫>�ξ�L��?��Ž$Ǣ�̔	�6)#�iS�?��?�/�\ʋ�6l��6>�^%?�Ӿm�>�~��Y��C��P�u���#=��><2H?�O���pO�>��v
??rb������ȿ{v����>'�?��?�m��?���@���>ǡ�?GdY?�mi>�m۾�pZ�ov�>P�@?@
R?�>~;�[�'��?�ض?e��?uY>t��?b*q?�6�>��q���߾�����Oq�/�<VR=�'|>�M>���w�$��H���w��w�^>���>��/=P��>���� ���0=��D�����g�=�>��> �>���>��>W�>�ͣ>��c;5�D=�/����J?KЍ?!����k�A�<�_6=Tm��Y�>�5?�*����˾��>MZ?��?�l\?x�>���9T���Y��r1���A?<a?M>���>���>@�r�z�;>� ;GOA�W:�>Q$�>����"�׾��~�.Q����>��?���>�ͳ=�!?�~?�u`>���>ˁ2���q��$��8�>�p�>�S�>�tv?dN?��g��� /���o��BS��>�6f?��?��3<���������J�j��x��>�z?|�g?gF�=U4?�S�?[�Z?�dA?�j�>SѦ=n���B>���>a�!?���ϧA�L&�K'�;[?_6?���>���ս�ּ����h��' ?%(\?�5&?[���1a�þ�!�<��$��M]�|��;LIF� �>��>sX��^�=��>s߰=�m�#$6�^�g<{ؼ=�|�>�'�=�!7������4,?,�'�7|��=,�o���I��q>�nn>|Aоm�K?�K?�Q�q����aN��!�q�R��?�e�?혔?gҦ�=Ck���A?x5�?�?��
?������ؾ�WѾ#����vx� ~�]5�=]�>b~����;�������߽
U.���?n��>H�%?�F?���>�3�>Y=���9I�ՇI�6!��I�QL���:�A�����Q2�/�ܽ�d�:L�����!��>�e�=,z2>�ڵ>�D}>���==&�>��5<u��=�����۵>:�>uQ�=F��>��U>����\�ʾ:R?
ǿ�`�'�p侓\��	D@?�d?���>��S��P��H���+ ?@l�?��? �s>uh��+���?Dw ?�����M	?�_:=o?k���c<�ʶ�1��b��o��>X���6e9��mL�2�\��?+?p�'��yǾ:"޽����P�t=��?�'?Q�%��B���t�1�K�4O�!|����b��ͦ��'�L�i�����0���b˃�$�,�By=]�#?@І?�d��C��Jh��WL�&8>#��>D��> }�>�R{>T��K�+�~�W�}�&�����2�>7xm?Ψ@>��`?�h^?��`?f�a?^�>?!^��@ɴ>S �p>�Q>�3K?0"?F�<?l(?s7L?pq>p>��% �eA¾��?��?��'?'9�>o/�>�AH��=<=�9F>+��<�Y>�]	�l�7=�X�={�����:�=�a�>��&?ʲ:�VF���ƾ�� > /?�
?�N�>�h��$�آ��� ?��?1w<�n �5����%�)��>���?.H	��=6��=\z�>�<\y��&z==��>��=�G`�a;=5$=�?,>f��=�e�=�柼ur=��o>�%��n�>�?|��>�V�>�4��g� ����$l�=��X>p�R>�>�6پ��������g��y>an�?�q�?��f=��=���='���lb��+��1����9�<��?RJ#?GKT?7��?w�=?rv#?м>�3�FG��{Z������E�?�-,?'�>9����ʾ�ᨿ�3�`Y?�m?F�`�����-)�����WԽ��>JM/���}����D�L����[s�����?��?�*B���6��u�h���O���}C?�8�>k��>�(�>�)�H�g�&��:>]�>R?��>ӝB?)h?��<?W��=��R�́���$��_o�=E��=�e-?���?��?tp?4��>g�>�ł��c��������_����a�ꖒ=P�>�>���>�t�>V�=�٪��G�7��3��=+BT>���>�,�>�͟>A$�>��=xH?O�>����} �ť��:]���,��u?�L�?w�+?���=/��ŇD�����`�>��?�u�?�)?��?�j �=�a�(��;v�爳>g�>�]�>���=�&(=�z>���>jJ�>m,�G���*9�DLZ��>?�DC?yA�=��ſw�q� Ao�1%���]<#��T�d�Vᒽ�\�{ͤ=�����i�����[����풾"���񲜾�8{�a��>�G�=d��=�^�=V��<�0żUI�<~�I=���<�L=2m���d<\;��罻VJ��Xp�rZ<LvD=�nл�ʾ�v}?^'I?),?=�C?/|>��>�}6�>�>\����i?u�V>?�h��H��p�9�7���&���Dؾ)׾&�c����4�>ŅE��o>��3>|��=�v�<7��=)�l=h1�=_iR��=���=��=S��=Gd�=��>�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>z�7>��>�0R�~`1�-�[��"e���[�~v!?��:�X�̾il�>�=!n޾��ž"2=/�5>BW=@��8E\�Z��=8�}��@=1�p=�4�>E,D>��=�꯽�+�=:+L=���=��N>\����05��}-��79=� �=5�b>e%>���>��?��/?fId?a�>��t���˾������>�5�=�$�>���=�UA>$��>��7?
wB?hI?�G�>�ѐ=5��>���>�H,�ol���Y������<=J�?`|�?��>�=�<A�8�}R�=i;��[��V?	R1?��?�7�>���A�Ῡf�-�$����=�K�<�	>vȼ���X=���k�]0'��9%>u��>=�?Վ<?��?��{>�M"<i5�>���=�Ս=Iւ:�F=A=D����=,k�u��=�n�<�=X��<�k���W��S��5�<o?�=DvS=��>��>�n�=y��>w�^>�ٚ� s3>(Xһ7�n�fU��鯾K��
u�]��� �6'��a�n>�:�>��D=S��1? ?r�:>��k=_U�?9o?¶> �E�A�#����対�4}�m�,>�f5>�I�Y;Y���a���+�<u�����>b��>Dg�>��o>[>*��8=�=�Z޾~�4��+�>G��?��O���p��Y������"�g��M;[/E?�;����=l�}?T�I?WM�?=��>3�����ؾ��->pZ��e{=�v�q�ժ��ʲ?l&'?S��>�꾕jD��=̾���ڷ>�3I���O�{���^�0���3÷����>��o�оe"3�Ff������0�B��Nr����>صO?�?>Bb�\U��ETO�����]��1y?�zg?f�>>I?�A?��wm�l��cn�=��n?���?�<�?K >,	�=6i�]%�>��?���?���?�{v?��:�n6�>E��;�S>|�ѽ�>�O>��='�>��?ԧ	?�?�>����D��w8��J��<<ϔ=@%�>��>��>ۼ�=���=���=��U>�d�>o8�>� _>�)�>�[�>X��u��[U+?Zb>JR�>u�+?nQ>Zk>� e��ѣ���`��p�����b)5�H;��~�=g�n����=�경W(�>#t��T�?��>��3��&?r}����:�}�4>���>TB^�4�s>[�(>�{>�L�>�
�>�Gm>E��=2 P>E�Ҿ�M>���� ���B���Q��SҾ8�y>(��x&�A����K�t`��+P�Ej�|��H	=���<�?������k��)�����/?�{�>r6?LL���Y��,�>{��>���>����w�������B�� �?j��?�:c>��>��W?��?:�1�� 3�AsZ��u��)A��e�Ǻ`��፿����͖
�'����_?��x?~rA?��<�5z>��?0�%��ӏ��%�>;/��(;��)<=S+�>z$����`�v�Ӿ��þJ0��>F>*�o?�!�??T?lNV�eĴ�4z>hcM?(�:?�.�?r;,?j�J?���?�?�C>��>�A�>�|C?�B%?�p?Ljj>�rC>7L�<��=kܱ�Z��O�޽��ٽ�'�:�;:=�oD=���:(�?=&�Q=^L�<���<�p\�'X����z�x;ɶu<1՚=x� >���>��_?8��>�َ>�;?����2�;����+?�J=l���q������z4��>��j?>�?�X?�R\>.�D�:�A�v�>�ʈ>>�/>^EY>=�>���t5�!��=Wq>�l>4��= [�8Á���nX�����<�8(>y�>�/w>m��<��>�Ũ�+�|�t�=�P�g��iGJ�@�#�~v���t�>&H?�?ۣ���q�a2��`�y�?3?m�h?�j�?t �>]M���U!�*;G�	<���>������.��Ǜ�����&S��%�=B%M>�5��k���>�N?�^Mž'����*�8�{���>}ࣾ �
�i����,澘v���e
�a>�=���!��:`��f調�G?�==�|����(���,R>=c�>��>���=�%!�'��w^žp#o=�#�>� �>sd�=�
�h_U�ݘ�V}�>��N??{?��s?�O��5����X����Xg�\�=c �>���>�?���>�q�=�Ğ��9&�S����]m��ֽ>{.�>%J��x��%�m���HM�<%�>|�?߄Ƽk��>+F#?�J?1�e?�s?F'�>��>��%���оC[ ?Y��?��>  ��}�z���H��)�Ǌ
?��/?�BǼY,[>��?X�?��?�N?d�?�IR>~>ξ�#�e*�>-x>byR�����x)�>��T?�
?5�t?�z?�y�z�E�+���j̛�n�>[�%=%"?�I-?�(?5�>Y��>2/�-��=�/�>V%�?F�t?ȞK?W͑>��4?a^�=�=D�½�>M��>y�"?�Rd?�Є?��6?'�?n�+�D���F�� �<�c�=O՞=����1�|�N�=^亽�m�=��P=�){:Dl;�9=��<��.�A<���V���m�>�Us>�Ɩ�r1>o�ž����XSA>�U��<s�����'p9�7�=|K�>��?9g�>�'$�H��=�M�>׵�>�H�N(?�?
�?��p:c�b�:Kھ�L�Ѱ>��A?�X�=i�l�D����u�qf=��m?bQ^?=�X�r��*�b?��]?'n�=���þ�b�#����O?$�
?h�G�H�>n�~?W�q?[��>@�e��8n�!��fCb���j�Aڶ=�p�>�V���d��<�>��7?�O�>�b>0�=w۾��w��s��?��?��?���?�!*>��n�4࿰]���E����]?�r�>r��#?���2�Ͼ�0���4��V��^�����[G���|��"�$�Aۃ���ֽ���=h�?�s?hCq?��_?ƹ ���c�^�N��P]V��+�S���E��E�b�C�}�n�H�m���C����F=h&Y�̺>�֎�?M�?�c����>�����}�ɤǾ���>��^�T`��m][��Mҽ!~=Iʽ�:��6������S?��>���>&�n?C�Z��<�3�5��Q`��i�L��=�:j>:��>۷?�2= �ż�m�<��վ`4��MRe��v>lc?��K?7�n?�� �G51�@���é!�*:3�\ ��#
C>��>H�>�(U�R��%��N>��s�&�(����	�.|y=��2?�Ԁ>��>g�?�?�	��᯾c6w�\^1��Ҋ<z��>)/i?�.�>�^�>�<Ͻo� ����>��l?���>Q�>����T!��{� �ʽ��>J�>���>B�o>��,�� \��j�����99��q�=��h?z�����`��>�R?	�:�H<�u�>�hv�I�!�O��4�'�~�>�?�Ū=�;>�ž�"���{��5���j?��?d""�u�%��>3�?�?�� ?��?�o>F��[�� ��> .B?��9?(�G??'|->qJ{=��z���P� j�>dU�>��#>���;Hk��N�9JK�q=w�<�\������3<�a)�G;�7L��dd>�LϿO�H����\J��`ؾ������������J��<t������Xþ섾F�,�ѕ��p�2��D�Kq�����o�?,`�?O�JL��U���U�u�2!
?����ը6=�"C��Y0þ��㾸:��V]�5�r�6h'���c���=?j����ƿ�ٓ�ZX侸D??��G?̀?Q���fI.����b�`>9'ɼ��>I������-�ݿ�4���[S?��>�P������a>��>�̶>�U�=\���W�=�>�JZ?���>ɯ|���3���D~�<��?"@�lA?̹(�dC�M�S=�<�>��	?�:A>u�/����u�����>Tߞ?���?�wH=�W�8/���d?��<a�F�������=���=�=�P�1�I>���>є�#{@�� ߽"Y6>�.�>{�!����^�o;�<��]>4�۽阽5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=s6��{���&V�}��=[��>c�>,������O��I��U��=Z ��>ſ`��O+���=2!����W�0����V�/�Wپ+���i��Z`�=��(>��>�_�>�c>I�k>�L[?�j?�A�>�>'�&���v�ǚ��eF=��=�
/��� ���=��5����뾀�����,�_	����L6�XTc=±W�҇���'�PW��H=���2?��4>p�ξc�C�d��:�;�E��%ױ��Z�@h̾��'�ik�Ç�?j�<?8	����N����T���X��3O?<��yR��,����=�ҝ��'�<���>%$�=�۾�71��bO�[0?r?���^#��8�*>�L ��"=��+?��?�(Y<���>��$?~�*���㽷�[>-]4>�L�>���>!
>��U�ܽ�D?uT?z� ������V�>����,�z�j�`=9N>A,5��/�H[>���<����>tY�Wq����< W?^��>�*�r�����d���#>=��x?G�?+�>�}k?}�B?���<%_���S��(��w=�W?i?��>�����о���C�5?M�e?��N>u�h�2��S�.��?��?{�n?�R?��0[}�������T]6?��v?�r^�qs�������V��=�>2\�>���>��9��k�>��>?�
#��G������Y4�Þ?v�@���?�;<� �"��=�;?B\�>j�O�??ƾ"{��܃����q=�"�>I���Uev����IS,�\�8?ܠ�?u��>;������X�>�%g�̂�?[w�?�=��!��<25��5{�a1�T�^>@�=*h�=��Ѽ�Ҿ�����Ͼ���~��{�/���f>u@��z����>�R�HK޿Zÿς��+��G��5\�>�`�>�ft>���myU���,��G^�oa]�`��뎣>��	>�ǽ̉��}�~�k5�a�׻���>kь���>�?I�j�����v�;	��>b��>��>�|��� ��Vz�?���s1Ϳˡ��݃	��W?�c�?`��?�?]mo���f�s"r�����+�B?z�j?6 W?�b�Cf�ӖF�]t?�>��B!V���T���A����>X�c?�Y�>�?a��?�=���=��D?/��bV��D׿8��)=��q�?Q��?�����>t�?c��>�������y���;B�@]����d?f_��$B�����F����t��E�?s-?��8�)��^�_?'�a�S�p���-���ƽ�ۡ>��0��e\��L��<���Xe����@y����?I^�?d�?���� #�S6%?�>f����8Ǿ��<ʀ�>�(�>*N>H_���u>����:�i	>���?�~�?Lj?��������U>�}?X#�>x�?K��=�g�>�i�=��
�-��_#>��=0�>�[�?�M?�O�>m�="�8�./�wYF�aIR�L%���C���>��a?�L?WKb>=���52�"!�eͽ�^1�4o��W@�ܡ,�ŝ߽j&5>q�=>�>i�D�Ӿ��#?�@���׿t敿��%��A?���> ?�� �	X�����<�a?w�y>ߩ	�n7���Ԑ�R59����?���?Rp ?�aо�N:;9i�=c�>��>$����µ�_`��g�S>�<?���M芿M�r�@XD>Hj�?|�@�ĳ?p_��	?��ZQ��K`~�����6���=,�7?Z-���z>���>��=Gnv�8�����s����>�A�?�z�?���>��l?L�o�T�B���1=�I�>��k?�s?�#q�󾫭B>L�?������_L��f?��
@�t@�^?���Z޿vm���6��W���#�=�3�=�l>���ǽu=��T�������%>A�}>��W>À�>��b>�o?>�S>\L���E!�uA���V��hA�x���D����^���:;"�T-��WT⾺��bD��E'���(���&��(�>�N?zO?�g�?���>��Y}������R=ؽ)�;*=D�>^P?C�V?�1?&4�=>E��i^b�Q�t��0��k؀��ȧ>�	f>ϳ>=��>Ϟ�>DG���l>�uN>ܼ>;�=`�v��������<�>�;�>���>�[�>]�>�^�=5������y��s�C���=,�?5"���O[�kf�����I�ľ�>C@'?�l�=G���|h˿1��
�8?���'�'�m�.Q�>@�+?^Y?��G>A�����<�.�=o�A��w"�F��>���ك�"�L�>��6?�g>�$t>E4�38�?tQ�X믾@�}>�A6?�z��&e;���t���H���ݾS�K>�r�>��F��p��閿�d��*h���y=nb:?�S?놱�s簾	�s��j��tS>0P[>��=��=�M>�;Z��wýJ�F��t#=!�=�E]>�Y?�Z+>���=֢>�M��֕L�·�>='E>��.>�>?]�$?�+�ꨙ�����Ee.�4t>Y�>���>�>�	G�u{�=���>8{a>�R
�5=������sB�zHW>�&��[�\�G�z�r�x=�_��w��=�Й=���"�@�82=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿx9�>/��>��ԃ��|���=O(�>�L?SW��,��J)��?9��>�����.�ȿ�dr�\��>�v�?A��?�g�����&�8���>?|�?��[?hfG>u]վg`��U�>�>?��M?�3�>������k?a��?R2�?sI>̊�?��s?�P�>�	w��{/��+������*�{=�{~;�p�>\�>�m���F����� U���j�k��a�`>�K$={�>gi�;���ö=��������@Zd��з>obp>W�I>k,�>� ?���>���>�=����쀾�Ж�t�K?���?����2n��P�<���=�^��&?hI4?Oi[�f�Ͼ�ը>
�\?t?�[?d�>G��I>��?迿1~��0��<L�K>4�>hH�>$���FK>��Ծ�4D�&p�>�ϗ>m����?ھ-���T��GB�>�e!?���>�Ӯ=S� ?_�#?��j>'�>�`E��8���E�&��>l��>|H?]�~?��?jչ�KZ3�j���桿�[��;N>��x?V?�ȕ>�������3�E��:I���Û�?)tg?�S�0?2�?R�??Q�A?�&f>���ؾ����]�>�1$?�&���K��� ��#_��?R�?�6�>��ܼ�)�4�<���p���U ?udS?��?t����`�Q�پ�o8=�x�ۚV<�H@<_�����>�o3>��>����=�|> �=bhv�j�/���>=�3�=�#�>X|O=�2U�PR½�C,?j�J��ă��=y�r��wD���>�L>A���^?S�=��{����>���E�U���?���?�n�? N��#�h��!=?7%�?�?�>������޾���#Aw��ax��[��%>|��>!�o����"���(����R����ƽ�#���?婚>~��>l�?��e>r]�>���x(�!_����<���x�b�9�a~J�E�6�c*��$��Y �"�>=0Vݾ�A����f><ex�0"�>�d?�6>r��>�1	?;� =z~�>�7�>�l�>7�	?�A�>G80>��>�ĳ<�a~��.R?����j](���GR��ZB?�jd?���>�b�6w���D ?~!�?�
�?��t>q�h�o�*�D?�E�>�h}��1
?��4=��M�v<���-5��>�����母>�ҽ��9�ȚL���g���	?�x?f*����;��ٽ�����n=N�?��(?�)���Q���o�ϸW�S�Ù��6h�:j��H�$���p��쏿�^��%����(�`r*=��*?j�?͌��!���&k��?��df>T�>K$�>%�>uI>��	�g�1�e^�M'�T���RR�>t[{?��>�E?�3?�LZ?�nA?;�>W��>\Հ��] ?�(8�6>c��>�G?r1?_38?>?�-?�0>�r��o����پݹ�>�a?Z�?��>�E?37��L
=/f����V����1��s�<aT'���*�2y3��Y$=	��>�U?x���8�:����k>(�7?��>)��>����&����<1�>ر
?�A�>� ��}r�`��R�>���?3��m/=��)>A��=腼t�Ѻ9I�=s������=����u;�� <i��=y�=@�v��_��`-�:њ�;�@�<�s�>��?���>6B�>�>��m� ����se�= Y>�S>�>Gپ�}��o$��[�g�Zy>Xw�?Yz�?��f=��=Ґ�=�|��iW�����#���n��<�?mJ#?�WT?��?��=?ik#?ú>�*�M��S^�������?.#,?&��>\��۽ʾ�񨿊�3��?�U?Aa�{���;)��w¾�)սJn>c/�j+~�x��AD�M��d���b�����?}��?��@���6�������Y����C?�#�>H@�>]�>��)���g��,��;>zm�>R?u��>�9S?Ni�?�ρ?4��>EP��V+����ܽ��&>m?П�?���?l&�?��>�_>�6ξ��)�V+?�s����h��ö�"g>7�=1��>���>�>P>fI>*���S�<!����u>�L�=��>n�>���>$[�>�,>>�]D?޳�>�E���l�nI��FK��M�
��Y}?��?�+?�Y�:T���;�o��E�>iG�?Eɫ?|+?X�I��*�=�+M��(þ�с� ��>���>K�>���=V�=�3=��>�C�>WS�b��8��3`���?"�D?Ǡ�=B:¿��o�|`���s����r�����V�ѩr��M�Pш=C���ۉ��K����]�_k��:��������Ӎ~�"�?�*�=���=(!�=�'<Ὧ��=ʆ=�F�<{��<�$�H�]<�4)�U8j��8���5<n��<#��<�f�O�˾�}?8-I?+?��C?�y>�B>zA3�ǎ�>�&���L?��U>Z�P�|}�� �;�ʸ��v��
�ؾX׾��c�{�X>5=J���>�83>_�=~U�<��=w�s=���=WH�^J=�S�=��=�)�=`��=$�>`;>�6w?B�������4Q�_罈�:?)9�>�|�=��ƾ�@?_�>>�2�������b��-?J��?�T�?��?�ui��d�>9��⎽`r�=����=2>��=B�2����>��J>y���J��*����4�?��@��??�ዿ��Ͽ�_/>��P>sg�=�la�:,������%�7�!��$!?$(��Xؾ�c�>v~�=�s��$ξK[R<4>Z�D=���Z���=�c�Q7�<�4}=�yZ>yE)>���=`/����=�Ԏ;31>u+>�T�}��7cE��\�=���=�>0�=�}�>W�$?�n<?�"�?)/�>�o��;ܾ"�ƾrt�>3%�>��b>p��='�>�)�>[P?�3>?}E?��>D&>3.�>�;�>�U��P��_���2����>e�?��g?�?3�=�䆾��(���/���=�
?�?CS?�Η>Z�	���)@����8�Zx\����q�0�r�"�l�z�#TϾF���j�!�=>;W>u� ?X�	?*��>�M>���>�B�>�i4>Ă5;¥���<i�!�T0߽R<>O�S�c,��+�������ս���=c��=�<�=�2'>N-�<p�d:	��=f?�>K>�<�>n��=�#ľ(;>G虾��_��P>��C�@�Y�;cy�2���
F��ˌ��C>��@>��=��ژ��S?���=Zsb>��?[{~?l�>�#��~���M|���w�hg����=�N>�6}��G(�(�>��J�ag�����>���>.פ>���=��$��TW����=�\�0Z�O��>��Y��T�Z�������D��r���7�_���p=�28?&���M�>�oM?6�Z?aL�?���>��m�d����,>:���/�>m�l�P����(<�?Jz�>���>� �spC��̾ۮ����>�RI��.P�����=k0��K�J����>����O�оg 3��T���ޏ�S�B���r��>�>fO?�	�?Tb�h��O���߫����?|6g?i�>�#?�U?ط���+�lQ��Kڶ=P~n?��?&�?��
>L��=��,����>T�>-=�?CW�?�`l?^a(�3�>�=�sU>��)��=7]�=�HB==��=��	?1�?�3?�ê����1�� ��Eb�&Q=�RQ=�Ǚ>O�>��y>�=Sc�=5f>�Ǉ>��>�_�>�[> ��>$f�>�@����վ#�?5�L��>��6?�6j>�>J����>�p>-���P��	��J☾�㒾��:���=g�9=���>�_ؿ颬?�M>���02�>b��=RL��F >���>������?,����>T��>zc>��>g/>[�(�q�þ���=���nP�AP��@7�������>r�\�'�E�w�澪���Vs�@g���%��g�t��iz�����pܼ#��?D�Ƚ&%����|���?B��>�t1?�Ac�:%�Q�X>�?ܤ�> ~�Mȏ�~��C�۾��?
��?�;c>��>F�W?"�?��1�)3��uZ��u�^(A�!e�X�`��፿����
�6��-�_?�x?+yA?�S�<":z>K��?��%�Lӏ��)�>�/�#';��?<=t+�>*��
�`�{�Ӿ�þ�7��HF>��o?9%�?rY?9TV��3���<>�9?'-A?��o?�-?e�,?�$���%?g� >qW�>�h?T�7?��.?��?d	4>�>{L��rE=�L�����&`���C��s�;t��[��=����bT<�n�=�fn�����i�f�A���E�>Ʀ<ޖ�=���=��>62�>+]?3Y�>y �>F@?��轤�%��%���9?=�ˮ���������*!ھ�U>�El?���?a�X?�m�>�5M�ɔS��>	�>�M>>]�v>�~�>�B���G��I=ߘ>>��=�[��t�Z8 �����3�;�j,>R��>:|>����r�'>}w���-z���d>��Q�>ú���S�'�G�
�1���v��Y�>��K?��? ��=�V����)Hf�,)?-Z<?vMM?#�?��=�۾��9�`�J�.C���>��<���鿢�|"����:�7��:ջs>Z*��.).��=��8��,;���!�`~���B2>�����=���`�8־���=a�B>53پ��3鋿Y񰿞�??d��<�g�����8���N�=���>l��>����4�G���5��|�E ��Vv?�O>a�<�
�T$]���!� r>�TS?;�r?{�?W�b�������Z��/�S�C��=�?�M�>fd<?�#�>[e�=yk���-������ao����>.�?��	[��Ž�u�X�E��|�>�7�>�2<\+?iQU?�?R�U?IW;?v�"?p��>Hu��ξ?k+?$��?��=�Fڼ� N�6�2�S�G���?��??�D9�w�>��?�o?	�?E@?� ?#�[>�2澿� �.1�>�c�>s�?��餿��>>�E?{��>o�q?�܂?Z�9=��M�ka޾0��/C>��D>��4?��?s?&�>���>pW4����=��?&n?[�?�H?�!>�f6?���=Z ?�K�I�>�#�>k<?�zc?
��?;�?Y�>s��S���z-1���ݼ��!>�S�=-\�=\��=I�=kۿ�ӭ3>6�T�9��=+�=���e����6��F���'��%^�>��s>���z�0>n�ľKK����@>iQ��0N���Ԋ���:���=��>��?���>�[#�ȼ�=Q��>�E�>����4(?��??�Q ;��b�0�ھ��K�-�>m	B?���=`�l�U���p�u��h=L�m?4�^?��W��%��P�b?�]?�g�=���þ4�b���龣�O?��
?��G���>[�~?�q?%��>��e��9n�����Cb�n�j��ж="r�>.X�H�d�?�>v�7??O�>'�b>z%�=�u۾H�w�)r��?��?�?���?+*>C�n�94�MK��BL���*^?�K�>���% #?h�&оv������9 ⾄˩�i���q%������F�%�-̃���ֽл=s�?Ds?_q?�e`?��n_d� >^��/���NV�-���[���E�K�D��NC��an��/�=����l���d?=_oy���L�JͲ?g?7�
��I?2�Z�/��3پ+ob>*��!�I=���=�!��BM�=�v��KT��+�jG��j�?ѡ�>I��>�0i?*�u��4V��0��$P�*��r-X>'�=��>l��>.�;�a��U��T��|\��2R��27v>-yc?��K?D�n?n��+1������!�3�/��d����B>5k>���>:�W�ߙ�D9&�lX>�t�r����w��	�	�N�~=�2?�(�>ƴ�>�O�?3?{	�l���kx�ԇ1�;��<{0�> i?@�>��>�н�� ����>��l?���>��>떌�mZ!���{�ŧʽ8&�>�>��>��o>X�,��#\��j��Q����9��u�=&�h?���>�`�F�>�R?'�:C�G<�|�>{�v��!������'�2�>a|?ǖ�=^�;>�ž�$���{��7����0?��?�ef�����0l>u4 ?��>���>.��?C3�>K���:犽�H�>�3V?}uG?"�W?mX	?3�=TU��:���,�a�շ�<�V�>=�> g�=�58>� ��c틾�Dk���b�y�5<$\� &����=���<��=���=y;>�ؿF�P���y����{��H�����]��MS�n���s$��/�����)�l��?��_�<�l��1���6*S�PrL����?S��?��ྠ=O����	f�Ku޾x��>�퐾�w��S���Ձ<`��E|��5��{�R��%6�H���^��:?�㾾�uſ>����[��?}aD?��}?_~�K�6�.�W�� �=�&�;詼;T���ܒ�M�ڿ�����C?U��>�ؾ_\�=
�c>F��>�S@>sx><����N������>��b?d?k���ʿ�����$����?F�@�|A?�(����&V=���>;�	?�?>[S1��I�E���aT�>h<�?���?�zM=S�W�I�	��e?|�<��F�t�ݻ��=�;�=�G=@��V�J>ZU�>��CSA��>ܽV�4>څ>�~"����]�^���<
�]>�ս�<��5Մ?+{\��f���/��T��U>��T? +�>Y:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?8ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=�6�+���{���&V�z��=Z��>b�>��,������O��I��V��=�T�>�ǿڱ%��U�m��;�a�<F�ow콪��;m�4��8�#�������܏>m>-�q>3�R>w�^>�m>e?��j?��}>�:>�*R�ZĈ�������=�F.��[o�"=t��fĽt�þt[�.��J�=���/����~{���I=�r�>=��V�j��P�#���\�>@��Q1?؅*>�;�Q�;�<�lž���$�p�0�˾�)�0j���?�>?������S�.I������豽�V?p:"��2 ��Ѡ���>�lƼ�E�;���>�N=�Ѿ�9,��2R�z�0?*�?�����`
+>�|���y=��,?�k?:�<v��>[P"?	m-���ٽ�-a>u&@>��>��>7�>[������2�?�T?�3���g���Ӑ>wNľ r}�iT=��>�8����O{T>���<�����oػT����q�<�(W?՛�>r�)����a������V==�x?'�?�.�>#{k?��B?�Ѥ<�g���S�0�pfw=��W?�)i?p�>/���]	о�����5?֣e?�N>�`h�z��g�.��U�$?��n?Z_?}t��vv}�F��:��dn6?��v?s^�xs�����Q�V�g=�>�[�>���>��9��k�>�>?�#��G�� ���yY4�$Þ?��@���?T�;<��T��=�;?k\�>�O��>ƾ�z������5�q=�"�>���ev����R,�f�8?ݠ�?���>������#��=Y���0"�?-6�?A����ǖ�G���,�����/�;>-�=E��=,�7=�<˾��i7־��� \���%�*f�> �@膽� ? �g�H��oֿ0I�����R�/�?��[>���=�E��g�m-���a�\�j�¾�Q�>��>8����葾Z�{�c;�oe��1�>�����>��S����ϛ��S*5<�>��>���>����ݽ�e��?�T��6ο*������Q�X?e�?$m�?&g?<(7<tw���{�d��*G?��s?�Z?39%�Y5]��l8�([v?��I���}��V�v�=��P?i�t>.��/.<�4��e�?��=�Af��oֿ�亿b�(��g�?G�?!K���>�r�?���>��	��n��4��yUU�x۽Ϭf?�_�>��ľV��Q}x�实�bx�>.V?Vfd��x�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?7$�>�?.r�=�a�>2e�=�򰾽6-�`l#>�!�=��>�)�?N�M?�K�>�Y�=��8��/��ZF�aGR�$��C���>B�a?��L?9Kb>���5!2��!�Yuͽ�e1�lS�hX@��,�>�߽)5>�=>�>�D��	Ӿ��?�q�I�ؿ�k��}'��34?�ƃ>��?�����t��q��=_?Gt�>B7��,��|'���l�d��?�E�?��?��׾�ʼ��>��>�=�>�ս[;��>�����7>8�B?J
�A����o�'�>x��?��@�׮?v�h��	?���P��Sa~����7�j��=��7?�0� �z>���>��=�nv�ܻ��S�s����>�B�?�{�?��>"�l?��o�N�B�^�1=/M�>̜k?�s?�Ro���}�B>��?!������L��f?	�
@}u@[�^?(�տ<.���}����I>x��=Em>��8�;&���k=7ݽ���@>&��>��R>`a~>9Nj>�[Q>g�/>J܃��%��M��1���N�=����R�Ud����q{����&῾"�оXӋ<c�ټ��@=m4"���潙ԕ���=��U?iR?��o?�� ?T ~�r�>]3��2Z=�#�2�=�"�>�[2?7�L?.�*?�f�=�0����d�>��v1��5����]�>��I>�H�>���>��>mi.���I>N>>,K�>�S >"�$=���5=��N>s�>5��>��>�	�>��<2����[���Q��_�2�720=>��?c箾�UD��F�����[;��bj>T�?��=Q���Y^ֿ�;���5?2���X��l~��(e4>H?;�f?�h>�Ҷ�e�݋�<��ҽ��e��=������'��gF��� >h�/?��g>�xs>�4�"y8��4Q�@��x}>1]6?����y9�4�u�t�H��	޾ yN>Ո�>��R��y�����p���h��{=�8:?��?!���#谾�s����m�Q>��Z>�h=���=x�N>sTb���˽�BG���$=-��='�_>�?V�.>h=�=�>�{���+L����>��H>?�5>�t@?Y�#?m_��8���D���)�w�}>�]�>�z�>�`	>�I��X�=E��>\�_>%��qWw�t����=��W>L���U�a�����Bf=�=��1	�=Y�=�S����<���=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�d�>���Z��q����u���#=1��>�9H?�R��'�O��>��v
?2?�]�M���k�ȿ�{v�j��>��?���?;�m�+@���@��y�>B��?eY?mi>�l۾�WZ�ƍ�>�@?rR?��>�9���'���?"޶?���?�I>���?g�s?�l�>$3x�7[/��6��S����V=as\;!e�>�Y>p���_fF��ד�+h��̻j�x����a>ř$=��>tE�g5���>�=���2K��c�f����>#*q>1�I>�W�>� ?�b�>Ϧ�>y�=�o��h‾[���Q�K?���?���_2n��T�<���=��^��&?-I4?�b[�u�Ͼ֨>ݺ\?k?�[?�d�>���(>��&迿~�����<�K>4�>H�>�#��sFK>��Ծ3D�\o�>�Η>����@ھ�,��RP��eB�>f!?���> خ=� ?��#?��j>�(�>9aE��9��]�E����>��>I?�~?��?�Թ��Z3�����桿��[�o;N>��x?V?�ʕ>Y���택��nE�BI�����h��?�tg?eS�?(2�?щ??\�A?8)f>���ؾS�����>�w!?����EF��	$���-�bR	?�?9��>-����	���#�7�R% �́?ߓY?�?���O*^���ʾO�=��N���j�+;�&���>�4>5�����=�>�f�=���A�{�=p|�=���>�Ĳ=x�K��f��,=,?�G�lۃ���=m�r�'xD���>�IL>�����^?Jl=��{�����x���U��?��?Uk�?���9�h��$=?�?L	?z"�>�J���}޾G���Pw�9~x�tw�T�>���>O�l���B���ҙ���F��^�Ž�~`���?>���>��?<Wu>T�>�\��?������>��I�e�n0��U���N��%���������Լ7��,����h>D�=�&�>�?�#�=�9>���>/��=}N�>��r>�>�}�>`|�>J��>��@>� ü22&��KR?#�����'�U�����h3B?�qd?�1�>�i�ǉ�����D�?$��?�r�?�<v>h��,+�fn?z=�>C��q
?�P:=e<�z4�<�U��4��/4��<�O��>�D׽� :��M��lf�^j
?�/?e��7�̾�>׽ ���(�n=�M�?��(?�)���Q���o�̸W�S�.���6h�Jj��O�$���p��쏿�^��%����(��r*=��*?j�?Ҍ����!���&k��?��df>W�>_$�>/�>)uI>��	�s�1�g^�
M'�I���eR�>{[{?B_>f8[?�J?!L?d�S?�,>'$ټ���W��>=8���_�>�+�>�92?KX+?s�??.�?b�8?yG�>��>�^�j�ξ� �>�N?��?f�(?7}/?����ݝ�=�'=�1�o�=��| >:�<(���,p(��$�;��=�D>�W?ߢ���8�	�����j>�7?�>b��>����!��`��<�
�>�
?Y@�>S���7}r�t`��T�>��?Y��|z=z�)>W��=V�����Ӻ�S�=�¼���=���w�;��3<8`�=��=�Br���T��}�:ev�;�<hu�>;�?���>RD�>t@��� �����e�=Y><S>6>�Dپ�}���$���g��^y>�w�?�z�?��f=B�=��=�|���U������������<��?�J#?�WT?	��?��=?�i#?>�>7+�M���^��m��n�?x#,?���>����ʾ��a�3��?G]?�:a����[>)��¾}ս߷>=]/��.~���_D�������������?���?��@���6�No辇���t[����C?��>^^�> �>��)��g�$�$;>���>�R?���>�q?^?�[:?А�>n���9��� e��o�m>�:N?�B�?�1�?�x?K�?�>2A����Y��Y=G�uw�a���~�=�7>��>�m�>�S�>���>����68,������*��>���>I��>�$?�U�>(Ԫ>^BH?���>�v��,3��ꣾq����UD��w?�j�?"^,?��=
��l�D�C���N:�>tt�?���?4�(?�M��8�=?�� ϵ�/s�_d�>z��>���>���=
zB=5�>��>@��>^��+G�	�4��,���?��D?��=�?���rj���޾�l����X�%�3�$Y�=6`F���=��¾�s�Z��ȇ��	�x���׾����J#�Γ���?A�=���<]�d<��ѽ��b=G��<n|�<c8z���*>�h�<`�<��*�~�f�n���1�=��=f�;p)���P˾�h}?�#I?�+?3�C?�z>��>�1�f^�>!���h}?y.U>\�P��H���d;��.��f���{�ؾ`I׾��c� ����>�H���>G3>v8�=��<��=B�s=�E�=5���H=���=_ �=H��=x��=�<>�p>�6w?W�������4Q��Z罥�:?�8�>s{�=��ƾr@?z�>>�2������xb��-?���?�T�?=�?Cti��d�>M���㎽�q�=M����=2>v��=t�2�T��>��J>���K��N����4�?��@��??�ዿϢϿ,a/>�-6>���=Se[�&�,�:���;7��#C���&?�4�����"�_>��=ɔ�	�ɾ�==��>tM\=G���qY�&��=�br�f��< �>=��q>҂F>j��=a̽m.�=���=a�=Y�%>u*G�`���Y�R��=���=�9>HA>�v�>��?*�?L~k?d��>��e�w����ܾ���>8ֿ>�`�>@ѓ>m%�>>n>[h4?*XJ?�U?�o�>��T>�@�>���>�?�DdS�����V��ƭ����?+}?t:�>�!%=~4��w4��?/�8W���?�]?\j�>k�>� �Q��J'(�Wi(���]��|�<S�f=Ţ��,L?�N�r�k����s�j�D>�>&��>+D�>t��>�q->-a>���>�,>o=�->�M��j�<���d̬=+��}ƈ���qx����<��e�7�>�2�n�A�����0e<�H�=_S�>�>8g�>3��=�ƪ�>�>f�O��v=�N|��I��|�%R���F��}��[� >l(e>��W����2c?��=*U�>ŗ�?��?Ax>�"!����e���e�>�w��?�=��J>r�-��#���4�z%P� ?ξ��>M>g{�>1����j&�K�P����=�����&�E]?b@^�T���~(�������0��v[����i��s>^�8?g�����>�v_?�Y?�Ġ?��>�Р��䛾\��=aA����0>2�)��׾N"<<�d#?��?_�>%���N?�{O̾*`�����>.I��P�������0����ἷ��w�>�����о�3�!b�����B�6Nr�W��>9�O?�?�!b�X��}QO����c����k?Mxg?'�>"I?�B?�����u�=����E�=x�n?2��?f5�?��
>���=Ȏ�����>�8?᭖?�f�?�q?ٸ;�_��>�:>;*�'>x[��}��=�>���=[�=�?P ?�
?�e�������<#Z�ó�<ME�=��>p�>�w>��=ۘm=�8�=
�Z>���>Ҟ�>��Z>X[�>p#�>wm���6���?�Ի���>�*L?w��>�jɼ+�u��X>��;>�J�����*����<��P5��<�@P=R�=�n�>�^ο��?~�L=J��V\?b��t6��*>eJm>*�¾>S'?��>G6�>�b?�:>Wf>Rs}>�>�KԾ��>�5��/ �ǘC�/>Q���Ͼ	C>�����(���	�CM���0H������M�/�j�i�����;��"�<���?����t;l�7q)�]����?���>�6?�ȏ�~����>r��>��>�T������Ǎ���ݾ���?��?�;c>��>E�W?"�?Ò1�/3��uZ�#�u�`(A�$e�M�`��፿�����
�H��2�_?�x?0yA?~S�<:z>M��?��%�Pӏ��)�>�/�#';�w?<=k+�>&*���`��Ӿ��þ8��HF>��o?7%�?nY?*TV����d�>�@?rg>?.�{?��1?�&?�&�~3?*�'>��?֝�>�~H?
;,?�B?T5]>�]>O�<�D�=�R��ט�	��~�/� 5�ڵ���	>��E�
�)�8�g>oҮ��V�<d�4��Z��1=�N=��G;�h�<S��<�N�>=�Y?{[�>J��>�4?П��26��W��?/?�q�9��?�����01��r/Ͼ�2W>��q?��?�<N?���>�[���L��� >���>z6a>y�>���>EZC��d:��Q��s->W�><�=�ʽ<nu������̱��%;>I��>R2|>N����'>�v���&z��d>C�Q�&���c�S���G��1���v��X�>E�K?�?֙=�S�F��Hf�3,)?Z<?OM?��?��=��۾_�9�O�J�9A���>A,�<�������u!���:����:_�s>t-��hOK���>k$�N�¾����#B3�.7پ�V>�׾�0ֽ9]ݾU�޾R���=�T>�b��⛎����� =?�Z=������Zj��Au�=��>l,�>� ��b����H���¾��=���>���>�밻~����M�6�	��i>�P?}`?���??wk�]�v�l�e��7��������=b�"?�3�>=�?��r>�X�=xh��=[�d<��l�S��c�>U{?"����+����7�J�!���>��>��=;�?�P5?�f?�i?��?���>��>o62�9����?��?��>�
#��/���8��t(��+�>�2??����?>�B?�j?B�&?ӖM?54?U]>�� �O�6�գ�>4�x>�@U�����-F>rwR?NY�>�uK?4�~?�!�=F��u�������=$/�=��.?q?��?��l>�3�>Px��D�=���>q�{?�>�?w`v?���=��%?y�A>��>�`Ѽ��>6��>��?��]?tUx?7DJ?s	?������߽V^���5!�P=�Ϣ=�;����=�~"=X�S�9ad=��+=Y��������l:�t�u;޺�;�U�Y�> �s>`���a�0>��ľI����@>;��GH��jʊ��:�=�=��>�?���>
[#����=O��>v@�>���w8(?�?8#?�;��b�:۾�K�:	�>�B?u��=��l��~����u�Íh=D�m?8�^?�W��/��/�b?8�]?�k�W=�[�þ
�b�و龢�O?��
?�G�Q�>�~?�q?ϳ�>��e��8n�<��'Cb���j�Զ=�q�>�V���d��=�>��7?xM�>�b>�(�=tv۾�w��s��?�?a�?���?s!*>��n��3࿔d��������]?�<�>!G���#?ɧ��R#о7�������1K������:���P��������&�-l��DԽ'ظ=[s?�s?��q?�Vb?Χ���c�֘_����IV��u�c��8D���C�S?C�8�k�w��=��1���ޞ)=mm�yz=�.�?�?� ��
�>B���1�������R>eǇ�%�V�	�D=�c��D=�<zi}�������j?�L�>-��>�Gf?��c�DI?��1K�%�>�����4�=�K�>7ɟ>�U�> Ἥ[����BؾJϖ���P��u>�c?<�K?J�n?�� �6�1�����!���I�<���iE>->�{�>۽R�����&��3>�>�s�f\�f��]g	�{�=�1?�|�>���>��?��?����쯾�\y�:�0����<!q�>��h?R��>�[�>��̽�� �q��>��l?`��>��>����fZ!���{��ʽ!&�>�>E��>�o>��,��#\��j��N����9�lu�=!�h?�����`�X�>nR?�:M�G<�|�>.�v��!�E���'�j�>�|?җ�=��;>�ž�$�k�{��7����#?]�?�_��X����>�K?r��>TȐ>w�?ʳ>P�����<�?��V?`0F?�~M?|��>�(X=a����׽f�?�7q�:�lP>y�`>v-�=���=d_�\Rm�=�P�ϛP��1�<����F�3<�~5:��<8o�= g1>�ڿ�ne�}d󾊗	�c�߾�|Ӿ��p���,�LW���l�������	⦾`M	�XK�_�d���>���1��EA����?�b�?h��c�J�����Q�U�~���|*?Ć������$��|�<���l_��ZK�D�L�{�c�-�A��	f��(B?ֳľ:ſ8p����뾹�H?�0?���?��jD�!��懼>��0�#D>�پKv��>�׿R�L�M?���>�;޾1�*��>�>���>Q�b>���J���>D!2?�A?��>��9���߿E߿��=u��?{�@[|A?��(���NV=��>��	?��?>�A1�pE����X�>�9�?���?�IM=m�W���	��|e?�c<��F�։ܻ��=8>�=�R=���`�J>�O�>4z�pOA��Uܽo�4>�Յ>hR"�����o^����<}]>��սsd��5Մ?,{\��f���/��T��U>��T?�*�>T:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=o6��{���&V�|��=[��>d�>��,������O��I��T��=�$��B̿T`��h!����=���<
�սV�X�)��M��5���W��:����=��=�>�0�>�={>��>#�^?�0\?x+�>T(C>��$2~��N���>Gw����V�C��\����z�����I<����Z���)4��M��[������0���I��l:�m6?��L>f�߾ �?�iN�;ef�9��&'<c��࿾�����f���?Lc;?ڋ���@�SN�:v><7�Խ�;W?��佫�����ߣ>�|�����<�ܟ>ҍ(=?ʾ!�'�M�N�Eu0?�[?�����\���%*>7� �&�=��+?��?ğZ<� �>�K%?X�*��9�Ye[>��3>oڣ>���>�8	>����W۽(�?��T?>��j���ސ>$`����z��a=.>+A5���[> ��<�򌾮,V��L���u�<{(W?ؚ�>��)���6b������X==²x?��?{-�>^{k?��B?�Τ<%h��3�S���>aw=��W?�)i?^�>Ї���	о.�����5?��e?,�N>Tbh����"�.�U�o$?�n?�^?�{���v}�]��z��|n6?��v?s^�ss�����{�V�x=�>\�>���>��9��k�>�>?�#��G������Y4�Þ?�@���?�;<f �D��=�;?L\�>��O�?ƾ�z��ك����q=�"�>���wev�����R,�^�8?ݠ�?q��>������=/�=#c���??$�?>��RU�<d��_�k�P7���J=�#�=�	�=�=���پ0���hp�����X��VX>��@��c�U�;?D���5#߿�߿�	���� &��?��w>��{=�"���>�W;<���7��e�^~���?�>�r>׬���瑾��{��P;����2�>'��؈>ȠS�����Ɵ��`3</�>l�>հ�>�Ү�d�#ʙ?�<��L9οٗ�������X?�T�?>f�?�^?�8<��v��b{�����G?�rs?Z?�%�rA]�
�8��t?x�:SW�M�P��E����>�??7G�>�-�nj>���>�?K~�<��:�,�Ͽ�צ�_��[ѹ?���?P������>~\�?!,�>�x
�ѡ���5�p���_�w���H?����I���5���C��ӈ��a:?/?<,n�,��`�_?&�a�\�p���-�
�ƽ�ۡ>��0�e\�K�����~Xe����@y����?E^�?Q�?6��� #�6%?�>`����8Ǿn�<À�>�(�>I*N>�G_�z�u>����:�'i	>���?�~�?Cj?핏�����U>	�}?���>A!�?)�=���>�x�=�y��%�@���">+6�=4}=��?�M?���>a��=o8�/��PF�{|R��J���C���>$�a?|TL?�b>Gm��12�?� �{̽t�1��@��?��)�%�޽��5>��=>t�><^D��Ӿ��?q���ؿ�i���r'�*84?���>� ?�����t����=_?�w�>�1�i,���'��JQ����?TG�?T�?M�׾�˼�>�>�E�>��Խ-'��劇���7>M�B?+�pB���o�y�>/��?}�@�ծ?� i��	?���P��Ra~����7�_��=��7?�0��z>���>��=�nv�ܻ��S�s����>�B�?�{�?��>$�l?��o�P�B���1=/M�>˜k?�s?[Ro���h�B>��?������L��f?	�
@}u@[�^?(�h⿃K��ؽ���iо���=:��=�d>�3��0�=A]K�TlA��I���y=��>��>���>�(�>:c>�,>F���^X ����R���:��������J������E��n��S;�{��iR������ͽ�Nٽ���|h�L�=��\?o�V?�=s?�*�>���$��=4����le�Uj	���=G֔>�=?�S?��)?��j=^��bum�������J���S�> '@>��>MO�>��>�E���t>[�>�|@>lM$>�ڢ=�
���=U�d>�>���>���>�5�>���<ô��L��ꥁ��1��PT��'�?��$��e��c��sR��K������=!rA?㚕=�Œ�9�̿C��%/1?V��!��X����j>=<?��T?�<>�̙��ѓ��D�<�_3=��0�%ؐ>��b����TA��g*>ݟ9?��g>�s>5�3��"8��;Q������{>V�6?"����y;�l6u�u�H��Jݾ�CL>�E�>*�I�b�s喿�g���h���z=�>:?A�?����ﮰ���t�?k���R>8C[>uE=�=�M>�?]��jý�G�}�%=LU�=#^>�?p,>�Y�=!w�>n���R�P��h�>Y4B>J!->�0@?�]$?[��Ж�p#��V+���w>*��>�`>a>HH���=3�>��_>��
�aU���'�A*=�@Y>W���|�`�ľu�9 v=1�����='�=b �X�<��t=�~?���(䈿��e���lD?S+?g �=2�F<��"�E ���H��F�?r�@m�?��	��V�?�?�@�?��I��=}�>׫>�ξ�L��?��Ž5Ǣ�ɔ	�,)#�jS�?��?��/�Zʋ�=l�}6>�^%?��Ӿ�h�>x{��Z��P��p�u�X�#=D��>�9H?hT����O��>�kw
?�?�\򾁩����ȿe|v����>��?Y��?��m�A���@���>y��?�fY?Tli>i۾r[Z����>�@?�R?��>�:���'�?�?�޶?���?��H>���?1�s?}|�>6x���/��M��ɋ����m=}Ʈ;v=�>.<>�a��\�E�_t��'��I�j�����_>��"=��>{��@����=�����䧾��a���>�o>�kJ>Q�>�?eh�>�~�>�=�h��|������G�K?���?w��N2n�dS�<�=��^�W&?�I4?F[���Ͼ֨>Ӻ\?N?�[?&e�>L��	>��迿�}��ȡ�<��K>r2�>KH�>� ��@FK>��Ծ�4D�+o�>�͗>[��?ھ*-���V���B�>we!?���>5Ю=ۙ ?��#?��j>�(�>CaE��9��X�E����>٢�>�H?�~?��?�Թ��Z3�����桿��[�t;N>��x?V?rʕ>b���񃝿~kE�3BI�<���^��?�tg?oS�0?<2�?�??`�A?|)f>؇�(ؾo�����>aU$?(�2��vM�؀��w���?¡�>�?}��17��B�<��^a�� �>�6Y?�S?� ��[�&�辞�==������+<;�ռ?���Td�=֒>��`����=1�=P�=pā�c���(#=�%>���><Z=��c�V��9@,?�HK�Hσ���=��r�"xD���>q�K>�'��I�^?�S=���{��������L�U���?���?�o�?`g����h��/=?M�?� ?B�>)����{޾���Ihw���x��k��c>���>�Mm�� �+���	���^L��Bƽ�*C�Ԁ?eN�>"��>�v?��>tf�>�����}!��k�Ӄ��s�y#C��+X��*I���u����,��+9=[�;g9��ֽ�>a̜��D�>6D)?>��=>a�>�A>P��>��q>��>e��>�i�>N$>�>���<�����KR?������'����W����2B?|od?4�>��h�(������?���?q�?�=v>�}h�f++��l?�6�>����p
?�]:=����<�X�����L(��R�C��>�G׽ :�yM��lf�l
?�/?FE���̾�Q׽�����n= N�?��(?�)���Q���o�ϸW�S�ə�j6h�Aj��H�$���p��쏿�^��%����(�kr*=��*?l�?Ό� �!���&k��?�vdf>:�>f$�>7�>uI>��	�f�1�`^�M'�B���FR�>t[{?D�Z><{K?!OD?�zF?bF?�;�=e�>�ƾ��>`5�=��D��r>��5?H� ?&T2?Z�E?�WO?I��>��=����V¾�>A�>93?��>�,?�>J�c�
�w�>h�=����6�Qg=����s�۽f�̻F��{��>jY?|����8�������j>u�7?�x�>6��>����7�����<��>.�
?�7�>�����yr��^��N�>���?���!�=��)>���= ޅ��Z��G�=�Q����=�߂��i;���<��=��=��m��$'�pa�:!�;�M�< u�>6�?���>�C�>�@��/� �c��f�=�Y><S>}>�Eپ�}���$��v�g��]y>�w�?�z�?лf=��=��=}���U�����G������<�??J#?)XT?`��?{�=?_j#?ѵ>+�jM���^�������?�!,?:��>����ʾ���3��?�[?!<a���;)���¾��Խ��>\/��/~�����D������������?���?A�?�6�~x�׿���\����C?~"�>�X�>}�>L�)���g��%��3;>���>}R?�>�>C�h?ۉ�?^�u?D�">��q�����a>���r�v>�`?�ʊ?H�?��z?0��>"�G>sF8�4����&�ն
��^�l�P��z��D=Q%T>n�>u�>���>�E�� ~�e��1ν;�ӎ=;��>���>f�?�I�>��&>G�G?8	�>���]s������΃��;�_qu?]��?��+?�w=�U���E�����X�>hn�?���?�*?S�S�N��=W-ؼ����m]r���>
�>#+�>��=_zF=��>�u�>�b�>���6S��]8�L���? )F?.��=������q�2����芾=`
�&�;��Z�U�=g8���;#�m�گ
�Z�̾>9h��چ��ó�E���K�x�j���zD?���=���<�>G(���)S;[�b;`BW=沌�l��<ay<=@
�<�3E=�*��
����i=�T=�/�oꃽ��˾��}?<I?	�+?��C?M�y>q3>�3��><u���??�V>o[P������|;�'�������ؾet׾�c��ʟ��F>�bI�`�>x/3>@a�=�'�<��=�ws=���=��P��=)�=�Q�=�b�=���=��>1W>�6w?W�������4Q�[罠�:?�8�>�{�=z�ƾ^@?��>>�2������{b��-?~��?�T�?6�?tti��d�>F��o㎽�q�=T����=2>j��=L�2�T��>��J>���K��$����4�?��@��??�ዿ͢Ͽ	a/>�KZ>K�%==e����e������Q��g,?�!��/�)^�>�i�=���Ծ)�W=���=�(s=0����]�L/>��"��^�<3H~=I�V>��=��=�H��̞=c&��F>�# >�u�=ñ���I�;�� >WǑ=;S>Vw?=���>Y4?��;?:vp?q7�>A����N���*˾�>��>��>>v�>��k>��>'p>?7]M?��Y?!DJ>9~>֏�>���>�T��U�$��?�q���^>W��?D��?.��>J��\�1��0�����r��'
? �?Z�>�2>�G�?��#��A�4�	4b�U��<�[/�"0���߼�N݇��)���a�?�=K��>.@�>u��>�q�>2�g>��j>��>�X�=��	��5�=Q3D;Uay<S��f�=?�۽=
e=��T<{��� �=����c�Pp��1�㼔A/�KI=���=R��>@g�=9��>7��=��޾�g>F����;Y��'׻�����W�0N{�u���W�N�'������=|i<>p�:J�Ȓ#?��=��t>���?��l?"Ϥ=����������B���1��k*����.>8K�R�'�?dA�wY��ʾ�A�>��`>���>��:=I��5M�1`.>И���J����>�Z����\�o�m�������(��W>k��S�=��E?غ�����>��T?5A?F��?fHW>�V�檾!>��羕�=V�7��E���bw�4�	?�%�>�>�>���:��G̾�'��Hշ>%AI�(�O�C�����0���+Ƿ� ��>�����о�&3��f�������B��Jr����>��O?��?4b��X���QO�������to?M|g?t�>�I?B?R��ov��q��^z�={�n?��?;�?B�
>�"�=�D���>;�?�-�?c��?�'x?��/�� ?���<�/�=�+�*Q�=
�'>Oz�=?�?>�?S�?�#?�Nƽ���h��ZپB!�?��=rB=���>s'�>�Qq>.�+>L�s=�_F=��T>��|>/��>\v>�Ƞ>fem>nҤ����� 	?WY5���>��0?��>�L�������&>�<E>�P���b\�V��x��sB>���p�!�=ސ>=g�>п3��?��<���? �����#3y>X�{>���0?�ޣ>�F�>��?4�>>�">�r�>/�AӾ k>��d!�F0C�9|R�'�Ѿ��z>�����&� ���u��#UI�/l���b��j��,��T8=�|o�<�I�?����k�M�)�l�����?�W�>�6?J׌����ƻ>���>"ƍ>�D��V����ƍ�pdᾊ�?��?�;c>��>I�W? �?ϒ1�?3��uZ�)�u�f(A�"e�V�`��፿�����
�b��/�_?�x?-yA?S�<):z>O��?��%�^ӏ��)�>�/�';�@<=y+�>#*��4�`���Ӿ��þ�7��HF>��o?:%�?vY?HTV��Aj���)>"�:?�1?�t?�1?�;?33�B%?�*7>��?%?�5?l�.?=�
?R�5>��=u4���)=�����	Խ�ν�����>=]�=41�97>)<�W=�ԉ<*��>�ۼ[�';�M���϶<�<=▦=F6�=a
�>�\?���>r��>*|7?i����)�����<�.?�K�=�������������>�n?s��?$6W?Aub>76J��sI��>g*�>��8>Ǿg>AW�>l��:�C�,r>=��>
��=5�X=�P�~o}�|��������=�7>L��>&3|>��ȹ'>hz���/z��d>�Q�ʺ�)�S��G�W�1�ցv�Y�>�K?��?Ω�=2\�+���Hf��.)?�\<?NM?��?0�=��۾��9���J��@�]�>6'�<���K���#��G�:���:>�s>.���k���>�N?�^Mž'����*�8�{���>}ࣾ �
�i����,澘v���e
�a>�=���!��:`��f調�G?�==�|����(���,R>=c�>��>���=�%!�'��w^žp#o=�#�>� �>sd�=�
�h_U�ݘ�V}�>��N??{?��s?�O��5����X����Xg�\�=c �>���>�?���>�q�=�Ğ��9&�S����]m��ֽ>{.�>%J��x��%�m���HM�<%�>|�?߄Ƽk��>+F#?�J?1�e?�s?F'�>��>��%���оC[ ?Y��?��>  ��}�z���H��)�Ǌ
?��/?�BǼY,[>��?X�?��?�N?d�?�IR>~>ξ�#�e*�>-x>byR�����x)�>��T?�
?5�t?�z?�y�z�E�+���j̛�n�>[�%=%"?�I-?�(?5�>Y��>2/�-��=�/�>V%�?F�t?ȞK?W͑>��4?a^�=�=D�½�>M��>y�"?�Rd?�Є?��6?'�?n�+�D���F�� �<�c�=O՞=����1�|�N�=^亽�m�=��P=�){:Dl;�9=��<��.�A<���V���m�>�Us>�Ɩ�r1>o�ž����XSA>�U��<s�����'p9�7�=|K�>��?9g�>�'$�H��=�M�>׵�>�H�N(?�?
�?��p:c�b�:Kھ�L�Ѱ>��A?�X�=i�l�D����u�qf=��m?bQ^?=�X�r��*�b?��]?'n�=���þ�b�#����O?$�
?h�G�H�>n�~?W�q?[��>@�e��8n�!��fCb���j�Aڶ=�p�>�V���d��<�>��7?�O�>�b>0�=w۾��w��s��?��?��?���?�!*>��n�4࿰]���E����]?�r�>r��#?���2�Ͼ�0���4��V��^�����[G���|��"�$�Aۃ���ֽ���=h�?�s?hCq?��_?ƹ ���c�^�N��P]V��+�S���E��E�b�C�}�n�H�m���C����F=h&Y�̺>�֎�?M�?�c����>�����}�ɤǾ���>��^�T`��m][��Mҽ!~=Iʽ�:��6������S?��>���>&�n?C�Z��<�3�5��Q`��i�L��=�:j>:��>۷?�2= �ż�m�<��վ`4��MRe��v>lc?��K?7�n?�� �G51�@���é!�*:3�\ ��#
C>��>H�>�(U�R��%��N>��s�&�(����	�.|y=��2?�Ԁ>��>g�?�?�	��᯾c6w�\^1��Ҋ<z��>)/i?�.�>�^�>�<Ͻo� ����>��l?���>Q�>����T!��{� �ʽ��>J�>���>B�o>��,�� \��j�����99��q�=��h?z�����`��>�R?	�:�H<�u�>�hv�I�!�O��4�'�~�>�?�Ū=�;>�ž�"���{��5���j?��?d""�u�%��>3�?�?�� ?��?�o>F��[�� ��> .B?��9?(�G??'|->qJ{=��z���P� j�>dU�>��#>���;Hk��N�9JK�q=w�<�\������3<�a)�G;�7L��dd>�LϿO�H����\J��`ؾ������������J��<t������Xþ섾F�,�ѕ��p�2��D�Kq�����o�?,`�?O�JL��U���U�u�2!
?����ը6=�"C��Y0þ��㾸:��V]�5�r�6h'���c���=?j����ƿ�ٓ�ZX侸D??��G?̀?Q���fI.����b�`>9'ɼ��>I������-�ݿ�4���[S?��>�P������a>��>�̶>�U�=\���W�=�>�JZ?���>ɯ|���3���D~�<��?"@�lA?̹(�dC�M�S=�<�>��	?�:A>u�/����u�����>Tߞ?���?�wH=�W�8/���d?��<a�F�������=���=�=�P�1�I>���>є�#{@�� ߽"Y6>�.�>{�!����^�o;�<��]>4�۽阽5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=s6��{���&V�}��=[��>c�>,������O��I��U��=Z ��>ſ`��O+���=2!����W�0����V�/�Wپ+���i��Z`�=��(>��>�_�>�c>I�k>�L[?�j?�A�>�>'�&���v�ǚ��eF=��=�
/��� ���=��5����뾀�����,�_	����L6�XTc=±W�҇���'�PW��H=���2?��4>p�ξc�C�d��:�;�E��%ױ��Z�@h̾��'�ik�Ç�?j�<?8	����N����T���X��3O?<��yR��,����=�ҝ��'�<���>%$�=�۾�71��bO�[0?r?���^#��8�*>�L ��"=��+?��?�(Y<���>��$?~�*���㽷�[>-]4>�L�>���>!
>��U�ܽ�D?uT?z� ������V�>����,�z�j�`=9N>A,5��/�H[>���<����>tY�Wq����< W?^��>�*�r�����d���#>=��x?G�?+�>�}k?}�B?���<%_���S��(��w=�W?i?��>�����о���C�5?M�e?��N>u�h�2��S�.��?��?{�n?�R?��0[}�������T]6?��v?�r^�qs�������V��=�>2\�>���>��9��k�>��>?�
#��G������Y4�Þ?v�@���?�;<� �"��=�;?B\�>j�O�??ƾ"{��܃����q=�"�>I���Uev����IS,�\�8?ܠ�?u��>;������X�>�%g�̂�?[w�?�=��!��<25��5{�a1�T�^>@�=*h�=��Ѽ�Ҿ�����Ͼ���~��{�/���f>u@��z����>�R�HK޿Zÿς��+��G��5\�>�`�>�ft>���myU���,��G^�oa]�`��뎣>��	>�ǽ̉��}�~�k5�a�׻���>kь���>�?I�j�����v�;	��>b��>��>�|��� ��Vz�?���s1Ϳˡ��݃	��W?�c�?`��?�?]mo���f�s"r�����+�B?z�j?6 W?�b�Cf�ӖF�]t?�>��B!V���T���A����>X�c?�Y�>�?a��?�=���=��D?/��bV��D׿8��)=��q�?Q��?�����>t�?c��>�������y���;B�@]����d?f_��$B�����F����t��E�?s-?��8�)��^�_?'�a�S�p���-���ƽ�ۡ>��0��e\��L��<���Xe����@y����?I^�?d�?���� #�S6%?�>f����8Ǿ��<ʀ�>�(�>*N>H_���u>����:�i	>���?�~�?Lj?��������U>�}?X#�>x�?K��=�g�>�i�=��
�-��_#>��=0�>�[�?�M?�O�>m�="�8�./�wYF�aIR�L%���C���>��a?�L?WKb>=���52�"!�eͽ�^1�4o��W@�ܡ,�ŝ߽j&5>q�=>�>i�D�Ӿ��#?�@���׿t敿��%��A?���> ?�� �	X�����<�a?w�y>ߩ	�n7���Ԑ�R59����?���?Rp ?�aо�N:;9i�=c�>��>$����µ�_`��g�S>�<?���M芿M�r�@XD>Hj�?|�@�ĳ?p_��	?��ZQ��K`~�����6���=,�7?Z-���z>���>��=Gnv�8�����s����>�A�?�z�?���>��l?L�o�T�B���1=�I�>��k?�s?�#q�󾫭B>L�?������_L��f?��
@�t@�^?���Z޿vm���6��W���#�=�3�=�l>���ǽu=��T�������%>A�}>��W>À�>��b>�o?>�S>\L���E!�uA���V��hA�x���D����^���:;"�T-��WT⾺��bD��E'���(���&��(�>�N?zO?�g�?���>��Y}������R=ؽ)�;*=D�>^P?C�V?�1?&4�=>E��i^b�Q�t��0��k؀��ȧ>�	f>ϳ>=��>Ϟ�>DG���l>�uN>ܼ>;�=`�v��������<�>�;�>���>�[�>]�>�^�=5������y��s�C���=,�?5"���O[�kf�����I�ľ�>C@'?�l�=G���|h˿1��
�8?���'�'�m�.Q�>@�+?^Y?��G>A�����<�.�=o�A��w"�F��>���ك�"�L�>��6?�g>�$t>E4�38�?tQ�X믾@�}>�A6?�z��&e;���t���H���ݾS�K>�r�>��F��p��閿�d��*h���y=nb:?�S?놱�s簾	�s��j��tS>0P[>��=��=�M>�;Z��wýJ�F��t#=!�=�E]>�Y?�Z+>���=֢>�M��֕L�·�>='E>��.>�>?]�$?�+�ꨙ�����Ee.�4t>Y�>���>�>�	G�u{�=���>8{a>�R
�5=������sB�zHW>�&��[�\�G�z�r�x=�_��w��=�Й=���"�@�82=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿx9�>/��>��ԃ��|���=O(�>�L?SW��,��J)��?9��>�����.�ȿ�dr�\��>�v�?A��?�g�����&�8���>?|�?��[?hfG>u]վg`��U�>�>?��M?�3�>������k?a��?R2�?sI>̊�?��s?�P�>�	w��{/��+������*�{=�{~;�p�>\�>�m���F����� U���j�k��a�`>�K$={�>gi�;���ö=��������@Zd��з>obp>W�I>k,�>� ?���>���>�=����쀾�Ж�t�K?���?����2n��P�<���=�^��&?hI4?Oi[�f�Ͼ�ը>
�\?t?�[?d�>G��I>��?迿1~��0��<L�K>4�>hH�>$���FK>��Ծ�4D�&p�>�ϗ>m����?ھ-���T��GB�>�e!?���>�Ӯ=S� ?_�#?��j>'�>�`E��8���E�&��>l��>|H?]�~?��?jչ�KZ3�j���桿�[��;N>��x?V?�ȕ>�������3�E��:I���Û�?)tg?�S�0?2�?R�??Q�A?�&f>���ؾ����]�>�1$?�&���K��� ��#_��?R�?�6�>��ܼ�)�4�<���p���U ?udS?��?t����`�Q�پ�o8=�x�ۚV<�H@<_�����>�o3>��>����=�|> �=bhv�j�/���>=�3�=�#�>X|O=�2U�PR½�C,?j�J��ă��=y�r��wD���>�L>A���^?S�=��{����>���E�U���?���?�n�? N��#�h��!=?7%�?�?�>������޾���#Aw��ax��[��%>|��>!�o����"���(����R����ƽ�#���?婚>~��>l�?��e>r]�>���x(�!_����<���x�b�9�a~J�E�6�c*��$��Y �"�>=0Vݾ�A����f><ex�0"�>�d?�6>r��>�1	?;� =z~�>�7�>�l�>7�	?�A�>G80>��>�ĳ<�a~��.R?����j](���GR��ZB?�jd?���>�b�6w���D ?~!�?�
�?��t>q�h�o�*�D?�E�>�h}��1
?��4=��M�v<���-5��>�����母>�ҽ��9�ȚL���g���	?�x?f*����;��ٽ�����n=N�?��(?�)���Q���o�ϸW�S�Ù��6h�:j��H�$���p��쏿�^��%����(�`r*=��*?j�?͌��!���&k��?��df>T�>K$�>%�>uI>��	�g�1�e^�M'�T���RR�>t[{?��>�E?�3?�LZ?�nA?;�>W��>\Հ��] ?�(8�6>c��>�G?r1?_38?>?�-?�0>�r��o����پݹ�>�a?Z�?��>�E?37��L
=/f����V����1��s�<aT'���*�2y3��Y$=	��>�U?x���8�:����k>(�7?��>)��>����&����<1�>ر
?�A�>� ��}r�`��R�>���?3��m/=��)>A��=腼t�Ѻ9I�=s������=����u;�� <i��=y�=@�v��_��`-�:њ�;�@�<�s�>��?���>6B�>�>��m� ����se�= Y>�S>�>Gپ�}��o$��[�g�Zy>Xw�?Yz�?��f=��=Ґ�=�|��iW�����#���n��<�?mJ#?�WT?��?��=?ik#?ú>�*�M��S^�������?.#,?&��>\��۽ʾ�񨿊�3��?�U?Aa�{���;)��w¾�)սJn>c/�j+~�x��AD�M��d���b�����?}��?��@���6�������Y����C?�#�>H@�>]�>��)���g��,��;>zm�>R?u��>�9S?Ni�?�ρ?4��>EP��V+����ܽ��&>m?П�?���?l&�?��>�_>�6ξ��)�V+?�s����h��ö�"g>7�=1��>���>�>P>fI>*���S�<!����u>�L�=��>n�>���>$[�>�,>>�]D?޳�>�E���l�nI��FK��M�
��Y}?��?�+?�Y�:T���;�o��E�>iG�?Eɫ?|+?X�I��*�=�+M��(þ�с� ��>���>K�>���=V�=�3=��>�C�>WS�b��8��3`���?"�D?Ǡ�=B:¿��o�|`���s����r�����V�ѩr��M�Pш=C���ۉ��K����]�_k��:��������Ӎ~�"�?�*�=���=(!�=�'<Ὧ��=ʆ=�F�<{��<�$�H�]<�4)�U8j��8���5<n��<#��<�f�O�˾�}?8-I?+?��C?�y>�B>zA3�ǎ�>�&���L?��U>Z�P�|}�� �;�ʸ��v��
�ؾX׾��c�{�X>5=J���>�83>_�=~U�<��=w�s=���=WH�^J=�S�=��=�)�=`��=$�>`;>�6w?B�������4Q�_罈�:?)9�>�|�=��ƾ�@?_�>>�2�������b��-?J��?�T�?��?�ui��d�>9��⎽`r�=����=2>��=B�2����>��J>y���J��*����4�?��@��??�ዿ��Ͽ�_/>��P>sg�=�la�:,������%�7�!��$!?$(��Xؾ�c�>v~�=�s��$ξK[R<4>Z�D=���Z���=�c�Q7�<�4}=�yZ>yE)>���=`/����=�Ԏ;31>u+>�T�}��7cE��\�=���=�>0�=�}�>W�$?�n<?�"�?)/�>�o��;ܾ"�ƾrt�>3%�>��b>p��='�>�)�>[P?�3>?}E?��>D&>3.�>�;�>�U��P��_���2����>e�?��g?�?3�=�䆾��(���/���=�
?�?CS?�Η>Z�	���)@����8�Zx\����q�0�r�"�l�z�#TϾF���j�!�=>;W>u� ?X�	?*��>�M>���>�B�>�i4>Ă5;¥���<i�!�T0߽R<>O�S�c,��+�������ս���=c��=�<�=�2'>N-�<p�d:	��=f?�>K>�<�>n��=�#ľ(;>G虾��_��P>��C�@�Y�;cy�2���
F��ˌ��C>��@>��=��ژ��S?���=Zsb>��?[{~?l�>�#��~���M|���w�hg����=�N>�6}��G(�(�>��J�ag�����>���>.פ>���=��$��TW����=�\�0Z�O��>��Y��T�Z�������D��r���7�_���p=�28?&���M�>�oM?6�Z?aL�?���>��m�d����,>:���/�>m�l�P����(<�?Jz�>���>� �spC��̾ۮ����>�RI��.P�����=k0��K�J����>����O�оg 3��T���ޏ�S�B���r��>�>fO?�	�?Tb�h��O���߫����?|6g?i�>�#?�U?ط���+�lQ��Kڶ=P~n?��?&�?��
>L��=��,����>T�>-=�?CW�?�`l?^a(�3�>�=�sU>��)��=7]�=�HB==��=��	?1�?�3?�ê����1�� ��Eb�&Q=�RQ=�Ǚ>O�>��y>�=Sc�=5f>�Ǉ>��>�_�>�[> ��>$f�>�@����վ#�?5�L��>��6?�6j>�>J����>�p>-���P��	��J☾�㒾��:���=g�9=���>�_ؿ颬?�M>���02�>b��=RL��F >���>������?,����>T��>zc>��>g/>[�(�q�þ���=���nP�AP��@7�������>r�\�'�E�w�澪���Vs�@g���%��g�t��iz�����pܼ#��?D�Ƚ&%����|���?B��>�t1?�Ac�:%�Q�X>�?ܤ�> ~�Mȏ�~��C�۾��?
��?�;c>��>F�W?"�?��1�)3��uZ��u�^(A�!e�X�`��፿����
�6��-�_?�x?+yA?�S�<":z>K��?��%�Lӏ��)�>�/�#';��?<=t+�>*��
�`�{�Ӿ�þ�7��HF>��o?9%�?rY?9TV��3���<>�9?'-A?��o?�-?e�,?�$���%?g� >qW�>�h?T�7?��.?��?d	4>�>{L��rE=�L�����&`���C��s�;t��[��=����bT<�n�=�fn�����i�f�A���E�>Ʀ<ޖ�=���=��>62�>+]?3Y�>y �>F@?��轤�%��%���9?=�ˮ���������*!ھ�U>�El?���?a�X?�m�>�5M�ɔS��>	�>�M>>]�v>�~�>�B���G��I=ߘ>>��=�[��t�Z8 �����3�;�j,>R��>:|>����r�'>}w���-z���d>��Q�>ú���S�'�G�
�1���v��Y�>��K?��? ��=�V����)Hf�,)?-Z<?vMM?#�?��=�۾��9�`�J�.C���>��<���鿢�|"����:�7��:ջs>Z*��.).��=��8��,;���!�`~���B2>�����=���`�8־���=a�B>53پ��3鋿Y񰿞�??d��<�g�����8���N�=���>l��>����4�G���5��|�E ��Vv?�O>a�<�
�T$]���!� r>�TS?;�r?{�?W�b�������Z��/�S�C��=�?�M�>fd<?�#�>[e�=yk���-������ao����>.�?��	[��Ž�u�X�E��|�>�7�>�2<\+?iQU?�?R�U?IW;?v�"?p��>Hu��ξ?k+?$��?��=�Fڼ� N�6�2�S�G���?��??�D9�w�>��?�o?	�?E@?� ?#�[>�2澿� �.1�>�c�>s�?��餿��>>�E?{��>o�q?�܂?Z�9=��M�ka޾0��/C>��D>��4?��?s?&�>���>pW4����=��?&n?[�?�H?�!>�f6?���=Z ?�K�I�>�#�>k<?�zc?
��?;�?Y�>s��S���z-1���ݼ��!>�S�=-\�=\��=I�=kۿ�ӭ3>6�T�9��=+�=���e����6��F���'��%^�>��s>���z�0>n�ľKK����@>iQ��0N���Ԋ���:���=��>��?���>�[#�ȼ�=Q��>�E�>����4(?��??�Q ;��b�0�ھ��K�-�>m	B?���=`�l�U���p�u��h=L�m?4�^?��W��%��P�b?�]?�g�=���þ4�b���龣�O?��
?��G���>[�~?�q?%��>��e��9n�����Cb�n�j��ж="r�>.X�H�d�?�>v�7??O�>'�b>z%�=�u۾H�w�)r��?��?�?���?+*>C�n�94�MK��BL���*^?�K�>���% #?h�&оv������9 ⾄˩�i���q%������F�%�-̃���ֽл=s�?Ds?_q?�e`?��n_d� >^��/���NV�-���[���E�K�D��NC��an��/�=����l���d?=_oy���L�JͲ?g?7�
��I?2�Z�/��3پ+ob>*��!�I=���=�!��BM�=�v��KT��+�jG��j�?ѡ�>I��>�0i?*�u��4V��0��$P�*��r-X>'�=��>l��>.�;�a��U��T��|\��2R��27v>-yc?��K?D�n?n��+1������!�3�/��d����B>5k>���>:�W�ߙ�D9&�lX>�t�r����w��	�	�N�~=�2?�(�>ƴ�>�O�?3?{	�l���kx�ԇ1�;��<{0�> i?@�>��>�н�� ����>��l?���>��>떌�mZ!���{�ŧʽ8&�>�>��>��o>X�,��#\��j��Q����9��u�=&�h?���>�`�F�>�R?'�:C�G<�|�>{�v��!������'�2�>a|?ǖ�=^�;>�ž�$���{��7����0?��?�ef�����0l>u4 ?��>���>.��?C3�>K���:犽�H�>�3V?}uG?"�W?mX	?3�=TU��:���,�a�շ�<�V�>=�> g�=�58>� ��c틾�Dk���b�y�5<$\� &����=���<��=���=y;>�ؿF�P���y����{��H�����]��MS�n���s$��/�����)�l��?��_�<�l��1���6*S�PrL����?S��?��ྠ=O����	f�Ku޾x��>�퐾�w��S���Ձ<`��E|��5��{�R��%6�H���^��:?�㾾�uſ>����[��?}aD?��}?_~�K�6�.�W�� �=�&�;詼;T���ܒ�M�ڿ�����C?U��>�ؾ_\�=
�c>F��>�S@>sx><����N������>��b?d?k���ʿ�����$����?F�@�|A?�(����&V=���>;�	?�?>[S1��I�E���aT�>h<�?���?�zM=S�W�I�	��e?|�<��F�t�ݻ��=�;�=�G=@��V�J>ZU�>��CSA��>ܽV�4>څ>�~"����]�^���<
�]>�ս�<��5Մ?+{\��f���/��T��U>��T? +�>Y:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?8ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=�6�+���{���&V�z��=Z��>b�>��,������O��I��V��=�T�>�ǿڱ%��U�m��;�a�<F�ow콪��;m�4��8�#�������܏>m>-�q>3�R>w�^>�m>e?��j?��}>�:>�*R�ZĈ�������=�F.��[o�"=t��fĽt�þt[�.��J�=���/����~{���I=�r�>=��V�j��P�#���\�>@��Q1?؅*>�;�Q�;�<�lž���$�p�0�˾�)�0j���?�>?������S�.I������豽�V?p:"��2 ��Ѡ���>�lƼ�E�;���>�N=�Ѿ�9,��2R�z�0?*�?�����`
+>�|���y=��,?�k?:�<v��>[P"?	m-���ٽ�-a>u&@>��>��>7�>[������2�?�T?�3���g���Ӑ>wNľ r}�iT=��>�8����O{T>���<�����oػT����q�<�(W?՛�>r�)����a������V==�x?'�?�.�>#{k?��B?�Ѥ<�g���S�0�pfw=��W?�)i?p�>/���]	о�����5?֣e?�N>�`h�z��g�.��U�$?��n?Z_?}t��vv}�F��:��dn6?��v?s^�xs�����Q�V�g=�>�[�>���>��9��k�>�>?�#��G�� ���yY4�$Þ?��@���?T�;<��T��=�;?k\�>�O��>ƾ�z������5�q=�"�>���ev����R,�f�8?ݠ�?���>������#��=Y���0"�?-6�?A����ǖ�G���,�����/�;>-�=E��=,�7=�<˾��i7־��� \���%�*f�> �@膽� ? �g�H��oֿ0I�����R�/�?��[>���=�E��g�m-���a�\�j�¾�Q�>��>8����葾Z�{�c;�oe��1�>�����>��S����ϛ��S*5<�>��>���>����ݽ�e��?�T��6ο*������Q�X?e�?$m�?&g?<(7<tw���{�d��*G?��s?�Z?39%�Y5]��l8�([v?��I���}��V�v�=��P?i�t>.��/.<�4��e�?��=�Af��oֿ�亿b�(��g�?G�?!K���>�r�?���>��	��n��4��yUU�x۽Ϭf?�_�>��ľV��Q}x�实�bx�>.V?Vfd��x�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?7$�>�?.r�=�a�>2e�=�򰾽6-�`l#>�!�=��>�)�?N�M?�K�>�Y�=��8��/��ZF�aGR�$��C���>B�a?��L?9Kb>���5!2��!�Yuͽ�e1�lS�hX@��,�>�߽)5>�=>�>�D��	Ӿ��?�q�I�ؿ�k��}'��34?�ƃ>��?�����t��q��=_?Gt�>B7��,��|'���l�d��?�E�?��?��׾�ʼ��>��>�=�>�ս[;��>�����7>8�B?J
�A����o�'�>x��?��@�׮?v�h��	?���P��Sa~����7�j��=��7?�0� �z>���>��=�nv�ܻ��S�s����>�B�?�{�?��>"�l?��o�N�B�^�1=/M�>̜k?�s?�Ro���}�B>��?!������L��f?	�
@}u@[�^?(�տ<.���}����I>x��=Em>��8�;&���k=7ݽ���@>&��>��R>`a~>9Nj>�[Q>g�/>J܃��%��M��1���N�=����R�Ud����q{����&῾"�оXӋ<c�ټ��@=m4"���潙ԕ���=��U?iR?��o?�� ?T ~�r�>]3��2Z=�#�2�=�"�>�[2?7�L?.�*?�f�=�0����d�>��v1��5����]�>��I>�H�>���>��>mi.���I>N>>,K�>�S >"�$=���5=��N>s�>5��>��>�	�>��<2����[���Q��_�2�720=>��?c箾�UD��F�����[;��bj>T�?��=Q���Y^ֿ�;���5?2���X��l~��(e4>H?;�f?�h>�Ҷ�e�݋�<��ҽ��e��=������'��gF��� >h�/?��g>�xs>�4�"y8��4Q�@��x}>1]6?����y9�4�u�t�H��	޾ yN>Ո�>��R��y�����p���h��{=�8:?��?!���#谾�s����m�Q>��Z>�h=���=x�N>sTb���˽�BG���$=-��='�_>�?V�.>h=�=�>�{���+L����>��H>?�5>�t@?Y�#?m_��8���D���)�w�}>�]�>�z�>�`	>�I��X�=E��>\�_>%��qWw�t����=��W>L���U�a�����Bf=�=��1	�=Y�=�S����<���=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�d�>���Z��q����u���#=1��>�9H?�R��'�O��>��v
?2?�]�M���k�ȿ�{v�j��>��?���?;�m�+@���@��y�>B��?eY?mi>�l۾�WZ�ƍ�>�@?rR?��>�9���'���?"޶?���?�I>���?g�s?�l�>$3x�7[/��6��S����V=as\;!e�>�Y>p���_fF��ד�+h��̻j�x����a>ř$=��>tE�g5���>�=���2K��c�f����>#*q>1�I>�W�>� ?�b�>Ϧ�>y�=�o��h‾[���Q�K?���?���_2n��T�<���=��^��&?-I4?�b[�u�Ͼ֨>ݺ\?k?�[?�d�>���(>��&迿~�����<�K>4�>H�>�#��sFK>��Ծ3D�\o�>�Η>����@ھ�,��RP��eB�>f!?���> خ=� ?��#?��j>�(�>9aE��9��]�E����>��>I?�~?��?�Թ��Z3�����桿��[�o;N>��x?V?�ʕ>Y���택��nE�BI�����h��?�tg?eS�?(2�?щ??\�A?8)f>���ؾS�����>�w!?����EF��	$���-�bR	?�?9��>-����	���#�7�R% �́?ߓY?�?���O*^���ʾO�=��N���j�+;�&���>�4>5�����=�>�f�=���A�{�=p|�=���>�Ĳ=x�K��f��,=,?�G�lۃ���=m�r�'xD���>�IL>�����^?Jl=��{�����x���U��?��?Uk�?���9�h��$=?�?L	?z"�>�J���}޾G���Pw�9~x�tw�T�>���>O�l���B���ҙ���F��^�Ž�~`���?>���>��?<Wu>T�>�\��?������>��I�e�n0��U���N��%���������Լ7��,����h>D�=�&�>�?�#�=�9>���>/��=}N�>��r>�>�}�>`|�>J��>��@>� ü22&��KR?#�����'�U�����h3B?�qd?�1�>�i�ǉ�����D�?$��?�r�?�<v>h��,+�fn?z=�>C��q
?�P:=e<�z4�<�U��4��/4��<�O��>�D׽� :��M��lf�^j
?�/?e��7�̾�>׽ ���(�n=�M�?��(?�)���Q���o�̸W�S�.���6h�Jj��O�$���p��쏿�^��%����(��r*=��*?j�?Ҍ����!���&k��?��df>W�>_$�>/�>)uI>��	�s�1�g^�
M'�I���eR�>{[{?B_>f8[?�J?!L?d�S?�,>'$ټ���W��>=8���_�>�+�>�92?KX+?s�??.�?b�8?yG�>��>�^�j�ξ� �>�N?��?f�(?7}/?����ݝ�=�'=�1�o�=��| >:�<(���,p(��$�;��=�D>�W?ߢ���8�	�����j>�7?�>b��>����!��`��<�
�>�
?Y@�>S���7}r�t`��T�>��?Y��|z=z�)>W��=V�����Ӻ�S�=�¼���=���w�;��3<8`�=��=�Br���T��}�:ev�;�<hu�>;�?���>RD�>t@��� �����e�=Y><S>6>�Dپ�}���$���g��^y>�w�?�z�?��f=B�=��=�|���U������������<��?�J#?�WT?	��?��=?�i#?>�>7+�M���^��m��n�?x#,?���>����ʾ��a�3��?G]?�:a����[>)��¾}ս߷>=]/��.~���_D�������������?���?��@���6�No辇���t[����C?��>^^�> �>��)��g�$�$;>���>�R?���>�q?^?�[:?А�>n���9��� e��o�m>�:N?�B�?�1�?�x?K�?�>2A����Y��Y=G�uw�a���~�=�7>��>�m�>�S�>���>����68,������*��>���>I��>�$?�U�>(Ԫ>^BH?���>�v��,3��ꣾq����UD��w?�j�?"^,?��=
��l�D�C���N:�>tt�?���?4�(?�M��8�=?�� ϵ�/s�_d�>z��>���>���=
zB=5�>��>@��>^��+G�	�4��,���?��D?��=�?���rj���޾�l����X�%�3�$Y�=6`F���=��¾�s�Z��ȇ��	�x���׾����J#�Γ���?A�=���<]�d<��ѽ��b=G��<n|�<c8z���*>�h�<`�<��*�~�f�n���1�=��=f�;p)���P˾�h}?�#I?�+?3�C?�z>��>�1�f^�>!���h}?y.U>\�P��H���d;��.��f���{�ؾ`I׾��c� ����>�H���>G3>v8�=��<��=B�s=�E�=5���H=���=_ �=H��=x��=�<>�p>�6w?W�������4Q��Z罥�:?�8�>s{�=��ƾr@?z�>>�2������xb��-?���?�T�?=�?Cti��d�>M���㎽�q�=M����=2>v��=t�2�T��>��J>���K��N����4�?��@��??�ዿϢϿ,a/>�-6>���=Se[�&�,�:���;7��#C���&?�4�����"�_>��=ɔ�	�ɾ�==��>tM\=G���qY�&��=�br�f��< �>=��q>҂F>j��=a̽m.�=���=a�=Y�%>u*G�`���Y�R��=���=�9>HA>�v�>��?*�?L~k?d��>��e�w����ܾ���>8ֿ>�`�>@ѓ>m%�>>n>[h4?*XJ?�U?�o�>��T>�@�>���>�?�DdS�����V��ƭ����?+}?t:�>�!%=~4��w4��?/�8W���?�]?\j�>k�>� �Q��J'(�Wi(���]��|�<S�f=Ţ��,L?�N�r�k����s�j�D>�>&��>+D�>t��>�q->-a>���>�,>o=�->�M��j�<���d̬=+��}ƈ���qx����<��e�7�>�2�n�A�����0e<�H�=_S�>�>8g�>3��=�ƪ�>�>f�O��v=�N|��I��|�%R���F��}��[� >l(e>��W����2c?��=*U�>ŗ�?��?Ax>�"!����e���e�>�w��?�=��J>r�-��#���4�z%P� ?ξ��>M>g{�>1����j&�K�P����=�����&�E]?b@^�T���~(�������0��v[����i��s>^�8?g�����>�v_?�Y?�Ġ?��>�Р��䛾\��=aA����0>2�)��׾N"<<�d#?��?_�>%���N?�{O̾*`�����>.I��P�������0����ἷ��w�>�����о�3�!b�����B�6Nr�W��>9�O?�?�!b�X��}QO����c����k?Mxg?'�>"I?�B?�����u�=����E�=x�n?2��?f5�?��
>���=Ȏ�����>�8?᭖?�f�?�q?ٸ;�_��>�:>;*�'>x[��}��=�>���=[�=�?P ?�
?�e�������<#Z�ó�<ME�=��>p�>�w>��=ۘm=�8�=
�Z>���>Ҟ�>��Z>X[�>p#�>wm���6���?�Ի���>�*L?w��>�jɼ+�u��X>��;>�J�����*����<��P5��<�@P=R�=�n�>�^ο��?~�L=J��V\?b��t6��*>eJm>*�¾>S'?��>G6�>�b?�:>Wf>Rs}>�>�KԾ��>�5��/ �ǘC�/>Q���Ͼ	C>�����(���	�CM���0H������M�/�j�i�����;��"�<���?����t;l�7q)�]����?���>�6?�ȏ�~����>r��>��>�T������Ǎ���ݾ���?��?�;c>��>E�W?"�?Ò1�/3��uZ�#�u�`(A�$e�M�`��፿�����
�H��2�_?�x?0yA?~S�<:z>M��?��%�Pӏ��)�>�/�#';�w?<=k+�>&*���`��Ӿ��þ8��HF>��o?7%�?nY?*TV����d�>�@?rg>?.�{?��1?�&?�&�~3?*�'>��?֝�>�~H?
;,?�B?T5]>�]>O�<�D�=�R��ט�	��~�/� 5�ڵ���	>��E�
�)�8�g>oҮ��V�<d�4��Z��1=�N=��G;�h�<S��<�N�>=�Y?{[�>J��>�4?П��26��W��?/?�q�9��?�����01��r/Ͼ�2W>��q?��?�<N?���>�[���L��� >���>z6a>y�>���>EZC��d:��Q��s->W�><�=�ʽ<nu������̱��%;>I��>R2|>N����'>�v���&z��d>C�Q�&���c�S���G��1���v��X�>E�K?�?֙=�S�F��Hf�3,)?Z<?OM?��?��=��۾_�9�O�J�9A���>A,�<�������u!���:����:_�s>t-������8�>ٮ-�W��+eG��e^�I���-���
�ݤn>f��Y�����U\>L�	>�{¾��%��A���ٞ���]?S��=,&���뜽��ܾ��<~!>d��>���=�y�lD)��ur��k�=�i�>��=�(��m���i8�'� ��-�>��H?�.=?��?��0�Dy���^�����T��mL)��P?���>�6�>�fk>~��<*� �e&�r|T�Ǧ����>��h>w�žY焿9���?�¾�yB�!�>6~ ?���>��>h�c?`.R?�/z?}$%?0?���>�ߠ�L�쾮;&?e��?fՅ=�xԽٲT��9��F��>�b)?�B�n��>Î?��?�'?��Q?�?�~>�� �}`@�O�>Jp�>��W��X��r?_>��J?���>RY?�ȃ?��=>��5�����t����u�=�>�2?�#?v�?�A�>���>򵡾4��=Ș�>Wc?o1�?��o?0��=B�?�F2>��>VӖ=���>.x�>`?cVO?^�s?��J?X|�>Rэ<�������Qs��)Q��|;��H<5�y=_j��s�/�M��</̱;�g��4׀������D������I�;-O�>{�t>������1>K3ľ|C��.�@>����p���튾�:�q�=wn�>>�?}E�>DB$�Ɛ=���>|s�>,�$(?��?oH?MR;��b���ھ�mK�z5�>V�A?��=ʼl��}��&�u���i=Ÿm?�n^? �W�S1���Z?]vX?�!ƾ��&�e茶���mv���P?��>����}�>܅�?�oy?�F?��4�a�g��3��3`��C��6�=�;�>����a��>}a)?�&�>�#>���=W�ƾ��埾�E?ً?� �? S�?�,>[�e�q޿����'ґ��=`?A�>�%���2#?���j1ξ����^_���ྀY���q���<���Τ�!�eł�I\㽉��=E�?��t?��n?I*^?�U �d?e�/�\�ɔ~�R�T�a�����/C���D��C���o���Ir��Z4��	i=rR�&�A�4��? K?1����?{ǔ��tԾ�'�ch>�N����5� ��==�����=�Զ=��J�V�j��ɾ(�?F�>r4�>.b*?cVW�d�J��%��-�u׾I+>k|�>��>"�>Y�D�2g�ԎL�@�ɾ�Ul��4h�Kڃ>3�`?�F?�}d?}���=�`ւ��7
�U���{���A>��C>W��>'���b�߽�\%�aB9��s�.������s�����=��!?�>>�j�>y��?A�>O��j���<��·3�����z�>�Ri?\ �>ςs>���I;.��p�>/�t?��>u"�>��~�z_���_�����@�>� >�X�>��>_u�ϴP��;��x����?��&�=���?���3�A�;�>sE?q,;iG=r��>��ѽ@�w�¾�/��Qn=�0?�=>��=.�����)ea�neڽP)?�K?&蒾��*��4~>�$"?��>�-�>E1�?�*�>UqþfE�Ա?�^?YBJ?rTA?DJ�>��=���x=Ƚ��&�W�,=	��>E�Z>�m=��=���ms\��w�U�D=ot�=��μ/P��~�<=�����J<��<��3>�ȿ�+�I��cy��N ��8�����핎�����? =/���F������q�2�'T�P�F���a��l{���#����?s%�?���%\ �n����������>=������=��־�|���̍�HaI�zs��"�%�q�^��w��-.R�E�'?������ǿ�����:ܾ�  ?�A ?�y?����"�Ԓ8�� >�D�<�7��d�뾧�����ο>���4�^?K��>@�J3��>��>P��>U�X>(Hq>����瞾�0�<Q�?ۆ-?Q��>�r��ɿ:���]��<���?-�@u|A?�(�(��9V="��>��	?��?>�G1�3H�� ���P�>�;�?���?^M=��W�a�	�<|e?�j<'�F���ݻ��=�#�=e:=���J>�U�>j���NA��Fܽح4>�օ>fs"����U�^��n�<d�]>>�սh#���l�?Id�yFa���B��j|���X>��=?�J ?-�l>��>6�i�,��&�t��x.?��?�K�?�K?ze~�B>��s�A?KjY?��?C,���t��u�>Lqh>� �(j��� �tv>+�>6>�� ����u�f���>��>� ���¿ %��Q�#��=�n=�o��ׅ1�z^E��O|;�k�� �J��pI��ֈ=NF�=�L>89�>��v>�T>Vg?6t?�F�>��>s���yn��-ƾ���2i��UYA�����CI?��!���y⾄��������{�����<�f��=NyR�[i��7o ���b�I�F�4[.?�#>F�ɾ�M�
�<��ɾ���3������U`̾��1���m����?�B?��!�V����c�U���mW?1��[�~̬���=�|���^=¯�>z��=P��!3��xS��o0?�n?�e���9��"=*>�� ��=�+?��?MT<��>�B%?��*�u��Z>�	3>?��>���>��	>l'��o'۽�j?�T?����g͐>[��G�z�ɫa=�D>@5�G�꼻�[>VΓ<���W��=�����<m�V?���>(�(������??�Ҽ-=�y?8=?���>"j?UB?�a�<�����U�6����V=`;V?rj?�%>㴄�s�Ҿ仨�\P2?%6e?2�R>ռg�r\�j-���z?��k?�?T����y�-o���0��8?�w?�6[�<1����.�#��`�?]�?u�>!��Jr�=?�,?,@�����n����'�.�?c�@� @#I�;%�\�F6|;�>��>A�v=�`��V��%Ծ@�=�Pm>g�=�`���;8�ۯ=�8?�/�?�0?p�辦>�"����?�_?����:=�D���[��{��G=��=Z�C�+�!�8E��{�.������豾l`��P#�>�4@��6� ��>�V=�2������-:y�����N���
?���>�R �"���ɵz��r��h�D�22�W �G��>��>����Sz��U|�
�;�@j��*��>��뼶1�>�N�s-��\����+&<w��>�8�>uڅ>�C��������?�����Ϳڹ����b�X?�w�?'��?b�?�� <�u�]i|���?��2F?m�r?(�Y?��IC[�pB3��j?�^��4U`���4�eHE��U>�"3?C�>��-���|=�>G��>Qg>�#/�}�Ŀ�ٶ�����5��?��?�o����>A��?s+?=i��7��[����*�i�,�~<A?�2>���M�!�%0=��ђ���
?F~0?�y��.�]�_?,�a�O�p���-���ƽ�ۡ>�0��e\��M��+���Xe����@y����?M^�?j�?���� #�c6%?�>a����8Ǿ[�<���>�(�>*N> H_���u>����:�i	>���?�~�?Sj?���������U>�}?m��>*�?��=�?���>�ɘ��С�mH>��&�Afj�bW�>x�?_��>m 3>h�Ⱦ��\��?e�9 �s˾��G���%>��>��Y?�Z�>ｏ�{�<�;ܾX�ƾ�����:>��1�1�����Id�>K��=�>�*0�����H ?3�tGտ1W���d�=�'?�lp>�)?L*��Cd�i��=[?m&v>ͺ��H��%���T�&J�?́�?9�
?��پ��CF�=-ۣ>���>�m�]������w>U�4?7t ��Ӌ�2y�Fr>�3�?�@�B�?�a���?r�
��w�y��X��4��C>+TK?3횾W|�=]�?�j>a~��ڸ�E�t���>�?�V�?G�>�b@?�_G��T
�:���Hd�>�ѕ?�#?�Q��[Q���"�7>����i����\?��@�E@[l?Pƍ�=(ܿ=g������E˾��a=\�=3W9>���њ=-�*=n߼M��G>0M�>Q]>�^m>)�U>M�<>.�+>d�����q����Ȏ��@9�������>�����X� �vJ �ȥ��)ԣ�Gd
���(c��E�B��6��[�T�>p�e?�b�?��E? 9$>襀�8?��Ӿ'௾Vu�=�mZ�:e?s�??v�?�w�?���=>���ڀ�����C�Ͼ�������>@g�>��>�H�>��>o_����=Rr�>i>[[2=���<���?��=�r>x�>�۽>���>�C<>��>Fϴ��1��j�h��
w�w̽0�?����Q�J��1���9��Ҧ���h�=Hb.?|>���?пf����2H?%���y)��+���>|�0?�cW?�>��t�T�5:>5����j�/`>�+ �~l���)��%Q>wl?�f>��u>º3��$8��P�����t{>4�5?�϶���7���u�¥H�(�ܾ)N>���>1H��s�%���\���h�K�{=ol:?C�?D���ా��u���<^S>\>�=7լ=�AM>a�g��ǽq�G�K	-=?��=�p^>BR?�+>��=Vڣ>:��"�O�ae�>e�B>>�+>	@?�%?M�㱗�疃���-��w>�5�>܀>�>�JJ�&�=�v�>ŵa>0_��i�����N�?��xW>'Z}�$N_��0u�&�w=C��F��=��=�� �`�<���%=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ#�>����Ԙ�Rƅ��x���<䃻>�K?���@�5�#��d
?t�?v�⦤��zȿ��u�F��>P��?.��?p�m��B��X�A�&��>���?��Z?��m>��߾��_�mg�>�=?M?�*�>���v����?f޵?>�?�Z_>}��?�wZ?;��>I"Y�|�*�ϔ���Eu��H={`ҽ�b>	>P��N�9��k�������|p�������>���<��>����r���9`=�$*<��������!��>!��>,�`>,��>S?���>�C�>���<�cؽ|�^���d�i�F?�я?�7����g��jp���E=�c6��"�>�,?d����ݾ|ر>Y8^?�s�?��a?<3�>�U�=A���¿��ž�4=�Dr>��>�!�> %��>��ܾMpY�*�>���>�m�;n�־y�l�*.=��>�??|��>E�=�1?%�?N�>���>�\\�g���T��� ?�O?��?E�?Y�?�睾��-����L��rX���>H5m?��)?�*�=�V��\��B��,w=N�=yK�?�R?ۚU��/ ?�e?U?U?b�=��S��d��%��=�?�>��!?����A��M&�z�y~?�P?��>�7��@�ս�Pּ���Y����?�(\?:A&?���,a��¾�7�<�"�N�U�~��;n�D���>w�>n�����=>=װ=�Om�VF6�%�f<�i�=z�>��=?.7��t���3?!�u���A�" �=l[�(#�Ŀ>��>������A?�����A������f���2۽ih�?��?.T�?���+<m��eJ?]�{?AS?�83?oYy���g��3	���P� Q�%<�>+��>p�9�]�7��������j@��u�̽����w?�˻>4)%?`?Z�>Uj�>@��E>5�j7���q澁�Q������3�Φ-�O,�j����7D���f�Ⱦ�����:�>��X�xz>VF?��.>��_>B1�>��8<C|�>��G>x]q>A�>r�l>V�$>�1�=ؼ�
8���FR?ͩ����'��������[.B?�^d?.!�>Eh�މ�����w?L��?�l�?��u>��h�P7+�Hh?fl�>�%��Il
?�X:=A��=�<|@�����6��"�����>��ֽ:��M�:Cf�op
?A"?!��[g̾+ؽ�4z�V��=d��?�^?
�3HC�d+^�`[<��HP�������y���R��u��狿��y��t���#��d�=�8 ?vq�?�0(�v�㾙���#�q�d�)���>��>%*=���>�[�>$�����*�@�q���C�_�����>���?���> �I?�<?W~P?dL?襎>�u�>**���=�>� �;$۠>e�>v�9?T�-? B0?9r?�f+?��b>��:����ؾ�?J�?G?�?��?�Ӆ��ýb���h���y�1K���
�=6;�<��׽�u��T=DT>�?2�=�V	#�>&־=>n)?��>�η>�)��Ū��_%�>��?���>\�#�qv������>�M�?�ۄ��RT=y�2>���=�K�=o�=�w�=!���^��=��+<�!�<�Q�B��=�9J>]R�;�0��~�V��b�=2����u�>(�?w��>�9�>*C��A� �����ǰ=�X>�R>��>=پ�t���$��u�g��y>�j�?�m�?c-h=��=��=÷���G������ｾ���<P�?OJ#?	=T?���?��=??k#?�>�3��L��!^���	����?.!,?ӌ�>��Y�ʾP񨿋�3��?�Z?,;a�i��8<)���¾��Խܱ>I\/�//~����+D�F(��@��~��i��?m��?�A���6�Nx�~���1Y���C?�!�>X�>��>��)�	�g��$��-;>y��>rR?���>�jL?'Et?!eT?�Xb>MC�ǳ���X�����#=>i�F?��?o�?f�|?��>�%�=m�5�������s4/���C&Z�S��<dM>���>��>���>]�=C����'���Q�C��=��><�>c_�>1��>��C>)J���~I?z�>j@��-�
��Y���"u���<7�?,�?u!$?���<|�)�*�J�������>��?_�?�p1?q>O���=K��<���������>QN�>H��>(��= '
<��D>`s�>%��>K�꽰��g�E�uf��F?�nJ?��=Fſ��q�8(h�&/��� �<�m��۪c�����\��f�=�ڗ����٧�[(]�����Ќ�����E���I~����>#�=���=�(�=!3�<�T�w9�<�XC=tQ�<4�=��l��u<��B�?r��ҏ��	Ի�F<44K=Ը�ĳȾ4"~?z�E?W1?��E?��f>GM>�3#��j�>P�D�?��P>@�k��s��+�A�ா���	�׾6�Ѿ��c�N��'">K�0�]Q�=Ɛ.>��=��<D�=LCv=�k�=�fm�R��<�B�=}��=��=��=e>^L>�z?vـ�JQ��3탿�+0�MOg?&=>)/=F'M��=3>c<->c��z�Ϳ�:�lCo?���?���?��?��c�GgI>O+��FqH�~*=��齡9.�����`=>�>��j>�1=��������=��?fp�?L?D���_�˿��=�7>�$>z�R���1��\���b�R}Z�@�!?;I;�1J̾7�>[�=,߾�ƾ8�.=��6>`b=@i�V\��=��z�Y�;=	l=,׉>��C>Ut�=2���=��I=��=��O>���^�7�]3,�k�3=���=��b>&>4��>y�?ba0?gXd? 6�>Un�lϾ_?���H�>��=�E�>���=sB>���>��7?�D?��K?���>ӽ�=�	�>��>�,���m�/n御̧���<��?�Ά?1Ѹ>��Q<��A�����g>��2ŽFv?�R1?�k?�>D
�#ſ�V�&^#��<�<`��>°�>D 3�g��=�|�>JS��h��7�o>�D�>���>�>Ti>l��=t�=�ì>�Y�=@���g�=���==f�;A�� o<=�=+�=�R=mS=���=���㽵���`��S��=E��<C�%>?��>912>21�>w�>����z�={�@��q4��L�=�M���V=�a�T�?d��1q)��J��\!b>���==�ɽ���@&�>�{�>��>�\�?.�|?�\��LF���s�?g��@줾�����o�>�eb=fHf���Q���|���w��2ܾ���>;�>�h�>6�n>8X*�1e>��s=)9���4���>�닾��ɦ�Yp�h������IZi�Rxκs%E?5���~�=�U|?nJ?{ӏ?���>�^��ݠ׾&*>
Y���}=ǚ�: s��%����??&?9��>b��#�D�Ho���ҽ�I�>�5�h�X������05�Q'$=D���a�>�R���N���n.�HX��ү���E��O�����>�L?�ҭ?�߃��Jz���S��4��-�v�	?Żn? s�>��>?����J����b����}=ưf?��?���?L�>s��=�X���c�>X%	?ܽ�?6��?5qs?�^?�=S�>@!�;� >x���3\�="�>Ӥ�=/T�=|l?k�
?0�
?Mr��?�	�&����GM^����<��=Ev�>Lf�>n�r>:�=4[g=�A�=�8\>Qڞ>bҏ>f�d>5�>�:�> �~�{~�H�@?��>��>�1I?ݻ>cO�=�%V��&�<��=�Z��D׽~^�����c�=l��;&ݧ����Mݏ>����┣?��>�V �qj?��)Φ��-�=馌>))��~��>:�?>��>J��>b=a>!�=��>���=�J���+�>lS�r4��o2�)3h�v���!�=Vd޽>�켍����s���r���M���\�HZ���t�m�'���=r��?	}����4��Z	�.~Ⱦ�
�>T�W>K;b?<m=�[��ie�>g�?��>��"���������Ҿɿ�?b��?�;c>h�>��W?��?�1�u3��uZ��u�q(A��e�*�`�l፿��
�o�� �_?��x?�xA?
M�<&:z>l��?��%�Fӏ�r)�>/��&;��?<=n+�>�*����`�ۮӾ��þQ8�GF>�o?%�?nY?lRV�f�m� '>?�:?$�1?�Dt?��1?j�;?�����$?1�3>�,?i?JP5?��.?��
?�2>-�=�xn&=�<�������Xѽ6.ʽ6����3=��z=jЇ�-�<;B=^��<��gټh�;Cࢼ��<�:=���=Q?�=���>"�]?�L�>p��>R�7?���w8��Ů�c+/?��9=?�������Ȣ�|��>��j?���?dZ?7gd>��A��C�>YX�>r&>�\>ad�>.}�=�E�_�=�L>�W>�ƥ=�XM�?ρ�4�	�����_��<�'>���>A|>O�����'>1%����y���d>�LQ�������S���G���1�ߢv���>0�K?c�?�1�=^J�h��VZf�2)?�b<?'?M?,�?���=�۾5�9�B�J��&���>G��<�������W��\�:�7g:��r>�-���R��k>}%��=޾�6n��K��'���=8����=�y���Ծ �x�>��=�'	>���� ��斿�����L?��i=W�����K��V��$�>vs�>G��>�f�J����(=�`9��9�=L��>7f7>ژƼ%!E�i�ў�>�F? ]?Lx�?�M��Ŗs� �C��� �/G���-���
?.��>k?[C>%��=���>M��e� *G�6��>`��>�l��uE��^��������%���>A�?T�>�;?	�T?�
?� `?��(?��?�܏>T1�� B&?6��?��=��Խ�T�� 9�JF����>y�)?�B�߹�>P�?�?��&?	�Q?�?|�>� ��C@����>�Y�>��W��b��=�_>��J?֚�>r=Y?�ԃ?v�=>]�5��颾�֩��U�=�>��2?6#?N�?�>]��> ���;�=ߞ�>�c?�0�?'�o?���=@�?�:2>F��>a��=ƛ�>u��>�??XO?4�s?��J?��>۸�<�7���8���Cs���O�5Ȃ;�wH<I�y=ؘ�>3t�K���<t�;Pg��3I�����$�D��������;�e�>��s>h���0>T�ľ�k����@>�]��_L��b���9��F�=���>;�?H��>Q�#�Rϐ=#r�>�y�>���G-(?��?��?(@F;c�b���ھ�aL��m�>�B?���=��l�o��Ҹu��i=�
n?�_^?��W�����sa?�UZ?@���]�8���ɾz�m�b��R?}�?��6�j�>ꑀ?tsq?���>2�i�|1q�dQ��zh_���M�%��=�ɗ>�X�k�a�L�>�5?*�>~�I>6k�=j�þ�(h��I���t	?(��?��?���?�| >��j�	�ݿ��羵ۓ�X�c?G��>�@��vv)?���@���s��{e��	y��v޼�2��͐��F����ڶ��4�2�=�?j
r?��s?��V?��g�e��eS��P����X��K	�U�E�+D>���,�*�k����l���!�@��h=Txz�e	C�vO�?X�$?v�*�D��>�$��-��QϾg�>>�2�����5�=�v����A=�qt=�g���3�:����!?9K�>��>�Z;?F ]���>���/���9�3���W(>�b�>ю>T�>��C<��2����=���)s�$ ̽I�u>{�c?��K?�-n?�� �2$1��]��'p!��2��C���XB>�>=��>&:S�h��+0&��s>�V�r�Sx��֑�k	���=.�2?Q�>q��>�Y�?�3?�	�����P}��}1�j�<�ú>�h?`��>�چ>W�ѽ�L!����>|1Y?�a>���>X_f�.���fV��w��mכ>���=��>Nɂ>��8�߀-�������-�'��a+>�u?+���"��ٸu>A.�?6\�=Cn�i>��'�'lK�� �����b7�����>�����>G���� �ʏj��=���X)?t&?����γ*�j~>�<"?�_�>e)�>�9�?�ߛ>�fþ˰ɺ��?��^?eJ?tA?Vo�>F!=����JZȽ��&��S-=��>��Z>o=l=��=�`�
�\��E���D=�e�=��ϼ�f��
7<匳��F<���<H4>� ο���=�	����͜Ծ+-��{Ȗ�����ou�����=ہ��������UԽ��Y��q��5��z��+�x�N��?ts�?���w��n��Wk��+D8��N\>���3�	=�z��gF�iƤ�������<��1B�=js�p�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >]C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾q1�<��?7�-?��>Ŏr�1�ɿc���z¤<���?0�@3|A?��(�r��2V=���>��	?��?>PE1��E�{����Z�>�;�?���?�iM=t�W�[*
��ve?,_<C�F���޻��==;�=7=���J>�V�>
���`A��ܽ��4>څ>p]"�u��,r^����<
z]>��ս�A���C�?��p��B�CvA��u��d�>�S?p��>=c�>Y��>�w;��!߿4���l�E?�t @�%�?<Y@?}x���gh>|뾥?�:$?���><�	�h���Ϡ>��H>\�4����G�G��4>yC�> .�=�!��S����V�N��<F�=��
¿�>4�3�'�C�=�6�=K�;�'�0����<K���|�/�H�ͼ�Ɵ=���=��4>@yk>�h>V�\>� k?�x?�ї>Zv�=�yB��*I�_�<�!y��ɖ�_lI�	�����ھnH�W�ؾ�F�Pc ��S	��N����<�$��=N7R��J���� �Kc� �F��,?��">�YǾLM�^[<��Ⱦ(���tĄ����H�̾u�1��Hn�0;�?��A?���aSU��H����nĽ�pW?���������$ �=�!���=;S�>Xx�=�Z�`�2�g�R�b�.?ب$?�ž������%>Gz���S�<\u?-c?���=���>�� ?��/�4@����=ML=w��>>F�>H�>��.ӽ�?e@?߭3��pþ�]�>�푾} ����=�X>"�Uv�;�g>��<�����c����/���<y�V?�f�>��)�����K��6���4=)=w?��?�n�>��j?^bB?���<î�aFT�3�����=��X?��i?ԅ>�1����ξ 5��6�3?�Qc?�R>c�c� x�j-�x�B�?*n?e.?a+���O~��+����v�6?>�v?�c��������.��H��>�>$��>�$��F�>I�%?��C��9����Ŀ"�6��b�?�e@�+�?�� �nQ'���M=��>n�>�*�&.b����$�ھ�E�=݁�>�^��1X��
0����P�L?�O�?H�?����������=�ٕ��Z�?��?l����Cg<O���l��n��5~�<_Ϋ=��E"������7���ƾ��
����H߿�̥�>AZ@V�V*�>D8�V6�TϿ$���[о�Sq���?O��>ӠȽ����A�j��Pu�X�G�'�H�������>M�>�	������~��w>������>��P��>��A�屾�R���:.<&Ռ><��>�^�>e/��St���Й?"n����Ϳ�랿[,���X?p�?7�?|s?��T<J�u� �����{A?�4o?��Y?q2�oU�15���j?NP��
Q`�ł4�$JE���T>�3?0W�>I�-��Q}=)x>ݥ�>8�>�/��Ŀ�ٶ������?L��?�p꾕��>z�?Rf+?�X��,���G����*�U{��KA?O{2>2}����!��=�j����
?�m0?���/���_?��a�5�p�	�-�r�ƽu�>N�0�%B\�l�) ��Ge������y���?8b�?��?W3���"��$%?�ί>͙���Ǿ?N�<���>��>WQN>��]�{u>D���:�)U	>M��?xx�?�}?��������!>�}?M6�>=s?�M>�Ъ>2��=����llI��:��.�_��>�vb?�?i?�\?G��>h�0�3�&�,p�[4W�ݱ���H�P�>�B|?oc? vZ>ƮW�&|�H?�2��X>8������Ab��￼�d6>���>b�>�\>������>� �?����Vؿ4;��wd,�#�2?�z�>q?k��Z!t������^?-q�>/N��7�����y���?8��?�B	?Yؾ��޼��>�u�>��>A�ʽ����������8>_zA?���-��O�p��>@��?��@���?e�h��?��%�Bㄿb���E��
��_N�=�<;?Kv��NM{>�^�>�^�<1Xk�kE���j��gn�>p3�?���?<��>�NT?N7A��+�-�k�N��>��?.U?�AϾ�#徫�=��=��X卿�+�P'U?��
@��@K_G?�񗿇hֿ����wN��[���l��=��=��2>?�ٽ�^�=F�7=N�8�
<��b��=s�>��d>q>6(O>�a;>�)>���E�!�r��Z���N�C�������Z�:���Wv�Nz��3�������?��4ýiy���Q��1&��>`���SIi?��?��{?�c�>����"?�����K�NJ>f&�=�1�>dK?FD�?��8?��t=L��5�t�"P����E���y{�>���>�ܥ>(/�>�J�>���
�>�/> 5�>��J<�3�=��A�5Z@�]�[>Ĥ�>x�>�{�>}C<>��>Bϴ��1��E�h��
w��̽/�?����O�J��1���9��榷�Sh�=Cb.?6|>���?пc����2H?F���d)�+�+�}�>�0?�cW?�>����T�?:>'����j�`>�+ �pl���)��%Q>xl?��f>��t>؛3��O8��sP�<��e|>�96? ���^9���u��H���ݾz�L>���>�k=��e��������i�W�x=�:?�P?ܑ��>���[�u�U0��RR>	s\>Z�=O��=CsM>:d���ƽ��G�~�,=wh�=��^>�U?Xr0>7ˁ=��>I=����T��>�pA>S;'>�	B?5*??���fI��*���#/��Bf>���>�&{>q�>�/P�qa�=�]�>м\>(9��ފ��m�e�G�SkA>�N�?�R�v�{��)v=ù���9�=bg�=���EXC�®=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿe��>�d"��u�������z����;�U�>��N?>�v�W�lz��O
?F��>���褿P�ǿ��u����>R��?���?`�o�*��JVC����>���?Ģ]?�e>���~P�_}�>�]5?h{J?���>%���A���?���?]��?�qP>���?/wl?��>�b#�Z0�Z���f����mV<��꼺6>��=�ٶ���A�����Q���жk��u�C#�>��=dt�>��y�о��'=i���r��q%��>��R>�A>��>�?�L�>j��>kx2=c,���t���c���K?���?L��e2n�GL�<˝�=H�^�,&?I4?�^[�^�ϾF֨>��\?�?�[?Pc�>b��I>��]迿:�����<��K>O4�>�G�>�#��JK>��Ծ	5D��o�>2Η>Q���?ھ+,��o.��KB�>ze!?���>�Ϯ=÷?�?.��=���>�:��z��1)(����>���>��a>s�7?�?Yy��[�/�{���L���;jw���=��?(0?�%'>�������X��9�>�6��+�?�x?���=W�=?wЌ?AG4?A�?{�>o/`�'����耽Й�=x_"?�M�9�A�� '�����
?�.?�/�>�~�E��ONۼ0�7F���?�^?M=(?19���`��I¾��<�a2���޹�&<\�(��9>�M>�[z��r�=��> �=�rl���7��M�<���=��>m[�=Ew8�G���v?,?gK��у��
�=D�r��gD�l�>��L>������^?��=���{�N
���k��	�T�1�?,��?`�?.(����h�a.=?e�?&?Gm�>�:��L�޾π�/�w��x�x�N?>9��>�r��G�я��'����C��G9ƽ���K�>��>�?2&?D�B>�Ν>� ����,�*a��z���[��C��7���-��B�U3���r<�?qƻ#ľTP��_��>�Lҽ��>�?~U_>�9m>:޸>�ͺA9�>�S>Dh�>�є>�	5>aV;>.L�=S[E�K^|�IR?������'�t�辪ư��B?^d?�L�>l;h�~������?V��?8h�?1v>@�h��6+��a?8U�>���le
?�j:=S)�& �<�>��������(��ߎ>&ֽ�:�;M��;f�y
?�6?v���_�̾Z�׽1ۚ��A�=�.�?�,?Um%��R�{xm���W�f�T�ٱ9���p��Ꞿc��)l��叿���v����'�oq�=��)?t͆?�O �x���ط���h���9�sr>��>���>��>��`>F���\1��]�W%$�懾���>�z?֙z>�]J?52E?R�V?oI?z�>MĽ>�;�����>�Z=���>R��>_�=?�3?r0?�`?܈)?pd>7
�qt��оH�?Ӊ?�`?+�?�?�k��푽�ɼ�Լ	Ad�S�v��?=q�<o�ｾ�S�dE�=�>6m? ���k8��%����e>�5?X��>��>#��m}���=���>�k
?�N�>� �0Ks���*��>V�?����7�<nE)>k%�=�=��� 6�=��=^�ɼG�=�p��Q
���P<�=�a�=�@;�#�hs��q�:��<��
?�U(?l��=?>���<3_V������ټۡ>������&=�ߚ�@/���	���*m�fm>�	�?Ee�?1~=4��=��>WѾ��þ�����ԛ�]D>�~�>eVJ?%Q�?C�?x�3?�;?Bק>0���ۤ�Py������O�K?P!,?ኑ>����ʾW�̉3���?�[?
;a�����7)���¾V�Խw�>$[/��/~�����D�=,������{��Q��?徝?KA��6��v� ����_����C?s%�>�W�>�>��)���g��"�>.;>���>�
R?3#�>��O?�{?��[?�T>�8��$��2Ǚ��GB���">�N@?���?2�?y?E\�>{|>s*�
E྾����( �@��p��ZrV=f.Z>�]�>��>�۩>��=G_Ƚ�����>���=��b>���>q��>��>Iw>�8�<o�G?W�>�n����y���^���X��Hs?Ϸ�?��&?��=�Y�^G�D���6#�>�%�?#��?�q,?p$X��_�=F���3���pr����>��>�m�>��=,yu=B�>~�>�P�>�]�S��8�CpU��?MH?��=%ƿ��q���q����Q+x<�m����c�C�����[��H�=����������`[�l����3��(����a����{��H�>�|�=i|�=���==��<M�ļv�<�nI=dM�<��=��o��X_<W::��Իp퉽�^���T<�eK=�)��˾֏}?nHI?۠+?�C?S�y>؄>u)4�Q��>�1��=?�%V>��O�Ob���W;�褨�����ؾ�~׾�d�$ȟ��D>I���>�L3>�e�={W�<8�=j�r=�Î=�4O��%=���=qH�=�d�=���=��>Kq>�z?�ʄ�DA���9}� ���|dn?�B@>�v��������>��=���J3���K��8�?gc�?W��?��>�t��
?{>�����1���	>u��=	�T>�<M�5=���>!=�Ծ,r����2�N�?IW@3>`?�|}���ɿLO}>�7>>r�R�`~1��\��^b�2�Z�K�!?�L;�U̾��>᰺=lB߾��ƾ>�.=m�6>�lb=e���S\�w��=c�{���<=p�j=�Ɖ>�D>�=##����=8IJ=��=��O>9���O8�o!,�k�3=��= �b>&>7��>��?`W0?zKd?�E�>I�m��,Ͼ�?��&�>�+�=�1�>N��=XB>7g�>��7?��D?N�K?]��>�c�=��>��> �,��m��T�f����5�<���?�҆?Iɸ>{S<O:A�Ú��l>�,xŽ)k?�R1?J?"؞>5A��࿑U+��3����H����)�=�"H�M]��/�9�S��$�=�K�>�M�>�?�>n�>q+>\V�=��>MU�>ـ!>��5�fd�<j��=��p=�4�fz=�D�<���=���J�<��K>�N&;%���b[!< ���1��<Ug����=�(�>W�=���>>�i>Y�����>�l4�yP�3a�<��˾�D�ǀj����r���Yν|�6>�=��q���N��>��>���=A�?$�p?�z<��*�f�侪���o���6��.=j��9�/R�x�-��'p��iV�ɾF}�>]Ύ>͟>�k>�
,���>�Vlo=�޾��3����>{䂾�I��)
�N�o����4E3j��=��"-E?�ԇ��{�=��|?
�G?���?���>r���d�ܾӳ >�v�y�<=[�>�o�HՊ�{�?+�(?=�>u�뾔,D��Ԣ��M=���>b/L���m��ԡ�_�@���S>vG4�dN�>� �
(����.���w����*�I��꓾p�>�"I?ft�?r���d-��`�^���Fs@<�/ ?�7\?��O>� ?1��>����>�
��;׾ˮż�i?���?z��?ٙ >=��=뵴��2�>�&	?6��?h��?zs?1�?���>ޏ;�� >Y����<�=��>�@�=���='s?A�
?f�
?	����	�g��Q��$^�!�<��="��>m�>ޤr>R+�=)�g=w��=P\>�͞>���>��d>
�>�c�>�*��y����?��s=@-�>��D?��=��l>�W,�{�ы;��W��dk��v���VT�0m!>�䁽Sk�Qƽ���>m�ȿJ�?�Y=3�1�?j��ȧ���<>�`>lĽt�>#��>[�>_��>��t>Z�>�c�>v�|>�(��c�[>H��N��S��b���'��P>,nP����Ó�Mơ=��ƽ�Q\�q����e���{�Og"���:XN�?+ ��$�8�B:��� ��8�k>��->�Ł?>�'=�"���{�>5P$?�]�:�Mܾ�ʒ��h�Ҿ��?n�?��>P�>ߖF?F��>��ɼ�W!�K�W�D�\��1f�������`��.����)������^?I�?|�H?9���<�>V��?Ge���Y�B�>2��[E.������>&���n��V�J�m ��q�s�M <�jJ?�W�?�l?,����i����>�Y�?-=r?�z?��J?U�?��w���?%�z>Ql�>YK?�tZ?ӫH?��? �=t�+>���=�<;,�#b��L�ڽ:ƽz��=�`�=�!�=<�==]���ҽh�}=�yݼ�Z�o��9�<#��<�v�=�>>vN�>��]?#��>%��>a�7?h���m8�����9'/?�^4=�R��扊������)�l��=G&j?��?w9[?%e>R�A�h�A�� >l\�>3$>�UZ>!��>u�뽢�A����=�s>|�>s8�=I&D�%/���
�`x�����<d!>Z ?�!>+���֖S>ڑk���)�G��>�=M���f��$Hc�W�H�ۄ��&��>}�F?0-?H ?>�N��2��3<?�W ?~�H??��=`��R-+�;?a���x�5�>�^O>�� ��S������s�A�����&=$ٵ����� �>����9¾��l��d�T����n<����9�=w���;X�J�秽=�Q�=���Re�{-������=�V?aN�=~����o���Ծ�l�=�.j>��>n��;�I+���%��N��R�=/�>X$>�@x����ZA�By�bń>�"F?3KZ?Ↄ?S�����w�V2F�s���!���՚��5?�x�>�
	?c�?>L\�=�ȱ�8���lf�s�H��F�>�i�>����G�[	���h��%��>e�?�>FB?\T?�b	?2�_?�&?� ?�O�>M?��뵾�A&?5��?��=��Խp�T�t 9�8F�k��>k�)?E�B�ݹ�>:�?ƽ?��&?�Q?�?��>˭ ��C@�Ô�>dY�>��W��b����_>��J?˚�>V=Y?�ԃ?��=>H�5��颾�֩�V�=w>��2?6#?I�?Я�>��>���o��=��>"c?+�?��o?xp�=��?#2>���>��=��>h�>��?BTO?0�s?��J?���>=��<�I��c=��*�s���Q����;1�H<�\y=�d���s�"����<�ɲ;�䶼�ր�O���D�������;l�>C�->�����]>�QݾM�s���n>���<��ž����H������%��>tz?A�>�@꽑(�=���>�o�>�@��C/?r?-�2?��p=l�f������L�>�J?�6�=�3t������u��{{1�S3x?)�Z?�k�����b?�^?�7��<���þ�Nb����׬O?��
?�bG���>b ?��q?���>� f��Kn����Sb�W�j�?��=y��>|*�V�d���>6�7?&�>��b>ޖ�=��۾��w�_�� ?/�?���?��?(*>N�n��<�`�����`�]?~V�>V���wU"?�b���Ͼk���������!���;��$c��=n���&$��ރ��0ֽ[�=�}?� s?�lq?�_?D� �#�c���]� ���V���0��qE��D���C��	o�����������;NJ=��q�A����?�'?W0���>=������;�!C>��������f�=*���c#@=��Z=�mh� p.�^N��� ?I*�>vH�>8�<?ȿ[��2>��1���7������3>�>d��>�T�>�0�:�d-�H,�R�ɾ�˄��vӽ6	X>�oo?H�d?{8Y?��q�/.m�Z?��4�|%���5>Z"Q>s8�>\T�{|��)+���L���}�	�)������}����=�M?��T>IPu>M��?���>���
���jҾވN�L�B="��>M�]?)��>-��>�����"�̨�>��O?(��>�[�>��-�r=��(k�2Ŗ��<?�@#?�?���>���,�Ψ���4��K���=�(�?؋��C�<�=1,?��a=��<={Pc>{'�<-l�Q�0��:V�ڝ�>�� ?�4���9(>�r��\���N��?�Z�YO)?�L?4璾��*��*~>�%"?�u�>f+�>�/�?;,�>ybþ��5�U�?��^?�1J?�NA?�Z�>:@=���@Ƚ9�&��,=���>E�Z>��l=���=���b\��u��1E=5��=�μ�V��ۄ<������I<ք�<C4>��˿�L)��� ��첾Zv��c8A�ɾꨮ�6bt���ǽ����Uk�J���B7�8�s������8��|����{����?���?3�y���6�PT���Ȏ�L%�&g>yy	�+O8�о?�g��6�@�ƾ�ն��V$�0�:��[���U�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >dC�<�,����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾t1�<��?7�-?��>Îr�1�ɿc���x¤<���?0�@�zA?��(����HHV=\��>�	?��?>�R1�=A�#���|Y�>a7�?���?F�L=��W���	���e?��<]�F�uYݻx��=/�=^	=�����J>�O�>���7FA��#ܽظ4>6؅>��"����Jz^�`6�<9}]>��ս�1��5Մ?,{\��f���/��T��U>��T? +�>?:�=��,?Z7H�a}Ͽ
�\��*a?�0�?���?$�(?6ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�҅�=�6ἒ���u���&V�n��=S��>T�>˂,�݋���O��I��Q��=�1 �Z�¿(�*�b���b�=�W0�pq������a������^��z�8�o׽�*O= ��=�wo>K�|>�r$>�o.>�X?��t?y/�>X?H>��὚����U��h�<y�+�/�8;�,��䚾Av񾶾꾗�	��9���)�����<�pז=hR�����~� � �d��G�Ve-?H�$>Eɾ�M�Oh%<��Ǿ���Z���A����˾%M2��^n���??;B?���Z�V����lc�eC½�V?%T��ڽ�����c��=�E��K�=r�>>�=r�㾃�2�8MS���(?�S*?OͲ�@a�Y��>��ͽ-;��?/?��=�w�>��$?��nǁ�M�D=w�>�b�><��>~��=m穾������?	�^?���=����"`>�\��𶊽�Z�=� ]�/��<ľ>�s�=\K���� ��m��J�=�\U?ٰ�>�y�������#�t�\��<Y�h?��?v
�>�q?��>? ��;-�辇�R�����:6=uY?3g?"� >�PG�h�ľ����h�7?Cd?U9>�ށ�~�پE�.�=7��?hDn?(�?��㼰Fq��ԕ�7�w�A?M�v?i^�h]��v����W��!�>�u�>y��>��9� E�>Hh>?,s#��Q������`F4��̞?��@�{�?-�4<�b����=�?���>�N�ž�ݲ������s=���>����v�N��Gl+�8�8?���?���>L���2�����=�ؕ��Z�?s�?J���}Ng<2���l�n��ۍ�<�Ϋ=s��G"������7���ƾ�
�W����ʿ����>Z@PS��(�>�C8��5⿓SϿ����]о�Uq�,�?G��>t�Ƚ������j�_Pu�Q�G���H������S�>.�>����"�����{�Ep;��ٞ���>��!�>w�S�?)��}���Y3<�ג>T��>�>!鮽�佾?�a���;ο��������X?e�?�e�?�q?AP8<��v���{����(G?O�s?�"Z?��$��%]��8�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�h�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*�F�+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.���a?s�o��s�[xm��_Ƚ���>�F��e���H���q����|�|鮿?�ݨ?�� @ɼ�?����VI7?���>à�Q�̾��
=m� ?h��>�܇=��>'��79�H19��O7>+� @v[@j��>nI��)r��.�>m!�?~��>���?�Ā>6�>��<>nd6���&��U�J��=I~�<G�?q?��>?��=#EE�N�E��7c�P�r����	K��ͯ>�&�?}�?�؇=3�޽�-�<;���Z�L����:�����S�=F��<���>���>.�=.�c�&A0���?q���ؿh���'�"%4?ĥ�>|?���F�t�;O�8_?�q�>�7��,��'%��|O�.��?�C�?��?.�׾��̼��>��>TX�>D�Խ$韽r�����7>ޓB?�B��E����o�+
�>��?P�@J֮?w i��?PN�^�z��1t��U<�(Y�����=Q?x ־z�b>:�?��<��w�填����?�>�F�?�q�?�I�>�;b?)`��,5�vZ���m�>��?�Q8?u}H�����">��]>�L*�L���b�:?��@� @��Y?b����ۿ)���H�Ͼֽ���2>��O>�J]>О�}f�=E��<O=k>��;93z>'��>٘�>|N�==�j>Vg}>�o��z������?��v�8��.�&]��������8�89⾟���ξ�:	����<=��%[��ԧ.�0_�;�U�q�?�?���?��>�]�����>#�T��B=���=%�-�!�f>��^?�|>?&�"?����� �ϛ���ؘ��z���C�R?kK�>��>�gr>�-�>�W{>J>n�0>Y`�>i�<��,=ଉ�1��=�Q�>'�>�u�>�t�>YC<>$�>:ϴ��1��p�h�/w�s̽�?J���&�J��1��w9�������h�=*b.?�{>���?пg����2H?F���D)�D�+���>q�0?ycW?��>�����T�v;>[����j�i`>, ��l���)��%Q>tl?+�f>�u>��3��d8���P����)d|>�26?�趾�B9�t�u��H��aݾ�GM>�þ>�(D��k�������qi��{=�x:?у?>���᰾�u��A���QR>t9\>�m=Wq�=�WM>�[c���ƽ�H��[.=߿�=��^>R
?�?3>�3�=�ǆ>aj��2	�Ff>r�
>�/�>Yv?�F?��!=�J���s֊�����>���>�r�=��9�7��=_�>ET�>��	>�:��f�dEY���>$�<^��}�k��*>�9���>K�4=�P��Ǝ�ioS>Ѭ{?)ɢ�W$s��Q4��EV�=nh?���>3
�>�}��Z�޻��N� ����?��@P��?�$���I>�.,?�?z����=F��>W�>t��*j7� rO?�f�=�#���	����~k�?�։?TT�c�o�IEk����=�N2?��^m�>���IH������#v��=k��>KiH?r���#�O�,x<��u
?�?�R�¬��Q�ȿ�v�G��>D��?P��?�&n�K+��Q$@�!��>���?�Y?<�j>Ll۾:xZ�0}�>9Q@?�Q?�]�>�W��&��?1�?$��?&I>���?��s?�o�>�Rw�M/�</��В��KC�=x�l;zq�>_X>E���D_F��ԓ��h��,�j����x
b>�v$=��>�$��)���S�=����@��.g�'��>��p>��I>X�>�� ?"[�>
��>f�=ˋ�[ꀾ ���o�K?���?����2n�#O�<���=A�^��&?{I4?�i[�X�Ͼ�ը>�\?d?�[?�c�>Q��R>��H迿R~����<��K>V4�>xH�>5%��WGK>��Ծ�4D�cp�>�ϗ>a ���?ھ�,���M��DB�>�e!?���>�Ѯ=r� ?��#?O�j>g�>XE��1��-�E�#��>O��>xZ?a�~?��?�ع��P3���衿և[��PN>��x?�O?���>ń���z��DE�G�H�,쒽��?`qg?��U?�+�?e�??	�A?�f>����ؾv���&�>��!?��úA��N&��	�g?�Q?,��>x;���ս�zּ���}{��O?I)\?:@&?���i*a���¾H0�<�"���U�4\�;��D���>�>Q���Y��=�>�հ=fNm��G6���f<�n�=P�>l�=�+7�Ux���.,?�AE�)����Κ=��r��]D�ŏ>ӰK>/t��s^?�!>�� |�)����g��
LU���?Gt�?V�?�n��֕h��=?�?��?��>�V���A޾�Qྔrw���w��o�U�>-��>��x��g�ӟ��r����C����Ľ:���#�>5�?�?�0�>�5�={��>st�uaY��}���#.��v���M�(���:��/��־�5��m>��� �,�R`�>�Q�5ZE>k<�>�6�>�q�>��>
摽(�z>�{�>ɻx>M'�>u�=�"=}��=�R,=-NM��sR?����9b��������K?z�y?W"?pP?�h7���w/�F�>O��?<�?��>� Z�K���O?�+�>Z�i��?�O�=qF�>Ï���Q���T-�+Py�9c��p�>��!��H��3E��e����>��?�?=�@����:<C���r�p=>+�?�F)?�)���Q�d�n�GW�5�S����l�`��e�$�j p����H������i(��`2=��)?{��?@� ����罭�
|j�j�=�V6h>�0�>K?�>�5�>�K>����(1�bL^��(�����W��>�){?���>��I?��;?�|P?%�L?���>M2�>���3]�>xY�;%�>.��>�9?7�-?�0?m?�s+?9nc>7%������twؾ9�?��?�O?�?�?��ֱý�ٚ���i��z�<W��#`�='�<G�׽�u�,:U=lT>�c?+���8�r���Zj>E�7?���>��>m��3偾���<|��>�
?{܏>IL��Wr�3�9��>�y�?���9�=ϔ)>'l�=����Ӂ�;��=��ļy��=Cc��9h;��E!<a��=Đ�=w�I��R��;��:�˖;���<0?�j'?��>�F>I���׽[�?ھ��=�Az>���>�?{>_���<��wP���Wz�(e]>���?>٥?������=�v���p�q��4�"�Ӱ��������>�Z?l��?��?B?h��>8�r>4U�������.�0z���e�>f!,?<��>���6�ʾh�	�3��?[?m=a����<)�~�¾��Խ��>RZ/��.~�4���D�!?��j��Jx��ћ�?���?�A���6��x辅����\��?�C?y!�>�V�>��>��)���g��$��0;>o��>_R?�#�>��O?�;{?&�[?�wT>��8�p/���ҙ�"	2�	�!>x@?���?���?Ny?�m�>��>k�)���>P�������܂��:W=�Z>~��>	)�>�>���=�Ƚ�y��f?��m�=ʏb>4��>���>j��>sw>̙�<PE?[�>���DAྒྷ���c�q��:=�Rp?��?�\?� �:ɣ�NO�!G��o�>�P�?{��?�!@?$����e�=洕<�iݾ���� ��>U��>O�U>>�>���=h�Z>���>�M�>�@��b���=�V}���!?��<?��9=��ȿ�t��]��M@����<�ߑ��E���w�t�U�k,�=a��|����p�T�c���!�~�䨹��̨�H~���>��=���='Z�=V��<�AA�YG�<���=�d0<:��<���iN)<"�1���f��z`�{��<��=.d���)��3ހ?��L?s>?�_?G�?>L��=��9����> ���i�?D�=>����Ⱦs�/�s���s���#��ە;��C�6���4�>AK��>�ET>Z�=�Ac�2"�=$�<A�k=̃��J�<kV�=y�=]�=z��=�(>L>��r?n"���я�+�u��㷾�p;?�7�>��F=sꃾ�?I`w=�0��cl���V��t?z
�?j��?�?!����[�>�����G�Q�7���">�(�>�R�� ����>�墽��K��:����ڼ��?`w@�S?ì���ͿO�N>��:>�^>liQ�o/1�([�	mZ���\�cc ?�(8���Ǿ
�>�<�=�ᾞ�Ⱦ���<g�6>��=�4�O�[�2)�="�|�\�4=_Gk=~D�>��C>7�=P˷���=j�Q=6��=p�T>�mһ7�2�3^)�9\'=��=�:_>j)>���>�	?��/?�Qd?p�>��l�*
̾�3��;Y�>���=��>��=��;>6��>@S6?a�D?�kL?���>!v�=���>�ݥ>iA-��qm��3���d��<�?Ӎ�?���>8݀<�4=�Ң���=���ǽЅ?�v2?h�?bě>����ɿ�^��_%���=י=��>��"�m3��,�<���=s�>Ө�&Xv>X�
?+;�>��=5�h���=���>z�=�߽�	�=�x=��.�~�սm[>�.��;b=�Q��AW���= =/��ۃ��~=���="|4�U�B��~�=c��>I�$>Z�>���=WS��_*)>���r�U���=cv����K��b�M�y��z,��t2�Az.>=�\>C[G�.|��0?���>g=>s��?�3h?��!>���G�Ծ�g��=p�:lA��=_�=X.s���H���e��P��������>�>v�>��l>��+�H?��=w=�%⾶L5��(�>�Y��������-q��;�������i�y󺻩D?�B��/Z�=�~?X�I?/֏?���>����|ؾ�/>����&=�����p�𘓽��?
'?��>�D�t�D�����Ӻ��|E�>�<!��
y��̞�4-�$KM>�ogn>I�3������$��r��g���J�����S�>8�C?�n�?������|�'E��L
�N��=�%?��[?:��>��>C��>T�!���۾��g==�?6��?�S�?��=��=@Ԁ�tf�>T�?�K�?���?~k?$@G�IF�>�黹�*>����Ѽ=�n�=5�q=b8�=�Z?��?�|	?�����6�%��a:���/���i=���=7v�>�@�>I,�>"��=B�f=Sq�=Çg>�c�>��>��h>5ڡ>���>�6�������$?nk�=Q��>=1?��}>�9=�æ�m��<��.���@���0�2�ƽ�+�kg�<ӵy;��{=<���[d�>��ƿ�ٕ?��?>É�"?�%=��5Y>�b>�Dֽ^��>��<>p��>j��>J�>�>U�>j�!>Ѭ�Z\>;}	�p��#0_��c����1�ohc>z�2�Vk��[S���-<!l����A6�Ph���|�-�@�-T����?�r;�a0���0��|��+/?�pn>�pi?�L�Yq ����>�?��=�,�U����q���m쾗>�?Ϻ�?���>�b�>��O?o�?I�N��H;���!�X�Y���A�Uke�m�Z�d7���̀����|9ܽ<TV?"hv?�Q?:ڨ�\��>h�p?��M�f�h�h��>�<�95+����=�K�>e��}̽�홾s5羦zw�$�_>�؂?&�?85?�P��Tan�$�'>��:?��1?�Pt?��1?��;?ݢ��$?G�3>�F?�d?Y5?��.?0�
?F-2>��=�Ʒ���%=�����H�нjʽf�nc4=2;z=�+�9��<um=9�<���ټ)�;���-�<u�:=�#�=�*�=��>��d?���>��>3�M?K޽�a/��2����#?YX=��ý�y;���ƾ�)��e~�_�K?�?��^?9�4>��%�R8�̫�=��>�'P>�2H>Ʃ�>��/��!���(<��>!��=*6�=_�[��8�8^�����l�=�1?>X�?Q�/>�px��X�>3����u�*{>�L5�9H
�����n�W�aX��Z�v��>�=?��*?�|�=f��2s�<�c�E�3?��8?.�B?@
~?���DL徢�@��=��L=��v>p ؼ��9�o%��I����V4�������>���uז�d֐>�Q ���]�t�X^�<�ﾽ��<���<M�=14��־\48��t>d��=mĹ�WI!����������X?썎=I.���gJ����<�/>ZZz>Ǐ�>}U1�b���@0�|"e�i�=��>��!>*\�B��XAB�'$�@�>�PE?�S_?�i�?����s���B�����Rh���gȼ,�?�j�>�b?�B>��=j���(�b�d��G���>��>��h�G��<��G$��_�$����>�4?�>b�?D�R?��
?n�`?�*?�B?�"�>���
���B&?懃?A�=o�Խe�T�2�8�9$F����> x)? �B����>��?V�?0�&?4�Q?��?�>�� ��I@�В�>\�>�W�Ca��?`>��J?���>�5Y?0Ӄ?��=>Z5�آ�~ʩ�>�=�>��2?3#?z�?R��>O��>󬡾+�=��>�c?�0�?��o?�w�=��?�22>a��>o��=���>��>?�WO?Q�s?��J?���>q��<c8��h3��*Ms�[�O���;wH<C�y=���:t�c7����<���;-m��4�����D��7��;%��>�gm>�h��X31>��ľO틾�d=>G$\�/���Ǎ�-E�!��=%��>��?H��>��vҏ=��>gn�>dZ��>(?.?��?���;�c�u޾WP��>@?��=�^m������jv��D=9m?��^?�V�����R�Z?XZ?/�;�0����|l��r����A?�'�>��z��>%��?�jl?���>�"���Ń�����6y�ƅ߽�.����>)]���Mb�/\�>��?-��>��x>j��<��ܾ��b���m���?�ɉ?H��?TK�?��T>��w����N���K��)^?0��>�?��& #?����-�Ͼ3P��f(��⾙��A���B���x��}�$�ރ��׽��=y�?js?�[q?a�_?̳ ��d��1^�*
��=kV��(�&�7�E��'E�őC�b�n��b�0��#����G=��~�͐A�R��?��'?E�/�؛�>����I��'3;��B>$����J�#�=u㋽(T@=�_[=B8h�TU.��4��
 ?e-�>Y3�>��<?�[�">�ٞ1���7������3>��>���>�N�>�G�:�e-����rɾ�����ӽ\�u>8�c?y�K?�9n?3&��A1�E ��l$!���4�s��@�A>��>�d�>��U�Oc���&�*�>�7hs������cf	�>-�=.�2?X4�>q�>�K�?(�?�#	�I�����z�t�1�j�<�L�>�i?���>��>�ͽ�!��F�>�LT?���>��|>Y���_!�5up�L���`�>k��>O3?��y>����A�y���n����X�:t]=!��?�����.E>��8? *>�E���7>��-�, $�ړ��'���>�>�X?:�/=Q8>U᭾�A!�R���z�P)?�J?�撾�*�,3~>�#"?~�>�.�>�/�?�'�>�rþ�JM��?��^?BBJ?�TA?9K�>,�=���O<Ƚf�&���,=���>U�Z>�"m=/u�=?��Sr\��w���D=�y�=�μ�Q��*�<���zK<��<��3>�Iο
1��[��]��̾�&�Z���Z�1�?z%�["�<�®���x�A��U#�ߗؽ9�=�0rS��g����Y�8J�?�@��!?��'����Ĕ��
�q�>���Z�-�%�k�Ɗ����þw����d�G��\����x��'?W�����ǿk���Ձܾ��? ?�y?B���"�8��!>^��<����>�������ο������^?��>`�5�����>�|�>|�X>�Hq>l��Ӟ��!�<�?J�-?�L�>'s���ɿ·���r�<���?5�@�WA?�4(�f�]Z]=�K�>?�	?4|?>��3�$��4��N��>���?�x�?*�B=��W�����e?--<��F�m���=<��=��=�����K>���>�T�P�C����,�6>�$�>�^,��E��\��<��\>�ӽ���	��?n]���d���0��u���>��U?o��>?��=e)?��J��ο�-[��wb?3��?�'�?C&?�<�� `�>.>۾��K?��5?�ݝ>��$��|u����=pܺ�
�N�S��A�U��s�=|��>�f'>�O-��J�u_U�{Mx�d9�=6 ���ÿ�h,��	���V=�T`�_q.��n*�7���f<3���k�ϒ��oz=*��=a8M>`��>�T>�e>�l\?tz?X��>���=rh��ޱ��Nʾ�민6�]���	���w�z�������/�۾���.}�������ͭ4��w>}h�����=%���|���C�� ?�OE>;���8�R�7�.�6g���P���{5�7���.;'u;�vFt�Q_�?��W?�S����M��l3����`�ҲM?S}齒�������->��=���=�W�>x�`=���T�?�6�W��0?),?l���ZB��K)>� ��C=n+?W�?w y<���>~%?�r+�����Y>��1>���>��>~h
>��-�ڽGQ?�T?��w���#|�>ڷ����{���g=c�>YG4�?�[]>k�<O0����{������E�<a�T?(m�>������H��%r���p =w�[?џ?�;?{�o?z*?#%��-�о��^�<�@���Q�ҸU?��z?���={}�9�߾�܋��b?̟2?�o>�>��� ��i��R�S�?��`?>K?�����򏿉˜�$b2�h7?qnv?E]��/��+j
�����eS�>�_�>`��>`�1��̩>�;:?h������/���:4��1�?��@�5�?��<�2�fY=k�>��>�/<�� ��}2��I�;K�;=?�>���T����_!����A?�`�?�	?� ���0����=�ٕ��Z�?�?|����Dg<T���l��n��G�<�Ϋ=���E"������7���ƾ��
����ῼ̥�>DZ@�U�n*�>�C8�Z6�TϿ(���[о�Sq���?P��>V�Ƚ����?�j��Pu�b�G�3�H�ť���M�>��>�������+�{�Sr;�}=���>��	�>)�S�D'��������5<��>���>��>�0���齾8ř?�b��9?ο媞���?�X?(g�?mn�?�p?9<��v���{�x��-G?��s?Z?�x%��=]��7���j?\���S`�g�4��FE��U>�3?�@�>S�-���|=&>W��>�g>�"/�1�Ŀ۶�'���U��?7��?�o�j��>z��?Xq+?�d��6���[��o�*��O2�h7A?32>����/�!�	/=��͒�K�
?g{0?y�� /�;�`?w�o���]��DT�#�����>��<q>s�>��������K��+�DR�?¿@��?��L��#�\*&?u�>�>�����81�>%%u>���=�>���>Z)>Dܾ��M�:�>���?��?	�?�'����P->�Cx?���>���?n�>�p�>��>��<�=h�[>�鵼�t�=W��>|�B?��?�F>�R@���Z�v g�^�����zN�B��>]�[?�hC?q�=]' �,U>����}����޽����~���hÏ:z�H=�D�>�>�P>t��V���>"?��a�п�=��ڌ��C?��P>�/?mھ�7��ʕ=�f?��n>9�!�쵿K���)����?d"�?^?LW��r5<�4O=��>hY�>K�>c���Q|�
�=*I9?��.�l����i}����>V��?�l@�ʲ?|�]�?H�����&Ƃ��
1����N��=�F:?���>�=��>��6>L���崿jy�		�> �?t��?�.?uR?�`�3,�,s �o=�>�^�?��?>f��gc���>}�>�Y<�o�� q��ܥx?a)@=Y@��b?�롿�pٿn������^�b>�j�=Y>�� �+si��hX<�`�<�[>=O>k��>
U�>J�L>�z>zH>>i>P��݈�t��/����0��7��������p�غ<��]
�����ξ!���/n��*I0�&�Q���6�J�$��O�<(~?���?�l�?���>.�@�1�#?�Ӿ>B�=���>Tր>��>��j?�e_?��?�갽X�Ӿ�e���s���6��[c�>�]�>!T�>���>�>�|��+h>O�->0��>�
_>K`a=���<Ї�=z�>Q��>�*?��>�0<>X>�����A�h�>�z���ν��?�����I��4��QB������y�=��-?��>���7Eп����ڦH?!���s��&+���>��0?��V?̔>z���u�X�g�>V���h��[>�� ���m�6�)�B�P>��?6�f>^�t>vg3�`B8���P�����r�|>_Y6?�Y��	j9��u���H��tݾ�=M>p��>��?��T��薿��~�3~i��0|=��:?�?{U������Fuu�I����kR>�7\>l�=8�=YVM>L�c��ǽ�!H�r�/=�^�=�^>h�?HC)>N��=��>�ܘ�'�U�B�>��N>x�">Ս>?�L"?"A�ur������;�-�`�u>Z��>��>�>�)J��]�=��>��d>����À~�<$�[1>��Z>��y�`0\���p����=�U�����=3��=o3���9��v+=u�|?����t�ٕ�Q��h&;?��?K�T>9Oq=��$�Lۮ��jžu)�?ߏ@Ls�?F?��X��X?橑?a���Nr>��>ur�>�������⸱>�D�*@�)Y��
�@:�?L��?%"K=���+\h��z/>�"?���b��>5��ĥ���Q��s����5��w�>!�S?��ξi���S�
��?���>w����0����ǿ��w�`�>
��?ፑ?��{�J+��
{B���>��?�\?��>#ƾ����/��>rr8?٬&?F�P>�8�A����?�>�?2ч?/FI>/��?_�s?S�>�Xx�]Z/�1������{=��m;���>��>����3\F��ٓ�'{��[�j�����b>��#=�5�>:��Q+���'�=�"��_J��VLf�>t�>ىp>lJ>ߒ�>�� ?�A�>��>�L=����DI��xٖ�z�K?ó�?<���1n�pI�<��=�^�&?'H4?~.[���Ͼը>$�\?P?[?�`�>"���>��迿��"��<��K>�5�>�F�>s��IK>P�Ծ(1D�cq�>Tϗ>��V=ھ�+������#E�>�e!?+��>̮=� ?.�"?�Rh>�y�>��D�5�����E�E�>i-�>3?a�~?� ?�����1�f'���O���	]�C�J>��z?|6?�ʖ>3����ߛ�Hˣ��V�A霽y�?�~c?d���W�?���?�\??]x??ڙd>I�Kܾ�S׽�0�>L�!?���`�A�_6&����kx?�0?���>nٓ�_oֽ�t׼���������?�%\?F&?��ua��þ�5�<H5 ��Y�c��;�
E���>�B>�����o�=��>��=��l��H6��zd<��=a�>���=�7�Y���=,?��G�gڃ�?�=(�r��wD��>ZIL>����^?�n=���{�u��{x��
U�� �?���?0k�?
����h�	$=?�?*	?"�>�I��|޾�ྛRw��~x�3v���>)��>}�l���Ꮴ�<����E����Ž9����V�>���>u!?�?l�>��>	�1���K��������Cj�.� ��0�."����&i��Ᵹ�[�<����%Y��q�>�K��7�>��
?�L>bWY>q�>����?Ġ>O�M>��T>�T�>�v>>��&>�(6>�!�=����H{R?��þ] '�����PU??"c? ��>,�s�������
�`?��?"�?4��>��d�w@+���?�?#�~�Y�
?ř=��;JM�<t���l�2� 
���y���>��ɽx�<��K���b��?`?v�L%˾^н
���S�n=�M�?��(?�)���Q���o�øW�S�ș�i6h�@j��J�$���p��쏿�^��%����(��s*=��*?b�?͌��!���&k��?��df>Q�>=$�>1�>?uI>��	�v�1�f^�M'�T���RR�>~[{?*D�>��J?�A?{hW?�M?H��>�<�>$l��6d�>Y�<p��>z��>�H=?�}/?[�.?�o?�7%?B�O>?c�����dؾ��?��?&"?�	?+d�>7����з���*��Y���d��u��o=��<Vս�Ng�'/=�rK>c[?�����8�����]�j>�v7?�w�>��> �U�����<U�>٬
?2<�>� �B�r��`��f�>���?��=Գ)>���=�����ٺFy�=�R��ę�=}р�r�;�Np <yĿ=�P�=�]x��O*�{��:M�;���<�7?U�?��>rV>�zB��OX�X��b��cf>m��<���>��@��S[���]���=j��?��?��-�#oM>�l���r�Y��"9����()ν�?�d?�@�?<M?���>�?�i�>�+�m탿�^� )��]�?� ,?�n�>���x�ʾ�娿��3���?"u?ZNa����Q)�?�¾�+սb�>�D/�\~�����$	D�fiv���#9��D��?R��?��?���6��q������X���C?� �>x9�>��>��)�
�g�L!�U_;>x��>�R?�"�>��O?6<{?�[?�eT>r�8��/��'ә�{}3���!>v@?Ⰱ?
�?y?�t�>��>R�)�n� X�����g������W=�Z>ؑ�>�'�>G�>V��=i�ǽ�M����>�+_�=ۅb>���>.��>��>L�w>�T�<�F?a�>����@b�gЛ��If���-e?�B�?�H?:"=� ���H��Z��C��>�U�?S�??d)?{��P)�=�0��4���}�����>��>��>ISZ=ֽ�=Lo>Jb�>p��>=Z��a��@��)��t�?�;I?d��=�9ƿ�Cr��r��٘���|<�^��]�d�����Y�-_�=�����U�6���;�Z�냟��7��@`=���y����>�w�=���=���=Zʶ<�μ�O�<-KG=~��<)�=��j�N�j<� 7���ٻ�d��R��m)W<�/L=ΏN�̾/}?�:M?�e.?{�H?�؂>�E->1:��k�>a�N��?�uc> hԼ�Y���E2�`#���O�۾p�پ��b�s����h>��u���>��2>?��=N-�<X��=I�b=~��=\�q���=�ѽ='��=�ȱ=�X�=(�>`+>��u?�.}�i��o����=��ؾf?;�i>�c����I��?q�<���AJ��=��
�u?���?�a�?!N�>
��0��>�F���p'�l�z�i��=��>><!�s�Q���>!�Ƽ+.?��Ф��Q�� i�?�e
@%J-?���I�ѿ��=) K>-�>Z9L��@*�\�M���>�Ά����?*2>�۾��>�h�=g��u�;��?=��H>��=��� ad�_;�=�,��\<�ѻ<��>�;>�ƫ=L�Žd��=��P=wy�=��n>E�t;[O��(�۽�}m<R��=��>	f>��>��?��.?��b?*d�>�d��Ծwþ�>�>�U�=���>Ocr=��4>�{�>�6?\_D?��L?���>X5Y=V��>iܦ>�Y,��o���d��Y3J<1t�?3R�?ʿ�>N٩<d6��<�X�=�H�ս�?*W/?!A?�>���1Nӿ����J2��D>�w�>�.�������<�[(>�P�=�O>��">�Z�>~��>�V>>�͒���=֊>[�>>�*>�� �/@>�����н��l<�Q��Л�%#0>,�c<����Ҍ=9x�>	��!�=��=YK�=�6�<0��=)��>u�>,��>��=-����'.>� ����O�_�=����E$>�x�c��y��01��/�Y�R>y�k> M��~���)��>��e>�kG>lS�?gLu?��2>�7�?L�Gǟ��LH��C�΁z=�> ��:9��:^���H���Ǿ��>��>p&�>��i>��*��?���V=�߾5�3��&�>,����8��Z�c�o�k*��*.���ok��F�#�F?����ʰ�=�}?cG?��?g��>�����վwi)>#����$=k'���f�kU��<R?�P(?F��>��̭E�	Q˾2´<�>�I��P��ȕ��0�5���ֶ�7ʰ>`%���dϾ�2��[�����a�B�s�s����>�P?)̮?�d�o퀿kO�H���E��7�?�yg?&�>�V?`\?/���<�����L�=��n?r��?�N�?�}>�Ƚ=�=���D�>�F	?+��?ṑ?�}s?uF@�W��>��V;�!>n�����=y�
>(�=�\�=�}?3�
?�
?�]��n�	���\��]����<,��=n�>�;�>a)r>6I�=3�g=���=��[>���>�Џ>p�d>��>�C�>�T��{���&?��=�Ӎ>042?�~�>Y=:��@��<jJ�	S?�}k+�zq��pPὂV�<�@�Q=�̼��>ˉǿ�3�?��S>��?�@���1���S>d�T>z޽���>�YE>&}>o|�>��>�G>�z�>L,(>�Ӊ�V�{>1�4�X>���s�>�o�9�	��{>o���ח�p����~�<�n�1�������c�������L� ی;P{�?�\���%���M���?R�k>��Q?�rZ�k���3H�>��5?�l�=����͕��Ғ��վ�n�?n @��>6��>��8?�o2?]H5�(N+��MQ�t&��QE���o�� p��瞿(Qr�n޾���<?nj?�?�B,?B�[CX>Ja?�U�(\����=2:}�>(i�A���X�>�ⴾ4��=uJ�����mfh��g>�8?v�\?���>��
�vB��v�>�Y�?*|v?r�?uUD??r�?P$����?���>�$*?�5?n�s?q(/?z��>��=��Q�H�,��1	�Y?ٽ�,���ޕ�p,��vL�>J�v>��C��)>ػ�<����&�ʼ+\�;��<4�ٽU���^�=i���
�f�=_��>��T?S�N>���>Ar+?J�=��F�#T:���e>튿��z���凾
^�sH�<����C?>�?�~~?�s���FJ��� �f>N(�>�$�>��:>)x ?�K�eO�����U>��>5���������޾<8Y��wQ>?��>�?�.�<����X3>��������$>�Y�=��4��kҾ�u���*��b2;� �?#�W?��/?�z=��ž_ w>baF�z6&?U�Y?�J?`P|?=�����?��Nc_�&�(�Si�>T�E�,�A�⭿7v��o��,K>G�>\.��uז�d֐>�Q ���]�t�X^�<�ﾽ��<���<M�=14��־\48��t>d��=mĹ�WI!����������X?썎=I.���gJ����<�/>ZZz>Ǐ�>}U1�b���@0�|"e�i�=��>��!>*\�B��XAB�'$�@�>�PE?�S_?�i�?����s���B�����Rh���gȼ,�?�j�>�b?�B>��=j���(�b�d��G���>��>��h�G��<��G$��_�$����>�4?�>b�?D�R?��
?n�`?�*?�B?�"�>���
���B&?懃?A�=o�Խe�T�2�8�9$F����> x)? �B����>��?V�?0�&?4�Q?��?�>�� ��I@�В�>\�>�W�Ca��?`>��J?���>�5Y?0Ӄ?��=>Z5�آ�~ʩ�>�=�>��2?3#?z�?R��>O��>󬡾+�=��>�c?�0�?��o?�w�=��?�22>a��>o��=���>��>?�WO?Q�s?��J?���>q��<c8��h3��*Ms�[�O���;wH<C�y=���:t�c7����<���;-m��4�����D��7��;%��>�gm>�h��X31>��ľO틾�d=>G$\�/���Ǎ�-E�!��=%��>��?H��>��vҏ=��>gn�>dZ��>(?.?��?���;�c�u޾WP��>@?��=�^m������jv��D=9m?��^?�V�����R�Z?XZ?/�;�0����|l��r����A?�'�>��z��>%��?�jl?���>�"���Ń�����6y�ƅ߽�.����>)]���Mb�/\�>��?-��>��x>j��<��ܾ��b���m���?�ɉ?H��?TK�?��T>��w����N���K��)^?0��>�?��& #?����-�Ͼ3P��f(��⾙��A���B���x��}�$�ރ��׽��=y�?js?�[q?a�_?̳ ��d��1^�*
��=kV��(�&�7�E��'E�őC�b�n��b�0��#����G=��~�͐A�R��?��'?E�/�؛�>����I��'3;��B>$����J�#�=u㋽(T@=�_[=B8h�TU.��4��
 ?e-�>Y3�>��<?�[�">�ٞ1���7������3>��>���>�N�>�G�:�e-����rɾ�����ӽ\�u>8�c?y�K?�9n?3&��A1�E ��l$!���4�s��@�A>��>�d�>��U�Oc���&�*�>�7hs������cf	�>-�=.�2?X4�>q�>�K�?(�?�#	�I�����z�t�1�j�<�L�>�i?���>��>�ͽ�!��F�>�LT?���>��|>Y���_!�5up�L���`�>k��>O3?��y>����A�y���n����X�:t]=!��?�����.E>��8? *>�E���7>��-�, $�ړ��'���>�>�X?:�/=Q8>U᭾�A!�R���z�P)?�J?�撾�*�,3~>�#"?~�>�.�>�/�?�'�>�rþ�JM��?��^?BBJ?�TA?9K�>,�=���O<Ƚf�&���,=���>U�Z>�"m=/u�=?��Sr\��w���D=�y�=�μ�Q��*�<���zK<��<��3>�Iο
1��[��]��̾�&�Z���Z�1�?z%�["�<�®���x�A��U#�ߗؽ9�=�0rS��g����Y�8J�?�@��!?��'����Ĕ��
�q�>���Z�-�%�k�Ɗ����þw����d�G��\����x��'?W�����ǿk���Ձܾ��? ?�y?B���"�8��!>^��<����>�������ο������^?��>`�5�����>�|�>|�X>�Hq>l��Ӟ��!�<�?J�-?�L�>'s���ɿ·���r�<���?5�@�WA?�4(�f�]Z]=�K�>?�	?4|?>��3�$��4��N��>���?�x�?*�B=��W�����e?--<��F�m���=<��=��=�����K>���>�T�P�C����,�6>�$�>�^,��E��\��<��\>�ӽ���	��?n]���d���0��u���>��U?o��>?��=e)?��J��ο�-[��wb?3��?�'�?C&?�<�� `�>.>۾��K?��5?�ݝ>��$��|u����=pܺ�
�N�S��A�U��s�=|��>�f'>�O-��J�u_U�{Mx�d9�=6 ���ÿ�h,��	���V=�T`�_q.��n*�7���f<3���k�ϒ��oz=*��=a8M>`��>�T>�e>�l\?tz?X��>���=rh��ޱ��Nʾ�민6�]���	���w�z�������/�۾���.}�������ͭ4��w>}h�����=%���|���C�� ?�OE>;���8�R�7�.�6g���P���{5�7���.;'u;�vFt�Q_�?��W?�S����M��l3����`�ҲM?S}齒�������->��=���=�W�>x�`=���T�?�6�W��0?),?l���ZB��K)>� ��C=n+?W�?w y<���>~%?�r+�����Y>��1>���>��>~h
>��-�ڽGQ?�T?��w���#|�>ڷ����{���g=c�>YG4�?�[]>k�<O0����{������E�<a�T?(m�>������H��%r���p =w�[?џ?�;?{�o?z*?#%��-�о��^�<�@���Q�ҸU?��z?���={}�9�߾�܋��b?̟2?�o>�>��� ��i��R�S�?��`?>K?�����򏿉˜�$b2�h7?qnv?E]��/��+j
�����eS�>�_�>`��>`�1��̩>�;:?h������/���:4��1�?��@�5�?��<�2�fY=k�>��>�/<�� ��}2��I�;K�;=?�>���T����_!����A?�`�?�	?� ���0����=�ٕ��Z�?�?|����Dg<T���l��n��G�<�Ϋ=���E"������7���ƾ��
����ῼ̥�>DZ@�U�n*�>�C8�Z6�TϿ(���[о�Sq���?P��>V�Ƚ����?�j��Pu�b�G�3�H�ť���M�>��>�������+�{�Sr;�}=���>��	�>)�S�D'��������5<��>���>��>�0���齾8ř?�b��9?ο媞���?�X?(g�?mn�?�p?9<��v���{�x��-G?��s?Z?�x%��=]��7���j?\���S`�g�4��FE��U>�3?�@�>S�-���|=&>W��>�g>�"/�1�Ŀ۶�'���U��?7��?�o�j��>z��?Xq+?�d��6���[��o�*��O2�h7A?32>����/�!�	/=��͒�K�
?g{0?y�� /�;�`?w�o���]��DT�#�����>��<q>s�>��������K��+�DR�?¿@��?��L��#�\*&?u�>�>�����81�>%%u>���=�>���>Z)>Dܾ��M�:�>���?��?	�?�'����P->�Cx?���>���?n�>�p�>��>��<�=h�[>�鵼�t�=W��>|�B?��?�F>�R@���Z�v g�^�����zN�B��>]�[?�hC?q�=]' �,U>����}����޽����~���hÏ:z�H=�D�>�>�P>t��V���>"?��a�п�=��ڌ��C?��P>�/?mھ�7��ʕ=�f?��n>9�!�쵿K���)����?d"�?^?LW��r5<�4O=��>hY�>K�>c���Q|�
�=*I9?��.�l����i}����>V��?�l@�ʲ?|�]�?H�����&Ƃ��
1����N��=�F:?���>�=��>��6>L���崿jy�		�> �?t��?�.?uR?�`�3,�,s �o=�>�^�?��?>f��gc���>}�>�Y<�o�� q��ܥx?a)@=Y@��b?�롿�pٿn������^�b>�j�=Y>�� �+si��hX<�`�<�[>=O>k��>
U�>J�L>�z>zH>>i>P��݈�t��/����0��7��������p�غ<��]
�����ξ!���/n��*I0�&�Q���6�J�$��O�<(~?���?�l�?���>.�@�1�#?�Ӿ>B�=���>Tր>��>��j?�e_?��?�갽X�Ӿ�e���s���6��[c�>�]�>!T�>���>�>�|��+h>O�->0��>�
_>K`a=���<Ї�=z�>Q��>�*?��>�0<>X>�����A�h�>�z���ν��?�����I��4��QB������y�=��-?��>���7Eп����ڦH?!���s��&+���>��0?��V?̔>z���u�X�g�>V���h��[>�� ���m�6�)�B�P>��?6�f>^�t>vg3�`B8���P�����r�|>_Y6?�Y��	j9��u���H��tݾ�=M>p��>��?��T��薿��~�3~i��0|=��:?�?{U������Fuu�I����kR>�7\>l�=8�=YVM>L�c��ǽ�!H�r�/=�^�=�^>h�?HC)>N��=��>�ܘ�'�U�B�>��N>x�">Ս>?�L"?"A�ur������;�-�`�u>Z��>��>�>�)J��]�=��>��d>����À~�<$�[1>��Z>��y�`0\���p����=�U�����=3��=o3���9��v+=u�|?����t�ٕ�Q��h&;?��?K�T>9Oq=��$�Lۮ��jžu)�?ߏ@Ls�?F?��X��X?橑?a���Nr>��>ur�>�������⸱>�D�*@�)Y��
�@:�?L��?%"K=���+\h��z/>�"?���b��>5��ĥ���Q��s����5��w�>!�S?��ξi���S�
��?���>w����0����ǿ��w�`�>
��?ፑ?��{�J+��
{B���>��?�\?��>#ƾ����/��>rr8?٬&?F�P>�8�A����?�>�?2ч?/FI>/��?_�s?S�>�Xx�]Z/�1������{=��m;���>��>����3\F��ٓ�'{��[�j�����b>��#=�5�>:��Q+���'�=�"��_J��VLf�>t�>ىp>lJ>ߒ�>�� ?�A�>��>�L=����DI��xٖ�z�K?ó�?<���1n�pI�<��=�^�&?'H4?~.[���Ͼը>$�\?P?[?�`�>"���>��迿��"��<��K>�5�>�F�>s��IK>P�Ծ(1D�cq�>Tϗ>��V=ھ�+������#E�>�e!?+��>̮=� ?.�"?�Rh>�y�>��D�5�����E�E�>i-�>3?a�~?� ?�����1�f'���O���	]�C�J>��z?|6?�ʖ>3����ߛ�Hˣ��V�A霽y�?�~c?d���W�?���?�\??]x??ڙd>I�Kܾ�S׽�0�>L�!?���`�A�_6&����kx?�0?���>nٓ�_oֽ�t׼���������?�%\?F&?��ua��þ�5�<H5 ��Y�c��;�
E���>�B>�����o�=��>��=��l��H6��zd<��=a�>���=�7�Y���=,?��G�gڃ�?�=(�r��wD��>ZIL>����^?�n=���{�u��{x��
U�� �?���?0k�?
����h�	$=?�?*	?"�>�I��|޾�ྛRw��~x�3v���>)��>}�l���Ꮴ�<����E����Ž9����V�>���>u!?�?l�>��>	�1���K��������Cj�.� ��0�."����&i��Ᵹ�[�<����%Y��q�>�K��7�>��
?�L>bWY>q�>����?Ġ>O�M>��T>�T�>�v>>��&>�(6>�!�=����H{R?��þ] '�����PU??"c? ��>,�s�������
�`?��?"�?4��>��d�w@+���?�?#�~�Y�
?ř=��;JM�<t���l�2� 
���y���>��ɽx�<��K���b��?`?v�L%˾^н
���S�n=�M�?��(?�)���Q���o�øW�S�ș�i6h�@j��J�$���p��쏿�^��%����(��s*=��*?b�?͌��!���&k��?��df>Q�>=$�>1�>?uI>��	�v�1�f^�M'�T���RR�>~[{?*D�>��J?�A?{hW?�M?H��>�<�>$l��6d�>Y�<p��>z��>�H=?�}/?[�.?�o?�7%?B�O>?c�����dؾ��?��?&"?�	?+d�>7����з���*��Y���d��u��o=��<Vս�Ng�'/=�rK>c[?�����8�����]�j>�v7?�w�>��> �U�����<U�>٬
?2<�>� �B�r��`��f�>���?��=Գ)>���=�����ٺFy�=�R��ę�=}р�r�;�Np <yĿ=�P�=�]x��O*�{��:M�;���<�7?U�?��>rV>�zB��OX�X��b��cf>m��<���>��@��S[���]���=j��?��?��-�#oM>�l���r�Y��"9����()ν�?�d?�@�?<M?���>�?�i�>�+�m탿�^� )��]�?� ,?�n�>���x�ʾ�娿��3���?"u?ZNa����Q)�?�¾�+սb�>�D/�\~�����$	D�fiv���#9��D��?R��?��?���6��q������X���C?� �>x9�>��>��)�
�g�L!�U_;>x��>�R?�"�>��O?6<{?�[?�eT>r�8��/��'ә�{}3���!>v@?Ⰱ?
�?y?�t�>��>R�)�n� X�����g������W=�Z>ؑ�>�'�>G�>V��=i�ǽ�M����>�+_�=ۅb>���>.��>��>L�w>�T�<�F?a�>����@b�gЛ��If���-e?�B�?�H?:"=� ���H��Z��C��>�U�?S�??d)?{��P)�=�0��4���}�����>��>��>ISZ=ֽ�=Lo>Jb�>p��>=Z��a��@��)��t�?�;I?d��=�9ƿ�Cr��r��٘���|<�^��]�d�����Y�-_�=�����U�6���;�Z�냟��7��@`=���y����>�w�=���=���=Zʶ<�μ�O�<-KG=~��<)�=��j�N�j<� 7���ٻ�d��R��m)W<�/L=ΏN�̾/}?�:M?�e.?{�H?�؂>�E->1:��k�>a�N��?�uc> hԼ�Y���E2�`#���O�۾p�پ��b�s����h>��u���>��2>?��=N-�<X��=I�b=~��=\�q���=�ѽ='��=�ȱ=�X�=(�>`+>��u?�.}�i��o����=��ؾf?;�i>�c����I��?q�<���AJ��=��
�u?���?�a�?!N�>
��0��>�F���p'�l�z�i��=��>><!�s�Q���>!�Ƽ+.?��Ф��Q�� i�?�e
@%J-?���I�ѿ��=) K>-�>Z9L��@*�\�M���>�Ά����?*2>�۾��>�h�=g��u�;��?=��H>��=��� ad�_;�=�,��\<�ѻ<��>�;>�ƫ=L�Žd��=��P=wy�=��n>E�t;[O��(�۽�}m<R��=��>	f>��>��?��.?��b?*d�>�d��Ծwþ�>�>�U�=���>Ocr=��4>�{�>�6?\_D?��L?���>X5Y=V��>iܦ>�Y,��o���d��Y3J<1t�?3R�?ʿ�>N٩<d6��<�X�=�H�ս�?*W/?!A?�>���1Nӿ����J2��D>�w�>�.�������<�[(>�P�=�O>��">�Z�>~��>�V>>�͒���=֊>[�>>�*>�� �/@>�����н��l<�Q��Л�%#0>,�c<����Ҍ=9x�>	��!�=��=YK�=�6�<0��=)��>u�>,��>��=-����'.>� ����O�_�=����E$>�x�c��y��01��/�Y�R>y�k> M��~���)��>��e>�kG>lS�?gLu?��2>�7�?L�Gǟ��LH��C�΁z=�> ��:9��:^���H���Ǿ��>��>p&�>��i>��*��?���V=�߾5�3��&�>,����8��Z�c�o�k*��*.���ok��F�#�F?����ʰ�=�}?cG?��?g��>�����վwi)>#����$=k'���f�kU��<R?�P(?F��>��̭E�	Q˾2´<�>�I��P��ȕ��0�5���ֶ�7ʰ>`%���dϾ�2��[�����a�B�s�s����>�P?)̮?�d�o퀿kO�H���E��7�?�yg?&�>�V?`\?/���<�����L�=��n?r��?�N�?�}>�Ƚ=�=���D�>�F	?+��?ṑ?�}s?uF@�W��>��V;�!>n�����=y�
>(�=�\�=�}?3�
?�
?�]��n�	���\��]����<,��=n�>�;�>a)r>6I�=3�g=���=��[>���>�Џ>p�d>��>�C�>�T��{���&?��=�Ӎ>042?�~�>Y=:��@��<jJ�	S?�}k+�zq��pPὂV�<�@�Q=�̼��>ˉǿ�3�?��S>��?�@���1���S>d�T>z޽���>�YE>&}>o|�>��>�G>�z�>L,(>�Ӊ�V�{>1�4�X>���s�>�o�9�	��{>o���ח�p����~�<�n�1�������c�������L� ی;P{�?�\���%���M���?R�k>��Q?�rZ�k���3H�>��5?�l�=����͕��Ғ��վ�n�?n @��>6��>��8?�o2?]H5�(N+��MQ�t&��QE���o�� p��瞿(Qr�n޾���<?nj?�?�B,?B�[CX>Ja?�U�(\����=2:}�>(i�A���X�>�ⴾ4��=uJ�����mfh��g>�8?v�\?���>��
�vB��v�>�Y�?*|v?r�?uUD??r�?P$����?���>�$*?�5?n�s?q(/?z��>��=��Q�H�,��1	�Y?ٽ�,���ޕ�p,��vL�>J�v>��C��)>ػ�<����&�ʼ+\�;��<4�ٽU���^�=i���
�f�=_��>��T?S�N>���>Ar+?J�=��F�#T:���e>튿��z���凾
^�sH�<����C?>�?�~~?�s���FJ��� �f>N(�>�$�>��:>)x ?�K�eO�����U>��>5���������޾<8Y��wQ>?��>�?�.�<����X3>��������$>�Y�=��4��kҾ�u���*��b2;� �?#�W?��/?�z=��ž_ w>baF�z6&?U�Y?�J?`P|?=�����?��Nc_�&�(�Si�>T�E�,�A�⭿7v��o��,K>G�>\.��2݈���>�N �
T���v����i��!�Ik�=���WU̾&��$槾�~Ӿ��=u�>�*
�|@&�g����S��U�l?󽬽��̾�	��-^߾Oɀ>�=n>��?�'��s�>������쾫4)>V�>\�>�t���-����D�_���q�>x9?��i?yw�?l)���ZU� �R�}���:<���J�J0?�J�>9�>��>MZ6<(�þ}��D(Z��4�8x�>:N�>ކ3��28�)հ�6��� O
�r}>H/�>.�I>�4	?�	P?� ?�8I?�0#?Hr?�2>ف=b�����&?�F}?0e<�%���+��!�"�+� �>ݪ(?#��h��>*�?T�%?>R8?bc]?K%?��=���!wB�C�x>Y��>�S�`����>�W?���>��6?�d�?=�> qL�x�Ⱦ4����5
>�%>�e5?��?gl?Ȗ�>��>p����=�A�>@g?���?��m?���= +�>jT>r�>�V>Q�>-��>P�?}�N?Րy?�tF?ذ ??}�<o��p	��u���
ݼ���z�!��)�=�E���V���{ü�Y$=�����4��2��Bh��f�O��㾼0v�<w�>��v>c��b�2>:ľ�\����@>����a㜾*`����6�+u�=}�>Ɗ?�?�>	�"�@2�=��>�M�>'���(?!�?>?-��;�a��VھI�N�l��>_�B?w��=��l��w����t��dT=�gn?�^?��S�=���'�f?mGQ?~����K��3��nKn�˻վ}i^?��?3���u�>SӀ?�v?�f?���
:�G���]���v�J!�=�K�>�b+��w��U�>�<?��>��e>|gx>Q�ھ�s���_���O?���?ǩ�?_?�?<�=b�o��6տQpﾬ����d?��>q����&?YcǼ�Ǿ���zFW������ͩ�q𵾕G��2����K��̃��,н�t�=�r?O�d?}n?��Z?j� {b��h��탿etQ�!J��L�;u0��G�t�?�WPk����������	�=��n���8�褵?4�"?��8�|�>u�� ۾��ƾ��>+����
 ��<S�̇%�5���a���$�j���*$"?#�>{��>�a5?�c^��=��B��E���׸>0@�>Ь>�j�>� �ۖK�-��6"� �����"��>�B]?�L?kB?-N�r�;�hT����'����q���R�>��>��S>e��clC���(�S�,��v>�&]��#��J-�uW�>��G?
�{=�Z
?�ڄ?�^?�(��p쾩n,�ՀD�6�S��?��O?
U�>p�?�&,�k����><�n?;��>�&�>���X'���~�] ��{�>B�>�%�>A��>���&\_�7Í�$
����9��	�==�a?��x�|��ҍ>�"P?Ge	��n=Kv�>ke7��z%�����o���>���>)�=�%[>�߽������s��X���-K?E$�>����z��� ?�*}?��-?��!?���?���=bo������rA?��y?!bs?C�u?���>.9�=��[>{�8���k�;�٘>9�>��=�r�<B�7��T���-� ��=+�=�&��rs���~��=0��o�>��=���><ѿ^9��uҾQ����6��Q"�n몾�WG����g�!���ؾ������@�<T1�CP��Y��+�Z����w�(9�?�W�?-�"��(�N��{���g�
�J��>U�b9��T�����r꨾��	��5E��*#���=��Jl�����r�'?Ӻ��Žǿ򰡿�:ܾ?! ?B ?�y?m�˞"��8��� >UV�<T.��М�[�����ο����v�^??��>k��,�����>饂>�X>�Fq>����瞾�7�<U�?%�-?���>}�r��ɿi���kդ<���?�@�\A?�$(�;��p�^=�=�>Y2	?-8?>/&0���X	��C�>c9�?��?pGO=j�V�K��be?�P <�G�M����=a�=ɕ=��t_J>3�>.��4-B�G�ݽ�_5>v�>���+��<�]���<��Y>�[׽������?�[�j�f���0��J~��>��T?l��>j��=O�+?oZH���ο��[�߇`?���?���?�5)?.Ǿ����>+ܾ�EM?p�5?c�>��&�.�u���=�|�CS���㾗�T��"�=���>�>��,�����
N��綼���=�� ��/ƿI5(��W�e=�kcb��l*�Ր(�q� =/E���{��.ǽ9�=�۸=6T>p'�>w:b>�Y�>��W?��r?�Y�>n_R>���i)����Ҿ-���q*^�EE�����n�"��v}���
��(⾣�������� ʾ#�:���=��L������D'��,m��I�w� ?��2>�վ��H�t��<��վ�����]�<G<��ʾn\1��r�+��?(�D?�F����K����v���ɽr�T?�Y��"��i��T��=����R�G=��>��=��F{+�{�L���=?=�?�M �OX����>Uʇ�7��=I=?�s�>�I���>�R<?����!�W��>z��=�B? ��>�w4>�y� _x=�,?���?ǎƾVV�����=�z���3%�s9�S"�>�R�<0��=�q>���=�W�����+�=�#о�(W?l��>��)�S��`�����z[==̲x?��?�-�>�zk?��B?ޤ<{g����S�2�bw=��W?*i?e�>c����	о)����5?��e?��N>�bh�����.�YU��$?��n?�^?�x��w}�U��]���n6?��v?s^�xs�����L�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?}�;<��U��=�;?l\�> �O��>ƾ�z������0�q=�"�>���ev����R,�f�8?ݠ�?���>���������=w_����?Ҝ�?೾�͏<�g�L�o��n���=���=a�м��ɽ4���A�~�Ҿ�&���f�f��>�&@���L��>F&8��P俴�Ϳ��Cf׾��R�)�&?�N�>�
����n�9�j��L���A��t����> 	>�K������z���/�H���r�?�JK�(�>��S���<���t��$�=�t>���>ou>��V�9	���Ƙ?|U۾�nڿt����]žbV+?f�?�s?;??���2�Ҿk�����= �e?�ӌ?wK}?��S����5Yܽ�j?`��gT`�L�4�IE��U>"3??A�>�-�ɿ|=�>��>wg>?$/�N�Ŀ�ٶ�������?L��?�p꾾��>���?2t+?!i��7��;\����*�h!+�B<A?@2>x���ȹ!�/=��Ӓ�л
?�~0?]w��-��_?.a��q�|.�xŽ���>D\/��aY�$ܼ�7!��je�s���]u����?�P�?t.�?����#�6�$?��>�s����Ǿ�5�<�6�>7��>�9P>Æ_�A&w>����@;�R�>��?r9�?&�?wo�������> �}?���>o�? ��=��?���=VN���A绵�>�����1$�um?RsV?�?��>� ?�9�UN2�4�5�����PF��4�>��g?^k:?n<*>�K�t�⼛�.���p�y�,��G|K��6ռ��`<��>���>ZZ�<�r��1���?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�c��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?bQo���i�B>��?"������L��f?�
@u@a�^?*��ٿj5����޾��b���>	�<x�>*����<�>�H�=&!X=�%>1>���=yXh>��{>�bH>%��><����[!�ì�>[m��&��������O��PS޾K������3r����"ؽ� �uP������8�콽���=�MV?��M?�8o?���>�f�� >�����C <��E��ɶ=���>u&3?�tO?��.?Av�=>����\�a��'����Tz�l �>��2>���>���>|@�>�m���s>%�\>��]>���=
|�;���<�'ƺp�}>���>
�>�*�>��>õ�<j�����,}�6 \�w�����?*��LOF�E�y�k*��P�T�Ks�>�"9? �]=����Kοwbƿ/(J?�y�	m��Ҿ�?�>�I?�֑?ݬ��&*Ǿ��W>�u,>zs�J�#��X>Mi̾]�>���e>, �>�Ճ>�7>��4��L>��T�c���m�>��)?�<׾x�UBs��)a���ɾ��>�+�>r�|=�h4������u�4�^��r=<=?��?�a��伾ῆ��C����>�o�>"Ğ�ܪ�=scm>�p�>d�!W����.=p|>�S>i�?��+>X,�=p�>☾2|F�I˦>�JE>��">�>?�X#?M������v��1���i>���>jV�>|��=�bK����=�p�>�+^>}_�Ҝ{��P�ԗ9�6�V>���GZ�Vs��:|= �����=Q;�=
��nD� �%=��~?XিF�����5���%|E??
�=���<�u"����꺾aA�?��@[��?~��f�U��2?5�?�͛��e�=�>NR�>��ɾ��D��?�Vý�����f�V�!��ˮ?� �?�.������Gk�2�>�&?�vϾPh�>{x��Z�������u�x�#=R��>�8H?�V����O�e>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9�~�'���?�޶?֯�?�x�>�?�_?_#�>�=�y�z���.����Q>��>.�>)p>�<|�|�l��8��=p����k���ھ�)I>�:=���>�૾�����)>B�Ͻ��L�Y��]u?"}�;��&m�>xf;?]��>�o�>���<��}<+��*3����N?��?����:|�Rx=�0�=u?.���?��B?�V�����>kl?���?%�e??��>�*�@����繿NC�����;.�>�Q�>�A�>��<$�>�qξ?l��t�>ȧx>uF�Ež�]���i<1(�>n&'?%��>b��=T�?��? "�>xξ>УB�댿#jM�N��>��>\�?KG�?O�?�y��8U1��.���+��[�O��F>�xq? �!?# �>'x��Hu���sa��7ͽ�Y����x?��e?i��� �?6҆?)b:?c�C?h&�>�󚽑�޾$U1��sv>\�2?���4<O�֑Q��|��Z?b�>?dX�>߾A�v�t<�=��l��ͫ�w ?��?�jW?h�9��w��������<����o;��)^�=79���&>f>�3���6�=;�>x�7�Q<ľס��=x��/M�=��>!(Y�����z�>�B,?5�;��1���E�=�er��RD�Cm>��L>Jt��J^?�;��2{�Ѭ�>L��S�}��?d��?�j�?P���.�h��&=?�$�?�T?Һ�>�b���a޾�?�p�y�(@y���=�>ڃ�>~PV��f����X��������˽�@��P�>m�? 3?"�>md�>�)�>�]��P!�;|>�b����K�r��y5��@A��&#��������彏߾d�����>ȧ߽���>ݏ?�*>��>�^�>J�$�@b�>@N=e^b>a9R>�i>��4>��<>ӷ��"�𽘮R?~���4�(�z)��䬾��C?�'e??��>�>5�58�������?K��?��? -�>��d�Q�)�Rl?$J�>��}��s?�3=����]��<������Y���p���9�>�)Խ�2<���L��b�s?�+?��mƾ�I���Um����<���?��9?%g,��dE��)z��m��Z���>��#�!�m�K�#��r����������#�S�=�c)?��?����=���fAl�Uy���K�O�O=1�>�y�>�i!?c�s>r,�ns���X����T��i��>g�r?��U>d�_?p<=?}�G?R|j?Y��>/��><���&��>H�<�#>���>�/%?�n;?P�1?@?J�4?"��>�X���B����?��?j�?B�>#�?,�����<Ń�����e�~L�<f��=(��<P�-�ڔ����ʥ0>�X?���٫8������k>��7?��>J��>���*+�����<�>��
?�E�>� ��}r��b��V�>9��?����=��)>N��=�����Ӻ�R�=|���n�=/6���w;�mq<׀�=���=!Qt�GR����:	W�;�t�<3d�>�?��>9O�>H?���� �������=��X>�.S>�>^Fپ�u��I!����g��!y>�p�?ap�?�rf=y@�=�q�=�����T�������-7�<~�?�C#?�NT?ю�?Y�=?5]#?y�>��nB��9\��[
����?)8?�`u=\�߾�\��d���?P�>��W���=�$\�3����=>�9�B��R�Y�L���[R��8��,��A��:���?Dޠ?d�`�:�N�>�z������^�1?�yO>+�#?��>��1vr�ӱj����>��F?lv1?��>� P?��z?~�Z?`aR>�M8�"ﭿ6(���g9��Y>yX@?Ć�?ޔ�?(�v?�~�>��>w)��߾�V��������)d����W=#^U>W��>0��>��>���=O�ǽ2ҩ�u%<����=�@c><N�>��>�}�>piw>蟿<+�H??��>Jjþ��E���u��[��v?2:�?A�(?B�<F��XB�˳�,�>k�?�L�?Y)?�;H���='�̼K���4�f��[�>aa�>J�>?v�=�&-=/>���>�N�>�����1p7�F�a�!W?��E?���=njſ��q��p�(>����]<T���`��f��[�U��=�����o�髾�]b�0s��©��v#��P���#�r�,��>V�=��=K��=~�<<:˼��i<-U=�ׯ< =eT��+<j�=�=T��l����3��i9;�%+=�߉����Ԯj?��b?��,?�q&?c��>��a<�=V�]>�$=� �%?a�,>�P�������Z{���Ҿso#��+�S,Ӿ��S�R�����=	;���=��)>�J�=bv�=���=���;�T�=�V�<"n�=43�<���=��=��X=w��=ޘ@>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��B����4�?��@��??�ዿТϿ6a/>��7>4>H�R��s1���\��b�G[Z��!?fS;��j̾>X�>��=@߾5fƾ�1/=Va6>w�a=����a\�/͙=ьz�=�;=��k=,̉>�D>l��=����9�=p�I=���=��O>�P��ٕ7�>�,�/Q5=	��=V�b>=)&>V5�>�-?B�$?��Z?���>܉'�ž��˾�2�>��=C�>���=��	>*7�>�r2?�:C?�H?=�>`�=�>���>b ���e�����7Q����E<4�u?S͇?���>X�f�@q��')���1�1�G�X?��B?��.?*��>y\���!�:��K����=bw!�
y�=3��*5�=�#��~��<v��=�с�p��>.�)>4D�>���>�_�=��>.�>��>Th�=8w�<J-� <ԥ��&;J#4=Ö́=�C��#�ڽ�l�=���<����������@S==���<f�={�>�Q>2��>aې=P'����.>������L����=/4����A�G�c���}�dE/��9�*C>~QX>з������?�Z>��?>!U�?8\u?
q">6�؁վ띿��c�ٳU�a�=V�>�`<�>d:���^��%M�^[Ҿ;��>�5>���>���>��G�'�#�b�:%$��#&�w
?o�ܾN}�r�+�h�o�����n���,�]��q�<��)?����U��=�P}?~�Y?o�?t\?�z7=�1��f�>�,����<����:��Q��=(��>��?�?+8��L�!���˾)R���z�>�G���O�������0����������>����nо��2�IO������$B��3q����>&�O?�?Wb�v���Q.O�����=����?�.g?���>+l?� ?餟��,������=�n?oL�?�4�?|6>�,���=_�?)��>���?w�?As?V	a�xc�>hT<�=�`�=�}b>K9v>Ź�=�X>w4?��?�"?*����%�;H�������}�}��;?@�<h{q>�r�=17�>�@�=_>�i0;�&~=�<�>�ח>�J=>8�>_B�>����t���)?'�=2Օ>�S2?ѿ�>�*4=���z�=�r��A���谽z�ག�%=���<��C=O��#��>��ƿM��?md6>���	�?.�������&>u>Ž���>�@!>[Ld>���>ަ�>B:>��~>��*>�GӾƗ>����T!��/C���R���Ѿ�hz>����)&�Z���R���cI��o��k[��	j�5+��F:=�w��<MH�?ш���k���)�*���v�?�R�>g6?�܌�A���[�>d��>鲍>�9��ᇕ�`č��k�u�?���?:c>6�>T�W?{�?#�1��3��sZ�	�u�x%A�he�S�`�4ߍ�������
� ��P�_?�x?<{A?YA�<�1z>^��?v�%�Aԏ�q2�>	/�%;��G<=c.�>���'�`��Ӿl�þ�7�B9F>�o?	&�?n^?c<V�{���n�>��;?�t?Y�?�7?��K?t�8�Y}.?�H>GG�>�9?4?q�??��?�A>���>:�>% >Z��<<���#余�@�([0�"=�d�=R�ʼD�(=a��<DD�<KvZ=��=�H�-7���Ά=�t�=7B�����=�_�>\(q?bn�>΃�>pMZ?��^�hE�jӠ�1[ ?�">�r�;�Y���Ǿ�n�@>ՁQ?�:�?��?䔧>C���'ٽ��>v\�>u4�>��>K��>��<{�$�u��=�ph=��N=��=_�?��]0�����c?�Ƹ�=���>�j�>|>/r����!>�Z�� nu�ۢe>�IK���,aV�M�G�@0�ÿv���>�5L?�R?��=4��+ʊ���e�� )?�<?��N?�~}?쮀=@ݾ{�9��L������>y��<���|j��p1����;�Hr8;v%u>6���mz�*>����Bz�p耿��T�����r^>�Q9��0>$3�������+ͽF,*=޲D>ů��-!��ƙ��?��=to?u�����ľ��n�!����h>#�>��>#�N��m��N�0����4�<A��>�`\>]�=����w�e���5��ք>�M?�[??�?kI[��q�
�<�����d	��1
2���?p|�>!�>4h8>�q	=w�ؾ��*]���E��z�>	r�><����J��ാ�>���"�>�~	?fW7>�?�X?\�	?��g?N! ?�?_:w>�-������,)?L�?��
='@��]E���.�ss:�u�?�+?��_�>��?�?w�6?��T?)�?6� >����A����>��^> �Y�fǮ� �t>��R?���>g�_?h��?�:�=uA�\-��z�{�d9>I�v>��A?A?��?�*�>��>���O�=��>Yc?21�?�o?���=&�?j22>)��>���=%��>��>�?�YO?��s?��J?j��>!��<v*��J5���7s��mO�5m�;�H<��y=B��9t��4����<�}�;bf���J��.�񼿯D���U��;���>��t>ꯕ�o�1>��¾����4j@>����<����@���T;���=w!~>��?�>�!��d�=J�>hR�>b��ZR(?�*?�~?�;wCb�>�پu$J�8��>^ B?�;�=?|l��U����u��*\=?l?��^?&_W����s�Z?�o?P0Ѿ��K�19��t�����ն!?�?@�c�K(�>�J�?
�}?.B�>>���X�}R����8�OՆ�s=�=/�q>{)��yM�
s�=y�*?���>T��>��>͔��`d�oӌ�}w?a�?	��?ȉ?��$>P�r�n�e?��"$���V^?��>�d���:#?El�=�ϾRf��kS����⾥Ӫ��⬾�㕾�t��[%�	{���(Խ@�=^?��r?Kq?D�_?Wf ���c���]����V��m����uoE���D�1C���n����fn��齃��bF=��z��B���?��.?e�@�3?�0���������ݨ%>M���T���̨�V��~���y9;
����\����k�>�1?�>#�>�(>?�9R�\J_���Q�cW�"�ݾ���>�_�>���>�,�>me=_������; ����%�t'���w>�d?*�J?J�l?����a{1�µ���f!���$�ځ���}F>�E>JK�>esU�g���C%��=�H�q�]���v����	�Z�v=\03?�ky>���>%4�?8�?t�	��e��j�v���0���_<�L�>U�h?�.�>
�>Y�ս{�!�޸�>��l?���>{	�>Ht��D`!�{�{� �ʽ��>�ҭ>���>�o>M�,�k#\��i��>����9����=��h?-�����`�vͅ>OR?��:�&H<e~�>�Vv�Q�!�����'��>�}?�Ϫ=|�;>�zž���{��@��`=?�&�>ap
��LH�{:�>v�\?�
?^��>���?�	�����9�=W�#?�t?�$~?<��?��>����W�=ɕ�%wq�J�ļ
��>��>rz�<�l��ׂ����x��<�$>� >2��h���CR������
�=k��P:
>:�ѿs3A���ž�Ѿ�?�z}�3���Q[=�ž�ࢻ��z�?������X�S�)9K� ���+z��]R�r=�e��?z��?�Y��h���Z���8���q��?)�;lTo�CyǾǤ���GU��z��n�]�s����X�������w���(?0痾E�Ŀ����ྤ� ?�o$?�t?*���<�4�:�~$�=�+U=Q벼i��M��?�ο�ݣ�x�Z?�U�>Y=��ҁ���>(l>E&A>ZmS>�r���⓾���<�?I�0? ��>2����ȿtU��$����?�@�xA?7�(����(V=}��>*z	?�?>X1�TA�����d�>�:�?���?��M=K�W���	�}e?.Y<� G�J�����=CO�={4=���~J>b�>;_�uyA��ܽ��4>���>2H#�i��9�^�Ͻ<B�]>��ս�6��1Մ?�w\�Af��/�Q���p>�T?t,�>h�=��,?�7H�VyϿb�\��,a?�/�?���?Q�(?R῾8ۚ>�ܾՋM?D6?���>a]&�N�t��W�=�9��}��S���V��=��>�w>��,���}O�7C��%��=ǳ������%#�).���t��>�Ǎ�}[ѽ�)߽�)W=3UN�9qF��F�KA���=k^�=η�>�5�>��>��X? �a?�4�>g>Y>��@�~؝��׾�9>�k������$����N��������ћӾ���I&����ښ���<�^�=��Q��揿;!���b���F��_/?d�>�eɾ�/M�f<��Ⱦ^���PUw�����.g̾��1���m���?rQA?^օ�Y~V�	���.�Θ��LsW?[�p���խ�P��=[;���\=�w�>g�=�7���3�NT��s2?r�4?�ɾj�N�\�>�ͪ�g�Z�r�!?���>�d�=��>,�K?� ���ۺb3�>N�o>�B�>�t�>�D<�b��c��818?�|W?DNp��u¾�_[>]ʾ<���\�`>�$(>A���ν�A�=7�Pi־�J^>�ܔ�	|"��(W?o��>��)�C��`��2���b==[�x?��?u+�>ezk?��B?��<`e����S��Pbw=�W?�)i?Ϲ>ő��1
о�����5?�e?X�N>;ch����p�.�TV�#$?��n?!^?rs��v}����
��-o6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>��������>�F��*��?��?�`�M���1��房�0;�\�=\ A>���=��>�������k���ʾe�������>D��>�l@Tn���Ĵ>�|a=#�����ֿ�����Jw��xt�\l?�8�>��=d\��a��P��F/��[*��kk���>p_m>cc�]�F�o��'�P�M�&�?�}�	4>>�-9�p�z�����,�_>f�j>I�>�s�>�T�7��<ܙ?�c ���ſ凲������q?Ɯ?�e�?0cW?��p�SѴ��5&�bx�=�q�?�z?e{�?S�I����g��S�i?Y����W���/�I��8U>�1?P��>{*��ަ=08>��>��'>��2��ÿ����w��4y�?Ӳ�?G��@�>U�?��-?�]�2���|ɯ��<)��d�9p�>?J�'>l騾�&��<�����%S?�.0?Pn۽�~��d?�3���n��|8��~ ����>�D;7�>ѷ�>��˾9�[��-~����;]�?���?y��?y�۽U�'��y?��>ȯ����i3�~�>sb�>�S�>-JȽ�0�>�&��o�U��=��?���?�?
�R��$���c>.��?7��>wJ�?���=�6�>1�=-ꢾpL��#H>��=���v�>�\Z?� �>,H�=:n!�s�+��6�G�N��h��G��y�>~�c?��B?f�3>T����k�e%��]����#�q�����,�E�����q>�>�G�=z�8��<ž��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*�hֿ����jN��R���%��=���=͆2>:�ٽ2_�=�7=`�8�=�����=h�>��d>�q>Z(O>�a;>�)>���I�!�r��Q���P�C�������Z�B��Xv�Fz��3�������?���3ý,y���Q��1&�@?`�="�==V?4�Q?�|o?a ?��r��>����HP�< M"�#ل=lF�>��1?��K?�f*?䴐=y���T�d�r���)���І���>xH>H>�>.��>;�>��R�d<G>!?>�w�>'�>�*)=�YJ�Cj=`�K>i��>�]�>Xi�>��j>{*g�௨��m��y�����C����P�?�վ�UG�m �������׾b�>7!?�+5>T5��P�ؿ?���LfC?Ƌ��;x������P>>#4?!̀?�O�<7Qj����A!>�n��T��w�>Á^���'�����wI>� ?}��>��&>F=.�#>�AQ�%d��GǮ>�-?�&ƾ����+s�_��L���WN>z3�>�;i=H�����`�|��:X��v=�	4?s�?]\-�t���g�c��U�����>n(�>�=k:H��=:��>ag����ɽ3�D� �N���>���>��?�M8>�<�=�*�>쇖�vcK�Lئ>
>>�z >
�>?��#?�����A��������'�#�q>�s�>+1{>�K>�U�B�=2�>�.^>�g-�Ts���+���I��N>Q6j���Z���e���}=ꟽ���=4�~="��� :��,0=ė~?jw���房g%�����yD?o1?Fl�=��M<ۏ"�m����2��0�?��@�q�?�^	���V�ĸ?�=�?������=�o�>zԫ>�;D�L�t�?�)ƽ�͢�Ն	��#��K�?.��?�N0�TË��l�77>\T%?��ӾPh�>{x��Z�������u�x�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?:��>C�?3�n?E�>j_�>��Z���ȿj���W>�I"�9� ?#*�>Z����j�<��y5x��yO��3y����>��<Ҙ�>��������>5�g��k��,�=�Ð>��(>P}�<Bw�>7�?���>�b�>��
=�b�=�aP���¾t�H?c�?��
��)i�j=���92�@��>�0?��
��ݔ�cC�>Rd?�Ix?ee?��><��}~��)~ÿ]a���Z���K>!�?|ۘ>���� ~�>zF�������jT>�J�>�TM�L^��H��E�҉>u7?Q�>��w<�~?~�%?�΋>^Y�>x�5��|���N�$�>�g�>@�?kǃ?�-?5�����3�����$C���-R��&l>�v?8�?�4�>^��s]��#=1� Ͻ�:�?�!f?Z1�}b?\��?JnA?g�4?p�>����ھy����i{>�N*?پ����<�3D�GN��ܝ?	;:?$F�>˶�7�ܽ�3�;�R�Ӄ��VT	?(�;?��=?!� ������n���o=�%=-��<L=�I>NUX>�46>80�͸+>�ɮ>@�<�䊾[�?=�୼��=O\�>�Ľ��ֽ�	D>�<,?|�G�sڃ�k�=�r�uxD���>�HL>�����^?Aj=��{����Ax���	U�' �?��? k�?���~�h�[$=?��?�	?�"�>J���|޾3��bQw�&{x��w�,�>��>W�l��徖���阪�WF����Ž�t\�Ah?c�?T�=?��>>T>ǝ�>��*��'�g�l��E�I��-*���P������8�����M�*<����d������S_">lѥ��^�>��>!�'>�Vu>J5�>X!O����>�3
=��=>���=�J=��>�;�R�Z�	bR?����(�)�{ޯ�n�B?�bd?xn�>��^�ȑ��b��z?*s�?A~�?
�x>�g�l�*���?]d�>���@�
?��<=����`�<=���g���-������̎>�{ս/�9�M�"g��*
?B�?bǇ�Nd̾Ytֽ����]�k=[��?<t)?X�)�IQ���o�N0X�oxR����i�f�Q��<%��Lp�.���.�����mt'��4=�*?�3�?���7��K���Ml�n�?�Ttb>K&�>k+�>Z��>K>9��T�1��^�#�&��V��U�>��z?��>�#N?�y7?I�L?$2H?Q��>yd�>>$���4�>>���>���>�4?��*?@�.?�?_�-?�#U>q�����p�Ҿ�A?\�?ς?��>R��>���� �Aau:�脼邾}���,O=(%}��(��?��e=i�]>	Y?�����8�����mk>��7?��>^��>����,����<��>K�
?G�>�  �P}r�(c�U�>k��?���[�=��)>g��=Y����Ӻ5X�=a���r�=�0��.|;�/s<ꄿ={��=�lt�$���@�:WՇ;�~�<'b�>�? ��>��>W��U� �o��8�=!�X>��R>4\>�3پ����[��}�g�<hx>���?~c�?�ie=t��=��=o���,x��
�kٽ�t �<x�??P#?ST?���?��=?�d#?nE> �L%���W����E�?`2?|]�=C���;ľ�=��p�@U"?���>��G����07�����>\��<C�1��;_� ���f"���=���U��m��?rJ�?�/$���<�����J����`��3?�!�>i�?���>�yE��Gl��TC�BU�<(PZ?o�c?�`�>��V?��q?r(I? 9{>2�;�z#��R���C�6<	U�==�C?���?���?"p?���>U�>�i)�`�ξШ�P@3�!��YC���.�=�t>�>�l�>���>r<�=;(��ⰽ@�8�#�=	߅>���> 
�>P��>+�P>�m-�$�G?
��>g������ߤ�z����<�C�u?C��?'�+?o�=5{�S�E�;-���]�>�q�?c��?R**?A�S�:��=�׼�ᶾ��q�B%�>�ڹ>01�>���=e�F=�T>"��>��>�'�d�l8�=M�k�?F?�û=ڦƿ�'q��~�`Q���K<������^�Ă�� �O���=U��h��Uݫ�{�Z��)��!��')�����9�^��}�>���=?>�X�=�V<r�����<_|=5<�	=��\��R\<)_����H��ɻWo�-�e=�3�;<�ɾ�*~?Q�H?8,?�QC?�w>�>�=����>N���`~?XbY>�`�+	���y;�y����y��ckؾ��׾-�f�?F��n2	>�DM�*K>�03>���=J`<�=��s=Ƌ�=`u%�s�=lg�=ű=�={��=��>Q�>�6w?X�������4Q��Z罥�:?�8�>l{�=��ƾp@?~�>>�2������wb��-?���?�T�?<�?Eti��d�>M���㎽�q�=@����=2>z��=u�2�V��>��J>���K��5����4�?��@��??�ዿϢϿ:a/>�p8>�&>8�R���1���^�)�a�=�W�L�!?�x;�&R̾���>��=�d߾�	ƾ�S,=�+7>[�a=���F�\�3:�=4Py��<=lh=�͊>��D>�d�=�����=�P=~��=X�L>yVN�m9���,��6=rC�=g�b>�U'>�>P�?�;0?�%e?���>�&p�
�ξe�����>�g�=��>���=ˡ<>��>�}6?�[B?��L?�t�>ق�=���>Ѷ�>�,���m����*צ�揵<���?���?GK�>;ـ<ye<����y<���Ž��?60?�1?xx�>�
�����sA�,N7�H��;��^�ln�<N{�ˈ�=�r�>Y�=L��9R*����>�>���=z	??��>��]>T��>��=��=��=�����=�2����<(���=���=��l=K&3�G剾& \<�J���@�5>�j�= ��=���>>��>Y;?EK9=�k��  <>�Q���FH��>6����A1���f���v�!!�+fv��=,>��Y>絏�iɛ�d?�G`>�I^>qA�?�W^?��d>�T�ž�W����y�鉺�f��<\=qK���6�Na0��kC�_/��B��>�^�=��>�M�>��>��`��v�=w#��� �x�?�ӾQ�%=����V��)����������a>��R?�ᗿ��>mY|?<�I?��?)�>T�����}m�=��N����$�>?۾L���"?P�?xJ?K���(:��G̾��^߷>�9I��O�p���0�l���ͷ���>���4�о%3�4g������ҎB��Er�y�>�O?Y�?�:b��W��oUO�.���'��bq?�|g?�>K? A?���bx�o���t�=��n?ٲ�?�<�?�>=��=劳�[C�>�T	?G��?���?Q\s?�?��3�>e͂;�� >ژ����=��>S��=R�=)�?�u
?4�
?P���w�	�����H�^���<���=/��>���>��r><��=��i=ⶢ=j�\>+��>7E�>˂d>���>���>� �����w:?�?>��>�lO?��>�i=G����$��
k/�����1@��-"����.����̝=�ր="��>�ʿ��?�R<>w����?xd�߽yD>V;'>�z7����>���=Ȼ>��a>�ә>�Xs> 8�>*F>BӾxw>e���d!��,C�S�R���ѾQ{z>����]&���ב���6I��m���f��j��.��;==��ν<�F�??����k���)�M���~�?�U�>�6?x֌�x���>���>aɍ>^N�������ȍ��kᾀ�?���?�;c>��>�W?қ?�1��3��uZ�ܮu�o(A��e�f�`�J፿1�����
�,����_?��x?�xA?C�<,:z>�?��%��ӏ��(�>S/��&;�D<=�+�>)��k�`�@�Ӿ�þ�5��GF>��o?�$�?$Y?{QV���m�7 '>��:?��1?�Ot?��1?H�;?ˡ���$?jo3>uF?�q? N5?��.?!�
?2>�
�=U����'=�7���@�ѽ�~ʽ���@�3=�]{=ݽѸ��
<F�=���<ǘ�ټ��;!(���!�<�:=��=S�=�>o�]?=c�>8i�>��7?���K8�SӮ�k.?��2=0���|��������>z�h?'�?��Y?W�`>��B�ZMB�v�>�t�>�X&>8i\>z��>̦ｗtD����=�>ug>�=�JN��v����	�m3����<��>ޥ?&2�>Tx	��4>��%d>���%>E�̽3����ܓ�#�P�־��l�>I�P?l�?��R>���7��po�I$?�ML?8Y?�W?n�u���ǾG)�z�i�ò%=A��>�w)��T����������X� \e> Fi>���%阾�]d>Bt��׾aur�s�K�gE�{�=�S�� �=*��bھ!r�z��=��$>F_��md��������XO?��<f!��{t����H�9>��>�>�3R��ᇽ�9>�@2�����=iR�>R�$>��!<:��I�#D��ʉ>�]:?�Th?y�?<S���i��{E����T��+)����#?3j}>��
?G��=az=��о4��i�L�W�>����>���>���P��䟾����Z��MZ�>��>J�W>�~?�^?�a�>��]?@�,?!/
?��>��½L���:�(?LM�?��==�����J��l5�ro?��L ?��-?��e����>�9?�?3�)?��R?��?Km�=C
��:�*o�>�O�>S�]����� i>�	N?{�>I�R?�?�Q1>�N=��Қ��wp���=��E>c7?�*?{�?=��>�#�>������=�\�>	}d?�v�?�t?M��=Js�>��(>4 �>X�=�+�>��>�2?�I?2�s?g�P?���>pu<�yԽ�୽�%e���������0;��=�L�&���o��܃=ž���J�gě�`Dx�t������JJ�<*E�>�by>���� �2>E,ľv��3?>}	��$n��0z��(�8��ٹ=TRy>ό?ڟ�>�J$�v�=u��>J��>���l(?�?3�?��-<�6`�(�ھWN����>)�A?�\�=�l������v�k^=X�m?�`?�LJ����#f?%nQ?����f=�*竾+�o��;˾Y�b?\?	�����s>�E�?�:p?��?A#��Y3�؃��J-y��~H����=��>��3���q�	ǰ>�E?�*�>܉b>kV~>�e�Kp���f���?Φ�?�Ʒ?%+�?�=;[��B�ȿ8��5���0b?+�>/ ��-�#?El����Ѿ������x���g���xi�����;ۤ�t ,��/��Ϝ�����=Go?�Vl?��r?ڋb?�� �h�	�c�C7��'lQ�M���p0>��hF�<�>���q�M���C������/��=O,m�UE�"e�?�g-?12n���>2w��q�꾇YǾ΋z>����ؔ��p��<u�ɽ���<b�7<V�V����R����,?w�>.�>�JB?��Y��II���B��uG����?,>���>t;�>M�>�I�;��]�R�"��ܾ1�_����k��>o??�3?��K?��6�G�Q������!��8Խ�C־Cȋ>�n>D�	>�#W�����x�*�KO��Q�D�������,����=fR>?L��<I�>�"�?_�?|C���ܾٿ���Q�.�ٽq*�>��O?�v�>�@K>oн2�8����>��b?h0�>&^�>Ƚ2�F�����@��~�>_�>da?�>O8���c��і�2C��cY.�9�(>RIc?j�K��z��ES>1�-?Ǜ�{�<�?�>��O���"�E��'�t����=���>5_>�I>r1����xUq�>���ɷ@?���>J��aY�k�p>��2?�!?@��>3ڞ?�I�>��7��Ӎ��[?棟?cit?��q?���>��q�Vl���<� 9��61"�%h> �>>;A0>5ɐ=�~H�,mƽ{�w=4�l=0��kR�����= �=/�ݽ��=��G>�	L>4yҿq�6��xվX�;Ҿ��$�ܘ�Ƽ���e�bh��{���ς� 2��x�O�(o�p��/�Qˢ���}�� �?�u�?]ܾb�������aҀ�P*�LD�>�����=&��^��J���� ��¾3%J��4��@*��-K�sN�[�'?����˽ǿᰡ�j;ܾ#! ?B ?%�y?����"�ƒ8��� >�H�<~,��Y�뾁����ο������^?^��>��U-�����>q��>��X>�Fq>-��X螾�9�<�?��-?��>��r� �ɿb���⽤<���?$�@�|A?O�(�/�쾠�U=���>	?'�?>R31��J�����^�>2�?��?b5M=l�W��	��re?�|�;�F�axܻ�=�Q�=qk=A��(�J>Tf�>yt�iA�l�ܽo�4>���>�"���{�^����<wi]>n�ս0|���e�?�2K��l��4���m���D>��U?Pd�>�F>�]-?��Q��6˿�HE��z?���?�m�?"�?)O��/ը>5�۾F=U?��.?�̘>Q���p�� �<�kX�A�u�����u?�#�#>���>��0=̦������R�;C���>�7���Ŀ��� �<8�<�"�˗6�����p��;�m��Ȕk�)۝�>��<r�=��j>���>�G=>�]N>}L[?
r?O�>��)>c;��B��7Pྥ���w��o�:��t�@j�9���\�-���Y=�����p�8���=X��儿4��[ml�R�H���0?��=��ɾK�6�& ;=������!<N1�⏶��A,�5�c�|M�?�A?p�c�E�Ր����s���b�q?��9��nؾ�:��	�=��y<83<w��>�T�=ށ;||�>�J��(?3_+?ŋ��||�b� >%��|鿼��+?T��> ;�!��>e�3?��s�v�P�ӡ�>��>�Z�>�_�>
q <f��곪�9�B?y�R?��|��s�W�>x����׾��
=�t>x�����I�8Q�>�n�;��`B�<�g��Ut�}(W?���>��)����`�����P==�x?ʒ?�-�>^{k?��B?rۤ<fh����S����`w=��W?�)i?��>����i	о����޿5?��e?D�N>�ah����X�.�PU�\$?��n?<_?\y���v}�w�����Vn6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?s�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>��������
>ɯ�4�?��?,.Ѿj�D;d�!�-�w��-��>E�=§\=�3.��(���=�3-۾ɋ�IXo�5�<�5�>��@/��2��>T��b@꿧�ɿ�����þ��W�M�C?���>T*9�������[Pt���b��?��⠽I��>E�3>���2�P��qz�N"I�㐊�p�I?�be����>�H�������j��0~��w�>?��>n�>�^���Vپ�9�?,���Qu���u����ԾdZ?y��?Dm�?�?s)�E�Ӿ�����>|fN?�I?f��?�^N���h��"�j?�_��YU`�͎4��HE��U>�"3?�B�>S�-�ô|=�>���>Cg>�#/�l�Ŀ�ٶ�}���H��?Չ�?�o���>o��?�s+?yi�8���[����*�A�+��<A?�2>����S�!�E0=��Ғ���
?V~0?�z�Z.�˸_?I�a�	�p�p�-��ƽ�ۡ>8�0�%T\�������Ze� ��@-y����?E]�?�?��N#��4%?~�>�����;Ǿ��<�}�>�,�>�2N>q_���u>��g�:��^	>e��?}�?cj?�������tY>c�}?nֵ>�:�?�V�=%��>Sy�=I����̉���*>���=uI��Vt�>�,P?U�>�b�=�0��.�c?�J�M�ul���E���>��f?��J?/�F>kُ������� �Y��Kc#�%|ɼ�y=��W�K鹽o:>��">k/>��K�0{Ҿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Ra~����7�U��=��7?�0�'�z>���>��=�nv�ݻ��R�s����>�B�?�{�?��>%�l?��o�P�B�X�1=0M�>Μk?�s?'Mo���o�B>��?"������L��f?
�
@~u@^�^?) �޿B2���[ľu$����=R�=�4$>���)��<rn;����U��<��5>:l>	�.>oWk>�c>3P>�Z0>�v������噿G�v�E�LO�D(�~�d�J��gb�vV�þD>��Y��o��&�������#��HĽE��=]?��K?aN]?/^�>ZX=�>d�Ҿ-����;z���<N�>P�?�CQ?]�7?��3�A�]��2T�톃�CƾD�9��)�>��J>G�>�t�>�%�>יl��r>u�z>��>���<�.P�2�b�ٮo=�9X>6��>�>W�>9�n>4E�=�浿n����+g��$V��u�X��?�຾��L����u��ު����=C�?�S>Ea{��6Ͽ-��
[D?�Jþ�s�v[�nI>��D?�]?y��=����$�gF>PJ/�ӿP�R&>����L���!���=�m?x�>�q�=��3��B���[���W�kR�>�9?�=�\$ ��Bd�Fx~��΢��p >؉�>n�=0�0�<���|���R��sI<��S?�F	?9���ξ�6n�θ��SȐ>1��>3�+��R�=��>Q�J�ӪF;�r���A7���=A�>�!?Q2+>i�=1��>����O�i�>A>;V*>O@?Ö$?�K������̃�Γ.�=�u>r3�>�ɀ>`�>�L�є�=�P�>ra>4��߁�3��Ѿ>�,W>��z���^���u���y=}A����=u��=�v���+<��&=�~?�c���舿X>뾉����pD?3?sv�=�W<_d"�����P�����?��@dt�?�I	��V���?�:�?(`��q��=.f�>	ϫ>��;\�L��z?ZƽFբ�E�	���"�%P�?��?-[3�|�����k��.>AN%?ҙӾPh�>zx��Z�������u�o�#=Q��>�8H?�V����O�e>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?toi>�g۾=`Z����>һ@?�R?�>�9�}�'���?�޶?֯�?�3r>{7�?w�^?� ?O�>��Z�����D����}�>��u=��>��{>`���[�N;��N���L�d�¾E �>�fe=��>ա����s�=��{�$���r�ܽP��>��>��Ź_�>�O�>�><>�ă=�D=U�������M?�Y�?�[�1cp�C��<���=��J�l�?+�9?�+��6ݾ�ѯ>��_?qƁ?c�]?	>�>�{��|��ḻ��Q����< v5>� �>�&�>��:�k�X>�پ��:�G�>�>����̾��o��;�ٚ>E!?@�>8�=T�?g�?���>	�>؄�(㖿}�b����=�3�> `�>]̟?��?����r�A�m^��Y ��6�_���>�È?6G?�|�>=c���ؙ�R�>�Ӓ��[��!z?�e?Uň�t�>63�?&U?��'?�o�>w�����J�H���&=P)0?�fj�lxd��F�9�>��
?��(?.U?�⽈s�{���G0�j�p�t�?�;?�P?��ݾ�s������'=���>�n=t�޺ڲD�k��>á�>^�V��7�=�ǚ>��ټk�׾�����=�J>L�c>Tq�U4��g�#=,?�G�dۃ���=e�r�xD�u�>�IL>���^?Rl=���{�����x���U�� �?���?[k�?���E�h��$=?�?N	?k"�>�J���}޾+���Pw�~x��w�:�>���>�l���D���љ���F��(�Ž/��Ϯ�>W�?D�D?���>
]>�n>�����K3���پ	�ؾH�}�6V��L�0��@�5*�)�ԾU�����]�}1��Žbv�>hj,=AMk>݌?bi$>v��>�A�>�=�Q}>GrI=���> �<
B#>�ͦ=�3$>Jo >�*=�LR?q�����'���ߪ���3B?)qd?�3�>DSh��������z?�?Tv�?w]v>srh�*+��g?b@�>����s
?�L:=5�*U�<~U�����H���-�|��>%׽:�$M��f�\g
?�-?�	��w�̾�1׽��l���<���?2LG?*|/�ªK�"4v�f��G����=�|���U���q:���n������ԇ�����K>��!?�J�?�5� 2�p�Q��р�4r0�;>�!�>Kg>R�?qR>���;f-�,�Q���#�����Y�>���?�uv>O�X?�A?#�H?��W?�9�>w�>�G����>a}=�G͚>c��># *?&�*?53?Ǣ?�a5?��>�&�<��;�׾%�?%�?I2?l�>i�
?�����e��O¼�Ƹ�~�X��E0�7N�=n2	<ם��d���᜼Fe)>oX?K��`�8�����/k>]�7?ǀ�>���>���7-��� �<a�>�
?�F�> ��}r��b�^W�>ˢ�?Q���=��)>@��=�����ӺpX�=~���?�=�4���s;��n<��=��=�4t�I�/��:p��;�t�<�t�>�?&��>�D�>�@��� �u���e�=�Y>�S>8>xFپ�}���$��{�g�}\y>�w�?�z�?e�f=�=���=�|���U�����R���d��<�?J#?;XT?X��?��=??j#?|�>�*�HM���^�������?R�3?"}=k�	����ѳ�"��˨?�\�>��T���M=A�/�	���#=(��=�X��~N�S����M�1q5����8��X��?͛�?��g�6��w:�Ǥ���T����R?��>~k?���>(��Hs��t:��>�"?��N?�0�>�'O?u�x?�b[?A(e><��m��(����c<^(>>@?�?�?T�?br?�K�>b>�&�.ھD"�v��~>��NV��*�)=��Q>\ɒ>p'�>6A�>ܼ�=��ͽN�Ƚ�2<�L�=�h>l^�>��>T��>]g>�A<�bG?��>����������ۏ��U�>�k�t?.�?:{*?j=/����F�{*���7�>M��?<�?��*?)DS����=B�̼R�����q��>���>���>���=�S=m�>j��>�O�>yC����R�8���D��y?Z�F?��=�3ƿJ�q��p����G<�ޒ�6�c��򖽠�Y��֧=�ɘ����Eh���\�������8���H6���|��~�>?�=�p�=�Q�=�$�<��ż.S�<�O=�W�<8=x]m�T,z<�b>�#���f���b�7b^<��C=����3�ɾVu?�[H?�+?"�7?�2�>3`+>��t��r�>KX��+?&�?>�y����žʃN��٢������@Ծ!⾨{�$��JI
>b���]>'0:>t��=�p5=y4�=9��=u��=g�<@�<���=ׅ�={�={>2>�+>�5w?���������8Q���罫�:?EV�>��=כƾ�@?^�>>!9�������^��?���?5I�?J�?�i�"_�>l��m��t�=���F2>�5�=[�2���>^K>����J��F3���*�?ӄ@�??�苿5�Ͽ�h/>��H>?��=X��5�x}k��P�љ=���(?��?���پ:��>��e=E'޾�|þ���<#�R>c��=ԇB��a��t�= �½�TK=�<N= \�>��f>1�=�V߽!d�=���<{�>[�0>�=�;���K�v���=�
�=BtO>Q�>u(�>3(?2*?�"Z?���>�ۤ���ƾql��H�n>S�4��b�>R��=/6�;�{�>+(H?Sd,?�Fe?s��>J�.=2�>���>�$&��AU�&�p��Z���=��c?U�?���>��:=Up�.�*��mU����?�,O?.:?��>H��Yۿ���[PJ��ܟ����o�="cn���<�P>�#���<x
�=�.�=��>���>�ˆ>�Jg=�.�=u�>���=�|�<��=��ؽƓ�Y��<��">�`�=�N}=��ɽ-�6<B7/=���<�O="4�<7락�EI�@$�=���=���>��=>9��>1�v<&���8�6>�䭾��N�W�>ꍳ�}j8���\�ܦr��q+��R����=��4>����4���2?�M>]�/>u�?ZVq?GWZ>�z����Ⱦ�t��1U�
Y����>I��=��0��*���A��B�?+侴��>�!�=j}�>^�>��0��� �ﲻ����B�\��>��m���Q�Hf5��#X��(���x����s�"wG�;�
?`ǐ���'>�m?V0V?�#�?�?�dU��Z����=u9��Å ��| ��\T�e�����>���><?h签p5A�U�Ⱦ�`����>�?/�'�N�씿�1��0������!ۭ>����qVԾuC1��O���z���"D��n��>��K?pt�?^�T���O����	K��s?�i?���>�	?�?�+��(2뾘�w��o�=uTn?c�?@��?�X>=^� Ғ>�3?^��>2��?y �?�#�?�����ˬ>SD��A=�0�=���Q>��*>���=��K?'�A? �3?�rR�Z�9��ӾT־wU��~����RB>�i>��=���>Ws�=]��=q�=�m�=چ�=�s!>�/�='�n>K7g=̵���O�[�.?..>��>f:?�>�U=$b��S\�>}#!��M��]�C���gк:�����6�=j|��F��>ECƿ~��?g�K>�Y���?�����4�_:�>�>q҉� ?������>��>nr\>�8�>�l�>jނ>�EӾf~>v���b!�,C�c�R�ҿѾ�}z>`���/&�<���~���EI�an���g�qj��-���;=����<�G�?����b�k���)�����s�?�Z�>(6?�ڌ������>T��>]ɍ>{K��D����Ǎ�/fᾊ�?%��?��b>��>d�W?��?'�0�X~0��6Z��Wu�h�@�%e��5`�]����ʁ��"
�VX���]_?�ey?t�A?Q{�<c�x>���?E�%����f�>�~.���:��w7=A�>�G��q `���Ӿ+ľ���e�D>�o?J�?9)?��R�x)����2>�;?��*?r�x?c2?M�@?(��*W!?AD9>�:?Ɍ?>&/?��-?2 	?�3+>Y�>O�<z�F=�w��p���Gxֽ��vW�� =�<|=;I��)%�{N=���<v���L���Q�;�Sּ4�<�7=ê�=�*�=�m`>g+�?��?!|�>7Q?l�&>|g�����n�+?�`��xX(��$e� o���ξh��>i�B?ž?٨�?\��>�����^���>� 0>�0�>�i+>� �>������Q=�a�=췝=͢n>�3��#~����ľ�v���o� u�>�v
?N�>=�w�)�<~K��ֽ'�<>������ɽ�����&?������m)�$-?�|d?5�2?���=�ܾBmһ sh��(?�@?͗T?�IN?�w�K+��m�.�|�_�;�/�>�r>�2�MG��T旿�<D��8�=b0�>ͥ�v�Y4*>�V۾��ν������R�>��� ?��L�>�M�.��*�q=O��=�*�>

�����D���F��Wfn?� ��=x�<ԉ�6���q>�w�>�h�>-<\��3�=�3�2#��wU�=��>Tn>�������-R�B���Ƈ>��D?�b?i��?D6U��xM�]L����z����<��?/ne>���>��=q�L=@����*�J�&K@���>���>��(�ǖI��f��IX�-� ��z>.a?s�L>�?�YZ?��>�\i?��'?o?���>��4�ž�.?x?�Y��\|�𽐽7�&���$���?��??އ��q�D>o�?�x?3?��i?[?��=c8���R��Mk>��>��w��'���({>�EB?	b�>�L:?���?�Ȟ>�\J�y�����c>;ҟ>��>��J?�6�>���>[�>i��>����(��=��>�c?%1�?��o?�s�=�?#C2>���>D �=e��>n��>�?2XO?��s?��J?}��> ��<�:��/���=s���O�@�;2H<�y=ɖ�m2t��I���<��;�d��/@�����^�D��쐼x�;+�>%�s>����0>�nž5���EZM>�z��ǘ��.u���tJ�s�=��>j��>K�>�	&�η`=
��>:b�>t��lr(?��?��?q�<��_��Qվ4�	ڬ>�=?���=�Gm�@꓿i*t� 	�=Wm?p�[?�O������ba?��\?�.�:��|��a�����J?�D?Z�G��2�>	�?�k?��>�_�~]i�]�����[��Uh�~�=n�>���a���><8?<��>��f>;ɘ=�\�k�x������?���?[v�?)�?T�>�es�V_�`�󾩆���{d?���>�ϰ��"'?��v���ܾſ���J���T��w��[<���E���뗾�qE��M�������=��?]�e?y's?��_?ia���g��+b��}���K�b��$�w�>�H*K�N�B�	�w�	��j��_⎾
��=�}���6��'�?E�-?֕T�v?S���K��buǾ4��='Ƭ��㽁L�=��y�=���p�g�n��ޡ�"�$?�ؒ>/��>��<?��a�ڔ?��:���I��	ؾ~E}>��>��>�a�>���4y�h�н0ʾ�m�}ۏ��*�>�*U?S29?�	Q?��E�\�I��:��ú��v)=.3Ѿp��>#�K>o�'>*3�4ս'���*+�U]��U��>c�M���W>�0?�b
>12�>��?�8?��I�dd��r�����S���-��>�|T?��?귛>���OJ��Z�>>�i??'�>���>yBL��S=�X����$��r�>���>�'?�4�>veG��JL�W���`ሿ�*,��JG>�a?XY��퀾�xk>PI?; �%s<s6�>@=1��#&�js���>n��^�=��
?�	�=K�&>�񆾙���ǁ�(h��6e-?VR?���b#L�TU�>X?��?Nrν;d�?�5,?o���s8�M��>y�?��m?[X?4$?M3�<�j¾�w�Aϼ�w
>�+�>bm>=�>�J�<�/V�Q���e��\!�=�#E>|d=��A�z��c����>5#D>�">��ֿ�$��qѾo���Ͼ^���ʟ�n޽Ng���l/�����b���i�wun��F��A6���ٽ��R�zL����?���?�α��؁�ݮ��І���ݴ?��}����i�8԰�ھN:���h޽:����k�^�^��S��q+?�g��
⽿��Mо+L+?��;?X�h?�	�Տ)��\=��cP=WF�=��d���В�(��������o?^;�>R7ܾ!Ge<?o�>�j%>̽>Y�p>����J����={� ?*�6?G?O���;��,���R���q�?�@�wA?�(�I��n�T=D��>�I	?G?>rn1�	����b�>+�?�?;�M=D�W�(
�Te?d<��F�3�ֻ�C�=1��={=��I�J>"Z�>�\���A��0ݽh4>g|�>ް!�����_^��6�<�	]>��ֽ^p���ӄ?�d\��f�y�/�>M����><�T?4�>��=�,?�:H��vϿC�\�p=a?1�?f��?m�(?�⿾��>��ܾ<�M?:6?���>�c&�ϲt����=�1�6�����@V�I��=I��>-{>4�,����>O�cɘ����=�����ɿd�1������>��<���½�q��N��﫾/ƽDpO�ב6�H�<�h>���>3=>!D>>uN?&$j?Ҷ�>J��=WY��Mg��î�n�缐���Z�Q��怾�~�� �����!�Ѿ]r����`���ľUN?�v�=@"M�e8��G�R�e��OG���0?�0>�{о��C�!{��b�ľ���l����!������!�+�d9n�K:�?��<?#����H��f�S�!� ׽�d?L$�,������ԡ=W�h��z=�L�>n�=����0��K��\0?}�?�U���q����,>����!�<b>)?+6 ?:�<1e�>г$?v�3���ؽ�6]>�9>���>(1�>�t�=��Z��r�?OU?o��P��3��>����S��n�n=>u�B��$�-Z>"�<&���Nƺh���Nԑ<vW?���>g�)����BA��0� ��<=0�x?�?Z(�>��k?�B?���</H��G�S�'��0w=��W?~ i?��>7�о�q���5?��e?��N>�Xh�)�龒�.�>e��?��n?mV?����P}�@������K6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>���������=*��� ��?�6�?������<����m����� y�<�B�=K@	��@�J�78��ɾ��
��-��R���(��>��@���3s�>pl4�c��ο�ǅ��;�kf�!�?�#�>��Dc����l�o"s�H���F�}����>0@>.�3�F�"�Z���-����>p�<٘�>�<��룾�̾ɚ�<��>���>t��>�ۍ���־�ǔ?{��lοd�����N$?_��?X�?m�?j������Ȍ����^=��e?F�y?�7z?� �������@>d?�8Ǿ.0/��(�S*V�&�!>��I?��l>:@�(�<�:^=���>�@�>�R��齿������1���?�{�?��z�>���?e�E?� ����A���41�Gj�<�I?y�.>�˽bS��B��cR�ho�>���>R >�u �*�_??da���p��-���Ž}ݡ>z0��\�o:����We�l웿[x�<��?�a�?:(�?����#���$?��>�l��rkǾ���<,Z�>�Z�>3YN>��a�Z-v>ȩ�{�:���>]��?Xz�?�o?Ɠ���ڦ�.�>y�}?��>K��?���=�5�>�3�=�Ͱ����FT#>5A�=l�>��?o�M?��>�_�=�y8��/�ăF���Q�$����C��O�>}�a?�oL?��c>d���z�/�0] ��-νL02����5UA�}�/��<�9�5>�>>�>JD��Ӿ��?Np�9�ؿ j��p'��54?/��>�?����t�����;_?Qz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�>;�>�I�>?�Խ����\�����7>1�B?Y��D��t�o�x�>���?
�@�ծ?ii��	?���P��Ua~����7�U��=��7?�0��z>���>��=�nv�ݻ��W�s����>�B�?�{�?��>"�l?��o�O�B���1=6M�>Μk?�s?�Po���b�B>��?#������L��f?�
@~u@^�^?+��ݿ���d�Ӿ�V��x�>|_�=��'>�鮼�'/���(��Y����(>hXM>>Lw>!�9>ؚ�>�y�>��:>1�K>&�~��(�:��0�|���`[��R���\�	��ȯ�<����v�{��N��싾8T���+��Т�h������="�S?@�Q?m%o?��>.#����>�������<o.&����=�Y�>m�-?��K?��)?�N�=Yb���hd��ʁ�I��t���jv�>W�V>r%�>�-�>ε�>,y�;t�5>�`A>�3~>bM�=S#= �Ի�2�<��D>L�>���>�ߺ>�Ȋ>���<�W��n���N��d|s���J<�ԣ?Kh ���L��a�����Cq��:B	>*�?��p���S�ͿY���Ae7?�	��z��f����>��H?�B�?M@����䍾d���ge��q��e�*>����)m���A޾���=m'6?��i>%bp>��3���9�eP�q���R@�>�6?&�� �?��ru��I��Dܾ�oO>+�>����~������=}��g��x=_9?n�?�E��K����n�f���'W>B[>�=Tl�=��N>Cf�WcϽ�C�KN;=2a�=;	g>d�?�3>�*�=8K�>.���?i�a��>׀7>�h<>_�>?EK(?�>��f���L��`.*���l>���> �>��
>UD���=�i�>��d>�N��ț���$�C:��qL>���k�Nk��AN�=�J��Ŏ�=��=n����G��8�<�~?���䈿M�7e���lD?�+?� �=��F<��"�9 ���H��/�?O�@�l�?��	���V���?�@�?D��
��=p}�>G׫>1ξ��L�Ǳ? ƽ�Ƣ���	��(#�cS�?��?��/�1ʋ�%l�@4>k_%?��Ӿ��>���H��&��^�u���$=�>HFH?u���W�V��e>���	?n�?��� ���C�ȿ�Xv����>��?�Ք?Ĵm��+��L@�K��>��?'�Y?(h>�jھ�Z���>hZ@?��Q?c�>kv�L'��#?���?3?�oV>�g�?g�g?M��>�
'=�K��֬����>T3���?�d>e��G�3�Ȝs�������X��Մ�#�>��=�E�>�$g�o��9|0>��p��<���Y?��/�>N�Y>��>m�>��?���>0�>͉�<N>����ɩ�3�J?il�?��2��͂��V�=�5>ar��z�>��`?��w>����&��>.d?=�?�5�?  ?��پE
��7{���妾,)�=w��=dE�>�[�>wGf=��z>����[D�6�>�u>���(�2x��Ů>�%
�="�4?���>H��=��?�^?�˨>���>�B*�8T��!�E���M>�P�>�0?��?dX?�'�r�%�)���^[����`����>۵}?�1?޻�>H-���ՙ��8>n�B�N�� �?�v?�l)���C?a�v?�4%?`�+?o*�>��+���뾼��~>r%?:�-���E��U:�~�}�?#V?�X�>�����q0�����,�v����?�:?�?� ��s�x��Ѥ��<��ۻR"��ô;i��=��T>�O>�����>7�)>>=X�^��0��̑ﻦ��<�L�>~F>��&����= =,?'�G�ۃ�q�=K�r�xD���>�IL>.��m�^?�k=��{�����x�� 	U�� �?��?8k�?���D�h��$=?!�?k	?m"�>lJ��~޾��� Pw�{~x��w�S�>%��>�l���N���ř��rF���Ž�h*�)�>�	?��%?=(�>�E�>P��>B���������D��q�F�O���?�����S�þ�\
<II�=~�۾�� �ꊘ>>�=�&�>/Z? �g=���>+ћ>D��Z��>}>�<�
�>�u�=p�>�3=��>���=�u���?R?����r�'����Bz���B?�2e?��>�9{��腿��g{?w��?��?�qo>��h���*��	?���>�&~��{	?y�2=�q2�_�<�ɲ�,�������(�|�>Xpݽ��9��gK��Ne�z?�?]�G�g�̾TK½�s���M�9n^�?f�8?�}/�3�8��g��y���9�_/�<�S�,�R���E��Ec�M���|������X�,Z >�,?:0�?4R�[h۾>M������\>���J>Nx�>`��>�$'?��=��5�(2'���z�/�������b�>"�?e�>�pA?�:?�M?ՂE?��o>T�>�������>+�q��h�>h��>��"?>�+?G,?�w?,)?�3>��9�����ܾ� ?�!?dH?�>?��>�{f�s&2���9l�t���lr|�Q=��;���î�F�,=��`>:�? �6�As;�����_>X#A?�?���>���@�����9�>�?�(�>�M�DGm�E�����>2ق?���=�C>Q��=��<�wz<_b
>��n��f�=W�<h���X=�s>��	<�����k=��ȼf��=Sa)>�o�>T�?���>Ic�>x2��� �q���O�=XY>e1S>,->.Mپ�z���$����g��Wy>�s�?�u�?�wf=iO�=n��=咠��^������	��F�<B�?�I#?VT?���?��=?V#?c�>��C���W�����R�?P9.?A�n>�������=����$?�o�>�+Y�x!7���*���ʾl�-����=��5��{��嫿|s<����=�U
�ZW���#�?Su�?"���c?�7G��i���)���??���>Wi�>.J�>�@��5[�p�#��`=l�?�kV?<��>�wO?�-q?<Q?�Gt>K��­�̮��i1|=a�2>��J?��?0��?��n?��>���=�������8�U������'����ۂ=��M>ǉ>��>��>�3s=�-彬��>tN�'�=�)Z>�^�>Л�> ��>��->��b���G?���>��������ˤ�螃� f<���u?ܣ�?��+?9=�z�y�E�6������>zs�?J�?#*?��S�ݯ�=�bռ6趾��q�;�>��>�9�>��=$F=�>��>�q�>8S�1I��k8��!O�?�F?ި�=ZHѿ�x�����34����&>�p���,���7�u͏����=(��B�E=Ųk��'��ƾ��P�q���$\���6_�c��>,� >Ș=��;�x�:�d)=KA�=mZ;n�O��7�'m��=?i1��"��V��������K=>��=�3x���¾$�q?��P?�"7?s�>?� �>�2�=�4���q�>"ɽ�?"�>����پ��@�%o���0��#	���f¾�a�;t|���=�`^�6o>b[C>]��=��<�n�=�e�=���=5 ��
�;=G��=Bx�=�Ý=ug�=��'>
��=�6w?A��������4Q�$Z罄�:?�8�>�{�=T�ƾS@?��>>�2������]b��-?}��?�T�?'�?�ti��d�>H��!厽Do�=����n=2>q��=��2�t��>��J>����J������4�?��@ٞ??�ዿТϿ�`/>�8>�>��R���1�&�\�:�`�1�W�E�!?�F;��4;p_�>�%�=w�޾�ž�&=CP4>[�a=����[���=�'{�8q:=X7j=��>�E>�ý=렲����=%�J=�`�=`#O>��j�!�8��Y2���9=�Q�=b�a>A
)>��>�?�T6?�u?Iظ>e�#��3�궾�܎>�|>�[�>_�ϻ~>"�|>�&?:
;?��E?E��>Yv�<���>V�>��8��l�7ܾ`��p�=�|?�V�?���>���<�P���~-�DA���N�C�?+n&?e?��y>+������;��� �y��=��;6k=͖/�,"���=��H��3�=��=>8�d>xA^>c�>�t�>���=�YI>��>Q}1>,���ǧ�<�;�@B=��#=��<P�`�kU�����5�<ѿ�<�xǽ�����?��(B=j9.=�ǧ����=�3�>�	&>p��>��=�ݯ�um,>Ub����J�@ۮ=F��@�@�a�K�|�k�,�?�6�U�:>qhU>c^u�����G?B
^>�!G>J��?�\t?�>����о���7�g�xL`�8¿=���=�;���9��J^��cI��̾�O�>�ID>���>a=[>ƌ@�W�'���H>)S�
+����>��Ծ���=|9�;b��ْ��1��Z	�w^>siW?�銿�	z>"Y?^3?Cd�?���>q=��5�TS6>R��a���E	�p�����=y+?�:? ]�>��e�I��G̾o��N�>�0I���O�V���,�0�U��]˷�R��>U󪾣�оb$3�Cg��3�����B��Gr�m��>s�O?��?l1b�W��JSO����=���p?�}g?�>�I?�B?$��x|��j��Y��=��n?v��?;�?�>n�=C<����>܃	?N�?�q�?+Ns?�e;�L��>^3;�a>�����=3�>��=�A�=6�
?.9?�
?�a���	������^�~�=	Z�=�ǐ>���>d]n>4��=!�p=�`�=xt]>O�>���>5�i>
��>2��>(������-?s->Cx>p�@?!O�>�u�=)�����	�\�޽���ל���½꯻f�彗ŀ�9�>��K<�+�>띾�K�?�^>�$�� ?�,��7M��o0>��=�l߽��>woC>O�>,��>x?>3�k>#/>u=;=C�ƾ�j>p���a!��L�>�Q��	;:u�>f���\�"��T����&A�/u��Ұ��#�i��Ɓ���A�S�+<͒�?���(�h��0�h��qT
?A��><r-?&d��G4�&��=�>
O�>���mZ���^���4ܾDf�?&Y�? c>Kz�>�X?
c?O0�
n0�.�Z��u�b�@��id���_�L荿t>���#�±���P_?��x? A?A:�<��z>�?� &�-����w�>�/��V:��:=Tu�>�V��Z�_��XҾ�ľ�g�!�F>�_o?0߃?�=?�
W�t�m�/$'>E�:?��1?Mt?��1?m�;?��� �$?e3>@?�l?	J5?8�.?��
?�1>���=]:���(=kC��=슾�ѽKkʽ���`)4=.{=�ȸɊ
<_~=���<m�qټD�;���T��<)X:=9�=J�=��>v�\?���>�b�>а7?�k��9��9����.?Q�+=�O��H\��{��P��8w>��i?�n�?ӳY?*�b>��A��qA��>�4�>�\%>ʭ\>ޯ>�3�\�C�$ �=�>�X>X�=��Z�3���D	�i�����<R�>m�>�?f>	=%��>9U}���g�\��=��>��Hξf�R�H�1h-��1���e�>!0;?�I?k�>�$ﾵK�*Ki���?��R?��[?�fq?4�Y>��뾉y��L7�`09��v>C���bѾ ������>L���<��>�� ���k,4=`6־�¼,�����f�!��|�>�k?�cq>�����#��:p=S".>M��>�9���'�ln���N���vz?�UǼ���)Ԁ��e�¥=�_�>��?Z.���;ݤ;�e���Y>���>w��>��U�1%վw�d��R�u߇>�6E?�R_? �?q�����s��C����cH����ڼ�#?�ܫ>f�?9�<>M$�=�����u���d�rdF���>3�>���W/H��=B�J{$�≋>��?[�>gb?�WR?��
?R`?p*? �?H�>�X��s�����??��|?�iz� 󭾌�.���!�s��?�?��\?�}��>�
?�{9?|&?��P?��7?��f��پ�s@��ׂ>���>�Jo��٪����>gQ?e�>2�?C��?��r>�(M�������>3��>.	>"�-?�?c?$!�>�>5=����X�=����Z׃?4q5?i�?�̻�>��>�D�>���>h�>�Dt>E�Z�"X�>�bn?��T? ń?���?Fn=�����2�\ �:t6)�r0�79ʽK]==
����<t-ڽR乆����U;�ع�*ǽ7'F=mz�=��.����>���>������I>K���w%%��L>ͭ�X������A�-{�=z�M>�:?N��>��0��U�={	�>��>���T;,?��?k�?�J�<�\H��]��i�Q�C��>s�I?R�>�x�����hkz����=w w?��h?���-ƾ�d?=v\?Vz�R�>���þ:g�����1S?p+?�8r�[6�>Ǫ{?N�o?;�>=0S��sd��%����^���u����=vb�>���i��.�>�O8?N��>!5e>�i>>��җx�����?�-�?z��?�q�?k>��j���ܿ�_��nC��l-^?��>�}����"?�	���Ͼ�U��ZΎ��7�A⪾O��L��}��6%�Ã���ֽ|ѻ=�?��r?Esq?W�_?�� �4Ed��e^����MV����U����E�R�D���C���n��Z��[���
���XF=��W�;eC�%��?�6?����>����R�7�Ⱦ3}>�0˾�P���<���O�#�>:y�[�1�e���Ӻ�Ɔ-?�gl>�U ?ߴS?R�p���p���]���[� �㾪�>\;�>�>�q�>�����7p��^-�i4��N�<�[Ͻ�x�>��^?�
T?�wV?����G�
�������=��Ǿ��>r�>�/>21��0������$D�5U�v�⾸B����#�m^�=�>?�E�=���>���?;~?�8��w귾�BQ�0s[���>�*?���>��>�#ݽ�� ���>6�l?h��>;Ϡ>K+����!�&|�_�ʽ���>���>�>(q>�,��8\��3���W�� @9�z��=5{h?�p���a�F�>�R?g8:9HY<̮�>�u���!��I��'���>�N?v'�=�;>/ž.���Z{��	��`�Z?U/?�=�e�R��Έ>��L?��>IH{>���?�K�>��K�z=
��A�?���?�>��?Sj0?�75�<�꾝��"սB�i� N�>ro�>�'�=���� T�{���5��o�=yV*>9�����=�=��y���=��̽	.�=M̿� N����z¾��� ���ʾ��ֽ���%G����r��l��H��k�\½U9e����������g����?���?�߯��IS=ب�f8��`*��l!?I§�����&5 �
i���r�@ž�k�����#����q�V�4?r��O�ĿOҟ�}�پ��?�9??��u?��$����m�����A���b�=&O��ō��f˿5����IT?�n�> !������>g�=|�=${>je˾5}��m`�=���>�8?��?�ƾ�K̿�iÿp���G�?\�@}C?��#�}I�O=B��>JN
?��B>B�+�'j��/��<��>���?�ߍ? <�=V��	e?�#�;��G�(�����=7�=	�4=�u�H�T>b9�>"���E� ⷽ&c.>[�>������^�f���;�4p>%l��埽5Մ?-{\��f���/��T��U>��T?+�>�9�=��,?H7H�a}Ͽ�\��*a?�0�?��?�(?Zۿ��ؚ>��ܾ��M?WD6?���>�d&��t����=�8�$���g���&V�P��=I��>)�>��,�����O�}I����=�����~Ŀ�y(��$�	��=Ԉa=�彀���ʻ̽K��=J��'�h���|�|��=\��=�>`Y>Fz>��8>��V?�m?���>Xe>�(�I�~��߾y��<�x���Z�Q�l�ݤp��U�ƙ���Oؾo����)����j���=��d�=R��r��:� �?�b�V�F���.?d�#>+�ʾ��M�� <"ʾ||����������2̾�1�%3n��ҟ?��A?�녿��V���������W?���n���Ӭ�Ӝ�=����#�=MS�>nŢ=���y?3��tS��e0?mn ?w��s\���>��)�ڽ��&?�>�;� ��>��S?9�2��G> ��>\�2>���>Gװ>sE��\vιmɽ�IE?��X?��m���T��`7>Sɾ��������>g�ʽ3��ϋ >9&c;o�Ͼ�w��ZA=LǼ�+W?z��>��)���o[�����==��x?��?��>�hk?��B?���<'O����S����Mw==�W?i?^�>�r���оz��ֶ5?,�e?��N>�}h����0�.�hX��?r�n?�_?���{}��������e6?��v?s^�ws�����D�V�e=�>�[�>���>��9��k�>�>?�#��G������yY4�%Þ?��@���?��;<��L��=�;?i\�>��O��>ƾ�z������/�q=�"�>���~ev����R,�c�8?ܠ�?���>������7�>+��WO�?0��?8ξ���}����r�\������=;ߙ=��<g���6����<���ھˍ�[���08�r��>�@|L�r^�>p�9��U꿩�̿>���̾5%�v-?�̪>[�'P��3s�C!p�mQQ�"�5��o�k$�>d�=8ل�b�b��W��k@�z����*?n���De>�"!��ޱ���N�*Δ=`�>��>��>��e�����!�?�6þ�ҿ�(���䘾R?���?T΁?��I?�����.��@��A�=���?�?�o�?�&�R�'�|�W��j?ﳪ��7`��4���E�"�S>\B3?���>x�-��3�=V>S��>X�>��.�h�Ŀ�ﶿD[��E��?ey�?
�꾬B�>B��?S�+?���������@+��X�9=A?�/>�����d!��Q=�⮒�[e
?�0?M���h���_?��a�8�p���-��ƽ<ۡ>S�0��c\�-9��x��rXe����?y����? ^�?t�?��� #��5%?��>�����9Ǿ���<
��><)�>p+N>�K_���u>a�'�:��h	>���?�~�?7j?��������6V>��}?�S�>)��?B��=��>b�=!����tr���>��=��1?�TX?;��>��.>=N⽑H/�IF:�� E�G���B�%�>�7i?ŸE?�uT>K5���U%�=�w�ۍ!�ѿ��	z��c�T\��jH>Z�>�>Q9(������?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�e��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?[Qo���i�B>��?"������L��f?�
@u@a�^?*5�޿5���˾���*��=Z�=�<�=�g���ϼ.h>rR=�׼�_t=��>�L�>G�j>�1�=6q<>Zb>`#��l�$�V����Ȑ���@��z���O���=��舾���\�{���¾X ����˼�ܽg����H~��ký�� >��W?/\H?l?|��>A����=�����;x�g�!�=oA�>3$?ӨU??3?aC	=1���X�2�����aQ�g)�>NXE>=��>0C�>儭>������}>[>$ރ>w�;=���<������=�.U>��>JP�> ��>%��>�pQ��֩�B���d������}�=(��?�6�J�m�qž��Ω>,E?�T>�!���ֿ�0��VA>?Da��6S*��ʓ���>�9?��?u�<�����^��͞>j���I�Y�7>}E�"��P@&����=�
,?ށg>9xt>��3� o8���P�:���}>.D6?���Te9�wku�#�H�S�ݾ9TN>ݸ�>�>�$r�8��8�~�Kmi��H{=�Q:?�k?�ﳽ�㰾�`u�b����zQ>:m\>�4=��=3�L>��f��ȽDI�a�,=�=�=	`>��?rN->��=��>����SN��>�sA>�,>��??�0%?/w�����څ����,��sx>w�>Tn�>��>e�J��<�=���>T/a>�����⃽����>�o�W>�>}�[�`��=v���=������=���=TW��ҽ<� �)=��~?�x��_䈿z$��\���iD?�,?�=E7J<T�"�\ ���C����?��@Zj�?y	�˞V���?X;�?���ſ�=�h�>Eԫ>�ξAtL���??.ƽ����s�	��:#��L�?�?T�/��ʋ��l�vh>�X%?U�ӾPh�>{x��Z�������u�x�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?�ٓ>R�?�[k?8��>b�=�Hl��ռ���{���j>�y��,��>MD�>��þ�f��t�v�m����=����S>��="*�>�I�[���B�#>��H<�y���=uP�>�=>�a�>6�>��>���>K�;>�Ң���.���_���R?8��?�z,�W�i���=p>h�k�߭ ?PD?ҚQ�����t�>G4P?Dg�?1u^?֣>]H⾫I��D����ƾ3A3�їM>�}?�>���X(�=����������6>^�>��=���Q���s=+l�>\?e�>X��<	�"?�?�>���>��6�RǦ��g��%�=��>��?��?9?(�t�K�/����e��ܾW��2>�ZM?�A?�"�>�G������R�O>|j�������܁?7Jz?�,����>�`?�+?	t?���>7�=uA྇̑���L>��-?�e�$�Q��Y/����k��>e?<�?�0�Vb�q�=�&4����P)?RS?�4'?��������Ѿ��=3u���N}��9|��V�:">E>k~��>D;=�<>��=K�������ǽ�!��sG%>�E);G+��Q:>k9,?��E��҃�|�=\�r�oD���>EL>�����^?�R=��{�:��w��x�T�� �?H��? m�?Y���p�h��%=?P�?�?�+�>�N���l޾���HAw��~x�&x���>��>D�m�'�<���*���*E��?�Ž��)��b�>��?��;?��>�-R>�>�1E���)�%�о�K�J�o��m)�Q�V��(��i&�����.^�i�YǾ��M�W��>oh����>M'?->�P�>�@�>��i=�-E>�d�>��f>8��>~�A>Y�>�>�Q
>�6B<fjR?�⽾	(�6������sB?�Dc?
>�>�T�@I�����$?\��?w��?՜v>tyg�'�)���?��>�b��;i
?��9=��k��<����y�� ��&�'�>��ս��9���L���d�P
?#?�k~�*�˾)н��/�1�k;=��?�zr?{Z��~[��js��=A��U�v6>W��)���;��!L�����to��,�*<�(?27�?fa�0aᾐȐ��އ���E��H=QQ�>c�>4�.?I�>1�������L���7�L����u�>.�n?��>��K?�;:?��O?�K?��>�¤>y�/+�>p��� �>���>��4?��-?>�0?��?av-?��j>�����t���оpR?dU?��?�S?GX?1�������{o�f�c��k��_l��]=~�<��ǽ�3^���H="i^>�T?(��!�8�����*k>Z7?���>7��>���\#���<�>�
?�=�>I����ur�N]�a^�> ��?R���[=k�)>N��=������κiY�=����/ݐ=a��K�;�1L<e��=V��=�yt�������:9 �;���<�n�>6�?o��>�L�>�5��6� �8��}k�=�Y>S>�>�Iپ�|��K$��i�g�8[y>�w�?�y�?��f=� �=-��=�t���N��b��!���k?�<��?FI#?]UT?ڒ�?��=?�n#?��>�.�%L��:\�����ܰ?�X8?8U>�6���ﾓs��¿0��R6?,2�>�i��Dؼ��^� ���u�>�S��ʈ�m����MR��'>�v�Q������?�?�5���3��s��^��e�B��D?=]">ky�>��?�>���k��6�u+>��'?8B?��>�Q?�z?�rR?��_>_v@��خ��.��k��<,N�=�&D?��?`ǈ?��g?�d�>{K>#�M��Qپ����U �-���W�n�#g�=�V;>R	�>���>}��>�
�=}�n��l���1�<2�=3�z>~��>��>��> �u>3�=\�F?	�>�龾*���o��0mk�'}�%�p?��?�u%?"�=P	�%?�8�ﾟ��>�?P��?d�+?̟U�`7�=�*��6c���Og�ܸ>@�>���>6߁=��o=��1>T��>�պ>�?���k^<�+{��?��D?���=e1ƿ�Ir�T:s�����w�h<�%��T�e����� [���=z엾
A��a���Z�FD���Փ�醵�W��L�x���>
Ċ=�v�=���=j��<�&��c�<G=��<��
=m�l�ӰY<EZ0��{ػ�t��3-g���P< rL=~p*��3ʾ+}?�5I?�i+?��B?�2u>M�>$s3��ݖ>�u���*?,�V>��Z�������9��b���ϕ��c׾�E־�?c�Ş�ϣ	>�iL��6>�h8>O�=�c�<���=��y=6��=I�H��|=��=ؤ�=�İ=&��=�>��>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��7>Q|>_�R��b1���\�b�#�Z�n�!?I;��̾�U�>f��=`1߾rƾT�0=856>B�b=bJ��\\�T
�=�#y��>=��l=h��>0D>?l�=\"�����=!qI=�0�=�$O>������7��W+���1=�x�=��b>7�&>���>�.?�"?Ǿ\?��>��N<�Ӿ;��o-�>��/=���>�la=�r<�P�>,oY?�A?&�b?���>a=3W>i�>�� ��H�?2��(⋾z�$>zq?��?��>+�= D���&�݅m�Z�	�223?57I?B 6?�S�>�V
�)��3<��=�����n��F���;!+�o�Ѽ7� ���=?����̛>$��>;��=r`�=���>Cՠ>�#�>>%>�h�;|˾=�f�=w_/>���\��;��=s�>y������ܖ=�_��1R�@h�Ѭt=��=��y�SD>���>�ڜ>:�>�L=����Q �=�7�
_P�˪�l`̾��T�ea����AR6�_�V��)>V>�� ��P���P�>D�|>�֒>ܽ�?lҁ?�l�>��=�� ��o��ys�x�$֟=SLR������F�5�4���@�]���>�+k=4J�>��>��]��*4��B�=2|"��k&�_y�>�?�� �q�E���\�짿,g������,�S?0���J�>!��??�m?ڏ�?1.�>�j*��.Ծ3J>؝�������!ɾ)�r���+?7J!?���>�T���e}�KW��ߑ��g�>E�<J�Pœ� 5�jm9<�2���c�>�ԯ�σ۾��3�?c��bT���8Y���l����>X
G?���?��7��C���pZ�_������>��a?�f�>�H�>Ol?����p����fM>�)m?;�?޵�?�}�=o8��[�>e�>��>I�?���?݈�?{A`��?Mϐ�LHK>�	>U}Q>O������=<,�>�7?j�?c�)?Ѱ��ƃ3��s��1��>i�L=2�=�L;>�r�=�Y>��f<,�=bO�=�_l>C3�>�b>"eO�@k�=\Yo>F���4����2?�>�GX>�A?Ş�>���=��ӽH	�<�SK��B�(}��Y����
��m�a�-=�={W��4��>�uѿy{�?0�B>�����
?]!���ֽ^-3>��Z>�̀�G� ?��X>zֹ>v��>��y>=* >��t>E��=�.Ӿe\>���Lh!��)C�X~R���Ѿq�z>����&����6����fI��\��%h��j��/��TF=�}>�<C�?j���Ŷk���)�*��҉?U[�>�6?�֌�Ј�ђ>��>Oэ>k\�������ˍ��cᾝ�?���?�7c>k�>��W?͜?��1��3��rZ�b�u�k'A��e�ʼ`�፿!�����
�0
����_?�x?�wA?9�<�0z>��?��%�Dҏ��,�>�/��#;�v<=�*�>(�� �`�ȫӾ�þ�;�lKF>C�o?�%�?[?MV��尿�W>��0?yp!?8{?E�9?�5B?:0 ��%?��>��?'?v�.?h"?g�?TZq>I >v�;�'�=���%���x��/�U�i�/�<l<q=r�ü�ߨ����=�V=����>A�2��ؕt;��<� =�d�=/�>�1f>:U�?ޭ?���>6
K?�F�=g����֝���B?w
�<�����_e�k>�������|>�p?<P�?�}?���>ѥ�� �Q��uT>�mn>�X�>)��=L�?��Ƚї��W��E"���YG>A�>��,���龡�ݾ��F�ܫ�p|>ֽ�>�y�>k8��J�$>6g��^�p�OIW>�G�4:���K[�wQE���*�� u����>��L?��?�̦=wm�J)����f��$?n'>?GN?�y?
�=�=ܾ��7���P�^�&� (�>�I�<6��1�����H;�$#Y;�x>����aȁ�R�B>"��ʰʾ��l�L�[����?f>i�"��������뤾�!���>��>w���@����i樿�c?�jL=%��Y� �#P=�Г>NZ�>ױ���=��#�":��|#C>��>���=�\��x��-�;��ž�~�>t�@?��\?�Ї?��o�����zJ��G�?��|û�G=?�$?���>�J>m�=n����
��k]�yt)���>��>n4���:��ٔ�?����	���l>��?B��=��>��Y?�f?��f?K�R?��?�A�>�@ �.���,?)r?�HZ=y��i�ݽ-�/���B���>��?��m�1,>j�0?��*?N=?\�s?���>��=C�4g��Ú>wxZ>�fA�t_���q:>�lJ?�y�>�Ke?��n?%�>r�<���Ҿ���b,>�0>�?��?�?�f>8�>-����w�=g��>^$e?���?�p?9.=���>��N>���>o�=��>�W�>�?o`K?��y?�pG?���>�x	=��޽���?� �0M6�ޓG�9h&�'�ƻ��r��Cq�4%0�w�<Z5V�0;���F�"���E9���b=F��<v9�>R?s>ޔ����0>�ž!�;�@>�Σ�/�������`;�{�=�ހ>p!?�#�> �#��Ԓ=t��>��>���(?2�?�<?�� ;t�b��۾T�K���>SB?5<�=�l��h����u�ޅf=
�m?�{^?\W������_?XR?|�ξ��U-��Z�������2z?H�?�jI����>�@�?I�o?�l?ݼ�V�?0��e�_��O��:�(>Ł�>.��qs���>n$F?*K�>r�Z>�O�<�/ɾ�Ӕ��4��W#(?��?T0�?�=�?�>��\���i��������^?=r�>L����z"?��0��*ϾV`��Ҿ��a0߾���������o1����$�涂�d�ӽ��=��?�Ps?�&q?�_?�� ���c��^�o�~���V��@��=��`D���D�C�R"m��d���������J*=�,{���?���?�'?I�Z�˛�>�қ�f�+��5�=���^���>j�<IO>�Lɼ��J�o�����ƈ?�A�>�3�>s�H?�xH�
�H��6��1��8�Q>/��>��>}��>1<`@/��T��$�Ⱦ�G��e���Zv>�kc?W�K?��n?:F��H1�=���.�!�\).�dR���C>a�>2��>XW����/&��F>���r����A����	�S}=�2?��>���>�C�?��?�J	�������x�]1�`��<1\�>SWi?�y�>��>��н�!����> �l?[��>e�>�����^!�0�{���ʽS�>��>��>��o>��,��+\��n��[���9�k��=ܰh?Ԅ����`���>fR?�)�:�yH<i�>�&w�Z�!���7�'�	>rt?���=��;>Jožz�|�{�W7��p)?uK?�����)�*k�>�� ?�t�>3�>��?U��>�ž�Z�;N�?�^?��K?wa@?�X�>j�<'�ɽ�˽6�#�4l.=��>+Z>g�q=�#�=>��Y�M&���D=�ù=��k�ʽ|z;����L<<���<5�4>gGѿP7>�T��|b�`Fᾃ� ��5��_����b�:�\�2�`�X���殾X����6�W��(k�ٯ��
}���"�?���?�6��@�w�[����������V�>��۾�н�����ʽ��2�	5���`��R���r���o��Us��A8?����%ÿ�l������9�>�c"?X??�[+�l$��.�M��=6#�>HBͽ?>�핿�eؿ�e��?�S?툿>� Ӿ�K=�m�>o�O>�{>��>�V��!F�E�U=e�?��?�F�>�>ľ��ƿe~����.j�?=�@�zA?��(�t��U=���>��	?��?>1�}>� .��88�>�8�?��?
-M=�W���	�"le?Ъ�;!�F���ֻ���=�ͤ=��=�@��rJ>�}�>"�� (A�^�۽ڵ4>B��>��"����s�^��Ǿ<��]>��ս����4Մ?{\��f���/�U���T>�T?�+�>$>�=��,?`7H�U}Ͽ��\��*a?�0�?��?D�(?�ڿ��ؚ>l�ܾW�M?]D6?��>�d&���t�Ѕ�=�+�\i��c�㾭&V����=���>@�>��,������O�:�����=����3���Ei
�w���v�=�i�<g��$����=(ʝ��p�x��������>�~D=3[>>�6�>�h>Dib>/�d?N�y?U?�{I>I!W������k̾��=H.h��5e����@N���?�����K��|�<�K���k�(�3��z�=��B���������d��O��,?�~�=����,5����<���r�����;����n�=�Ax�x�?��7?,-����B���JH�V��wQ?�U��۾L7��q�=v�=�G=�o�>��=������7�E�C�?/0?l_?�[��*퐾[�,>iv ��k�<�O,?qG?S��;�5�>%?��%��v὜�_>��4>v¢>�X�>��>D5��|Nؽ��?�;T?A��kg���Z�>I＾�iz���Q=��>j�2��'���|T>2�c<6����e��J����<G+W?���>~ *���u���S��z==��x?�|?y-�>�qk?��B?z��<�S����S��"��Iv=�W?/i?��>����C�Ͼ,���V�5?פe? O>�h������.�z]�a?��n?CO?����k}�e������p6?4�v?dd^�k������EW�E"�>���>J�>F�9� ��>�b>?�#�y;��򡿿�S4�Ҟ?��@z��?��A<Ţ���=xc?���>h�N�2ƾ�=��lP��"�p=L*�>�0��dVv�A ��d,�J�8?�u�?���>+R���t����=P暾�l�?�^�?{ﲾf!j<K��no�:^�<,�=�GĽ~�b��4���C���پ��'���o�X���>A�@���z?�k����l�ʿ����O��-��m�0?���>jc�E�⾑�\�ïf�.Q�?�9���D����>�
>�je�x���&m{��a)����=t��>�H�=ly��5?k��/{�+Z=����42�>�3?��>I\��	�����?Mg��eÿ[����_��c9?�ؿ?�gP?��-?V�>��_����=\�=��)?`0?v4�?f��=�a=P�<-h?�����J�DZ��X��ם�ZU%?���>��(��z;>(��>�>k�<N�s�ȿq�����֧�?���?Я�����>]��?�wH?�C��0���3Ⱦ�V۾���=�&'?w�>�4��R�K�q�K�-w����>��K?�,�=����]�_?+�a�N�p���-���ƽ�ۡ>��0��e\�N�����Xe����@y����?N^�?i�?Ե�� #�g6%?�>d����8Ǿ��<���>�(�>*N>cH_���u>����:�i	>���?�~�?Qj?���� ����U>
�}?w)�>�
�?���=�+�>���=	˰�-�A�KZ$>,2�=N�F��^?�M?|��>ȷ�=��7���.��9F�YR��O��C�% �>��a?�xL?�Jb>mŸ�&#0�L� ���ͽ�;2��T鼤�?�n�-�k���.4>;�=>j>��E�0�Ҿ��?Mp�5�ؿ�i��Hp'��54?4��>�?��f�t� ���;_?Sz�>�6�,���%���B�]��?�G�?6�?��׾2Q̼<>6�>�I�>f�Խ���@�����7>9�B?3��D��t�o�c�>���?	�@�ծ?Wi��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?kQo���i�B>��?"������L��f?�
@u@a�^?*�Ϳ�Y���%�;浾t�>�r�=��>��1���0=A��>T&�yQ��~᛽�>[��=!g>.�U>�R�>O�>sx���"�/���哿�"����О���v�0��|�ʼZ�*�il��a���|S=(i`�m�[��S&��zF�X�h��=�T?R-O?^�k?�?��s��� >&��*�=�EN��~O=+��>D@5?_LI?�.?`6�=����6f�g)���O��΁��_�>,�N>t�>���>[�>�9<x_C>�(>TZ{>{'>_ =�3�y��<4�I>��>"��>�˵>�^�>�˺=ⲿOG��@s�죨��("�(��?�O�'+�ҵj���C�N:���=��?���z@��ʿ�朿�5I?v������2ľ]�>�??K5�?r�<�����?������f��&7���=P5V��Da�,O��L^>��?�h>tt>T�3���8��$P�����Gz>�<6?;k����<��3u��uG���پ�oL>G��>v�Q�)��	��Z�~�\g��z=ߖ9?�X?����؉��9Ro�т��[�R>�Z>s=+D�=��K>>�r���нA�G���#=|��=C�`>�N?��+>;�=5ԣ>�o��'�O�M{�>�~B>K�+>��??6%?/��A^��d���8.��v>�H�>G*�>�U>�WJ���=^s�>� b>����ヽ�����?�=�W>�}��O_�`*u��'y=�����}�=�m�=�@ ���<�)+%=�~?���(䈿��e���lD?S+?^ �=��F<��"�E ���H��G�?r�@m�?��	��V�?�?�@�?��I��=}�>׫>�ξ�L��?��Ž4Ǣ�Ȕ	�/)#�iS�?��?��/�Zʋ�;l�}6>�^%?��Ӿhq�>�~�T[��y����u��h#=M��>�6H?;c��b�O���=�_s
?�?�S�����ȿ�v����>� �?Y�?F�m�*=��<@���>���?�nY?�Oi>r_۾�ZZ��z�>V�@?�R?0�>�;�&�'���?�۶?X��?��I>�\�?�Us?��>}�s�`�/����Sh����x=���;偒>l�>Y����TF� �z��Ąj�n���'e>��(=�l�>�v��滾�H�=����t����\�l�>�)p>8O>�$�>� ?,�>4 �>�=�}���y��>q���vD?�x?T�Ѿ�*U�ށK>�.=�����$?�1'?�鶾T�����>��c?���?:��?���>��쾒���8Ͼ�?�ɾ�˪=[H>��>D��>/*u<%M�=a)!�+�+��_ʽ�|>OU�t��& �8�M�%F�>�@�>zL>��(>�c?}�$?�P�>���>O&�	H��i;S��]�>�B�>�V?	��?:2?�Q�L�+�I������{�Q�ԁb>!N�?'�?!b�>Vo{��k��hn:��H��ƽ��p?A��?�l�}�2?�Z�?|J%?a�A?}� ?��绹m���<���>"�!?��
�[�@�]r&�rK�F?p#?�2�>�ۑ������2@����gv?��[?y�%?����+b�eƾ�E�<A�%�7ꃻ)T�;�7o�k�>�� >hl��S��=�'>چ�=�l�`K9���;ɷ�=�M�>;��=�@6�2����-?	��= ���w>Pa�c�%�:�>տ?�.&��o?&k�����>���̆����W6�?�*�?�y�?A��=�sd���{?Ǆ�?DH$?q"?\6Q��/��-��;׾Iܾ%֠���6> M+>�5��0��[��Ñ��uzv���������>DD�>v��>���>�>�>?��>?ͭ�)�A�n���H3 ��h�5� �+`�Q�2�0�.��J��Gҽ!|��a����|��^C�>�Q<��>ET?3e4>�7�>N~�>�B��`�b>�>8��>��?�i>�>j#�>�C=��h�eLR?�����'�l�辸Ű��!B?ibd?�'�>�Yj������� n?���?hn�?�v>{h��4+��V?F�>_	���d
?��:=�^����<�2��An��������ӗ�>�׽�:���L���f��J
?Q)?�ޏ��g̾��ֽ5_��)�=���?'�>?�4��pL���o���_�G5[�(F�<s������\%���d�������H����`���l=�r)?3p�?W��w�ξ�kK��.v�T�B��g>'?�G�>R� ?Ե>���d�F�ߪH�T�%����;�>ZɄ?g�y>*p`?OhG?�Y?��X?k��>,�>�ľv��>p��;�L�> �>�?�`?rn0?�w?A�'?�ҕ>npѽ���վɥ
?�?A�#?v?�x?=ў��J�y]�=�γ�Aye��H���r=4=n�������W�<@�j>��?*[�c�6�Nh����e>�7?�?�>��>WZ���k���V�<(v�>��?*��>�� �m�r������>f��?v��]H�<��+>o]�=ĳ��HF���S�=^?ļE+�=��q��/�|�)<��=S��=��n8�;4��;BI�;���<�t�>;�?��>�D�>@��X� �����b�=Y>�S>�> Eپ�}���$����g��Zy>Iw�?�z�?�f=��=ə�=�|��`U��&��$������<	�?�J#?�WT?���?��=?�i#?+�>5*�M��t^����� �?A.?�>�y���־�ը��b2�Q�?���>�Pc�T�6+%�++�����	�=�o3�1A��;߱�r:@�c��<�9������i�?֠?gL@��8�/!辗w�����}HC?���>O­>�7�>��)��h� ��	T>?�W?+�>ÍM?�x?"!`?
OR>�@��W��wA��\c<Es!>�M?��?K��?J�v?2��>̟>\�(��w���W���L���fn��U =x�Z>���>�%�>U�>p��=�������t&8�GS>$�>�  ?N��>���>JaX>V�/�-_U?6TZ>���\�!��-�_M�py�>�q�?�x�?u/?E	B���<�K�,rž._u>�`�?�n�?�a1?T���9s=rB<�a��#�<���>���>��n>g]�>�2L>��>>��>��>����r���'%�G=�]$?�?o�>�ſ&r���o�����&�<ؚ�� �f�𙽼�X��¢=ŗ�� ������;V��L��vɒ����'�I|�Y�>$�=�~�=CE�=�M�<���f�<	\I=^�:<G��<��j�X�w<E"1��bE������}���V<>;I=��s���þ!��?��Q?Y76?��N?Y�>�k>>K�ӽ�ڠ>n�W�r�?j&>�󟽠�Ѿ�u��ܯ��]�l�>T�������bt��᣾9�>��ڼMN>(1{>(>�:����=#��=�,�=m�L;��C="|�=���=���=�С=��=�e!>�6w?X�������4Q��Z罥�:?�8�>i{�=��ƾq@?~�>>�2������yb��-?���?�T�?>�??ti��d�>L���㎽�q�=H����=2>q��=w�2�T��>��J>���K��F����4�?��@��??�ዿТϿ7a/>Qk;>�->L�V�-�mP@�9�[�er�4T'?��4�����q>�M�=�Ͼ؆Ǿ|��=�M;>�;%=
�B��*_�-��=G�u��K	=p�a=�s>s�6>�x�=l���=3#9=��=^*M>ܝ򼚂}��啽��=��=|H>�])>$��>�?�/?Šb?��>T�m���о�h�����>镮=�|�>���=��A>�µ>��7?*�C?�J?���>
�u=Uܽ>�+�>�k-��>l�7������f=��?[�? ع>�6�</�D�_���<�u�սt�?Q�2?:.?ٞ>�0����{"]�vK���=i�#���r���gN5�0G=G\���LO���<�+?��L>��>���>�>��/>���>�sX>���=I�=M��-�,��k����=�/�=��.�^yK=^����=��=:�V<�5r��==jr��L>=�\�=�r?׌>t�>P��=aㅾ|M>��v�js.�(��<�ň�U�C��mk�S�}��������>�g�>E1�,�����?:Hu>� >�<�?*�?3$="L������旝���w�Y����c>cjj=O�,�eC���l��H=�E���]��>r{\>,Q�>!�!>�w1���2���/=U>Ѿ)R����>t���o�ٽӀ����������������o����=�gY?����
�=�as?FA?u�?&S"?s�ݽY!��rǽYh��>{b���0�
���>�G-?� ?d�>A�}�]��F̾D���ݷ>�@I���O�W�2�0���H̷�Ԍ�>������о�#3�eg��m���[�B��Lr�,�>�O?s�?a;b��W���TO�"���+���r?�{g?��>,K?�@?�)��z�q���o�=��n?̳�?�<�?D>�O����q>�/?cN?c��?Mƪ?���?�R����>oH>�K�=F����)<��K�F3�>�f>΀?�Ͽ>�?�!��
�qE�#{������N��k�=���>�>�v�=��=�>	>$>�>T3>y�y>�1>Ԅw=ը�>ز������l(?�2�=�ȅ>�3?��>dpQ=UYνk2<N잽`�R�����X������|;�"���m|=��漆��>p�Ŀ���?�"e>P��C�?����(���[>#U>
ý���>{�O>�,�>�i�>큩>LC*>a�>��>b���� >������@CN�U@d�������>K�;�j�m�ϾN	��х�]����la���^K��솽���?aR�B�m�I�$��&3��0?�)�>��&?���Zi�@>��>?��>?���{ ��Њ�s�¾fk�?�F�?J;c>��>l�W?�?��1��3��uZ���u�i(A�e�l�`��፿����t�
��	��V�_?��x?(yA?�M�<-9z>��?i�%�-ҏ�*�>g/�
';��;<=�+�>�)����`���Ӿ;�þ6��GF>T�o?%�?EY?UV�Q�P�&gg>dO9?i=@?��}?�@F?#�S?+�8�.�
?��I>ks�>�V?-\;??�>�R�>"�>pl�>
֗��,>�գ���Ͼ�x潵*��G�:�n=-<�O��N`0���	>g2�=��=E�s�(>�=Zt��e
��&9>K�G>�|�=�k�>�d??U��>$m=?N7����,������d/?/�h=�����3Y�������R>h?�w�?�i[?M*g>XI�wxJ��� >wˉ>��9>"dv>E��>�t���=�!�=F�>�H>��=^�W���u����s�����;��">���>�~>d%��45'>�z���+y�[�^>��M��x��6�Y�j�G�}�0�!�q����>StL?��?�Ι=1�!���Ff��)?��;?�KM?)}?I�=��ھ9� �J��U!�]`�>
n�<=,���䡿��9���޺F-o>�螾�B����>s�Ͼf|��w��6�.�/� t<X	��G�:>������ l�tr	>�+�>l#�ũ�|*���Oɿ$�}?��=]�農�A������"��e>�Q�>��0�����j�������!>6 �>@�=��ս����dCH�׋���>d�=?��c?��?�C���g���A�6�վq1���PM�R�?㈫>�B?٨H>JD�<S_о!3���S��1,����>d��>@�'�u�F�>/��[��J�#�+2	>���>�-�=�R�>��M?���>�??�r,?�~?��|>���;�� �%?�i�?�|�=�!��)�F���6���F��,�>�&?{	8���>l?a?�<#?��O?y?f,>Pn�Ӷ=����>�E�>BT�sR���xk>@M?|�>�[?�=�?�M>><�7�篾��w�(��=��=o�/?��"??�?��>���>D����V�=�H�>�	c?�&�?��o?�=�?��1>^��>3.�=�h�>��>��?iBO?Žs?��J?(��>��<!���9շ��Ss��X����;�BR<_y=� �VRq����1y�<���;�a���邼�$�G�\�����;�
�>��q>�"��0/>%�ľÞ��N8C>�	������#����7�}�=��~>�v?�ّ>��$���=ײ�>���>a�_�(??�?�P;�b�1�۾��J���>�aB?ߤ�=�3m�5����u��tw=Z%o?�1_?+�T�����ob?L�\?a��RJ:�nN¾s�h��6�g�O?�C?'H�^��>R�?�Mr?a��>�|e�3o��-��+�`��f��q�=��>���v2e��I�>kE6?���>�R>T�=Jܾx�kP����?���?Lݯ?߉?�&>5Go��߿�F���+����]?�o�>i���#?8���6�ϾE�������(���䫾�*�������$�-���Hmֽ�R�=�?�)s?�`q?��_?:z �s�c��*^����ڀV�=8�g-�V�E��E�rqC��n��c�m��8��G1G=���v
=�93�?��'?w�4����>^��5+뾧aξ�wD>���Z���=,����>=Ο[=�Gk�2��쯾C� ?��>fZ�>�;?�[��4>�_�0���6����N0>���>��>�x�>�e�!v'�� ܽ�ȾY|���ܽ$>ٗa?�/J?b~n?���:t0�~��EV!��@�ԡ���A>�B>".�>1�P� +���'��:�Olq�	��݌�[�e�f=�)?#�>�A�>���?�?˷	����{ǁ�pV5��@�<�[�>��[?C\�>���>�����h�>M)c?��>]�>%����"��$o��5����>�8�>���>�Մ>���:�L��͉������+�T��=x�i?M1t��K\��YX>?�;?��=XT�<�ow>:��x�ڧ�N�o�x��=�� ?Ϛ�<�]U>о�i��t�~�e.q��L)?u;?������*���}>�!?�s�>�%�>�%�? |�>\�¾��3��x?��^?EJ?2+A?�>��=�ܱ�GȽ�P'�j�)=��>�Z>�]l={��=Rg�t�[�#���D=�=kaӼt���U<�=���E<��<�r4>��ԿP�8���¾�����Ӿ؝�f��䵷��Q��b}��1ƾ�����!]���=��Խ7dO��➾2����1�?��?�|�A\x�2����|�b�o=�>����2��)����D��`^����K�������yI��Hj�cw�ۮ'?�&�\����)¿џ �� C?}[W?RM?�@��ge��O��ˎ>q'!>�i >3������ؠԿ=�o��-S?*&�>���h�;��>�Օ>&��>6t�>��8��j�T�a�
��>�3*?��>�>������ʵ�g�=��?�� @xKA?��&����[=8��>)?��;>��)�'��b��2��>�0�?�ԉ?��==E�U�H�.��,d?�;,
B�ۻ�!��=ʣ�=��<t��yI>�S�>��'��YG���ؽ�@->���>���?��X�F�<��S>�|ҽ����5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=u6�����{���&V�}��=[��>c�>,������O��I��U��=;j �L�ÿen#�x�ͪ�=�g-=ǅL��{��A�' ,����ߤ^�k佟��=-�3>�-t>�5�>�%?>�7>X�[?�r?��>�P>�9P�����ܾ���=\tw�I�����V�'���z�����jؾ�� �>�0Y��о�j<�'L�=XQ�)���P}!�Gb�X�G���-?p� >�IȾ�FM�t�<��ƾ���|�$�ƺ��4-̾sC3��cp���?��@?����ЛV�����q��>��&�V?�@ �}=�������=����!=�ߚ>o��=(⾾�2���R���1?c�?�ؾI��F�a>��,���>�( ?[�?����G>�*?��|�m��a�=�|,>��z>���>_z>�ȭ�$6м�8?SJ?�S@�񾀾�Z�>U�̾���� �2>h�8>��3f�=��>梂��6�����Y��=���1+T?�>\���C�_����d��\lC=�v?�?�;�>�n?��C?pN=y�ؾ�N���+�Y=�3O?�h?Ҁ
>Q>���Ծ驾B�7?,O_?->G�����۾*�2�;�� ?9�i?j�
?�jm<�/���������5?;n?:kM�Dʇ��K⾞W����U>�� ?��?��-��p?#D?A[��I��3���\g+��z�?��@Y,�?wVj�6쟽W�H>?+?�k��c����K�-ŭ�Ҽ����>����\�|�T�9�p���P^?�l�?�?Z�6�����"�=<���X��?:�?ݬ���:�<��zcj��- �/y�<1�=|%����!D�ס8�O�ƾ/�
����y��櫆>�@0������>�5��⿦�ο�Ѕ���̾l�r��2?qy�>��̽XǤ���i�f�s��wF�4!H����P�>1<>)���T瓾`\|��M;�<Q�����>@��Z�>�eS������,�u<�Ӓ>�m�>���>V&���ž��r�?!;���Ϳ�.���w��Y?21�?�߄?�??��;�cx�5ky���"��F?�jr?��X?N�1���W�(��x%e?�پT)[��mM��?�Fka>b�L?q��>��5<�=���=U6�>��>���1p��)g��ȅ���Q�?��?ױ̾|�?;��?c?�O�g>��ޓԾ�'��>���?�ʿ>���3�7���>����3?��o?��ļ�:�[�_?,�a�S�p���-��ƽ�ۡ>��0��e\�;M��U���Xe����@y����?F^�?`�?��� #�`6%?�>x����8ǾW�<���>)�>s*N>9H_�òu>����:�"i	>���?�~�?Kj?��������)V>�}?L�>x�?�d�=tD�>�7�=���"-����> i>��O�E�?�GN?���>Ǚ�=��7��1��LE��tP�.�O�B��
�>~�^?��H?@o\>X��UY�C+$� 齍[2�F`��IB���I�$�ݽ��;>
�=>f>ڂK�:Ӿp�?� ��Mؿ�җ�F�)��4?v�>��? $���x�:�B��N_?�*�>���`ֳ�s������?��?a�?��־��ż��>��>9�>94ٽ�ܛ�و���=>TC?���'���so�qR�>!��?�@���?��h��k
?:�t���w{�����|D�9>��8?�xW�>]��>�=6�u�*����u��L�>��?�?IT�>�Pe?Id��6��g�=09�>�-_?EG?�p<�o�7�m>\P?t��b򐿏~��2g?�5@c@	]?������ؿFr��x�֎���7�>� r>Ḣ>�9����=�{>�yX������="��>��>��>^��>�q�>���=YK��y������ӎ�o�*�Ŧ��x�Z������܉+�<�V��U.��>�ؽ�_��kf<�&��Dʽ,���S�=\�W?�nQ?��o?��?��]� �>1���܄�<n��1�]=A'|>�k7?b�D?�W'?H�s=�5����c��G~�����W ��k=�>it8>U?�>�H�>x�>�K�<�DJ>�BB>�}y>���=��N=�T��y�
;9�P>�g�>���>㔴>d�q>��=����Ʃ���e!���m���?�����_;�������+�̓�_^> �"?�ٯ=�e��ZsͿ���pI?Q��� a�`+=�G?�3�?!�=ge�-�B��՟=�@p���X��>�_&������:0��	�>�V?��f>yu>�3��d8���P�S|��(h|>26?�嶾�B9���u�q�H��bݾ�@M>Y¾>�]D� k�*���3�.ri�=�{=�v:?|�? 2��᰾�u��A��!UR>�1\>z>=�i�=:UM>oqc�S�ƽ�H��x.=9��=�^>�4	?NhD><)>�`�>�W�������v�>�D�>;�>�5L?��L?�96=\���gk۽�H��p�=��>�'�>��>>�S��縼�Zy>dҀ=�Ȥ<�E�q�6�Gq��郕>X'���ZJ�Ɠ�;+��SkG>U�#����4��_u>�j~?�����و�!a������D?G�?4{�=�`<W#���������[��?0�@U�?
�W��?�>�?.<��+��=�F�>e��>�̾t�M�_T?x�ýJ�����nm!��ԯ?��?C�/�D�����k��a>��%?��ҾX��>���c_��84���u�k�$=?��>�
H?����S�S��l>�(p
?7$?��񾕅��6�ȿ��v�oj�>A��?W۔?.�m�o ��8J@��B�>R��?5�Y?�fi>@�ھC[�C�>ƴ@?��Q?���>���	(���?��?EŅ?�TJ>�%�?Mt?	~�>��|�,.����������or=:�;^j�>���=�ｾn�E������_��\j�3l��\c>$=��>��F����	�=I����ͧ�Xh���>�ym>e�H>휞>J ?0R�>�!�>o� =X���3܀�3���y�K?���?����2n�eS�<_��=^�^��&?_I4?�d[�o�ϾRը>�\?F?�[?�c�>+��A>��&迿~����<Z�K>�3�>�H�>�#���GK>9�Ծ�4D�ip�>�ϗ>� ��q?ھ -��t��FB�>�e!?��>"Ү=,?-{?��>���>ГI�Gc���9���0?ޡ?J�?���?�i)?������|���ҹ.�o�u>}�o?��?�Z�=�E���i�_�>ñL�� ���0v?�~}?D=<�H%?�s�?HI?uep?��>.e�>�����d=kM>��!?Y���@��h&�E���?F�?�)�>�T����߽�)��ɳ��}���)?k�Z?&$?7��'+a�-���bT�<S�@�׋ѻ2Q�;����E�>��>'���Lɳ=8�>�<�=5Zf���5��"4<k��=+��>�8�=��5�����e�&?|�%=H�n�s>\�O�����m>A�Y>���# A?.���1��a�¿�r���Z^�ʫ�?��?eW�?�d�w�Z�� ?�ȍ?��?���>�)���6g���O�q+�������"=h��>���['�<��ϲ�!����4���y;n�?'�#?�V?/?�>��>r�f>2� �Bq?�] �=��D�l�*�۾
�3��F�/@0��G��e�/��+�=ᛦ��U���Pa>�z=��>A^?8�e>��>�j�>��/��Q>�E�>��>+�>�
2>�6>��=wE��$�=�2P?N2ؾ�y)�Uv�m�¾��I?��o?��>����_�� C�,�%?��?�ٛ?��W>�t��3�2Y?�b?��k�5H?�V=�b�=sԠ=
�ѾZ6�۬R��νf7�>	UP�cL>�Y�H���Z��>�F?1�=�r��j�˽r*���o�=�U�?�+?s)�tL��m�IQ���S���#�l!j��Τ�]�*p�������s(���&�$S=�3)?��?����h�-�����l��<��^^>Z��>e6�>��>!�Z>�
���2���Y��h!�^bz���>{?߯�>�xI?&<?�P?aOL?�:�>��>@¯�,��>�"�;�C�>t�>c�9?��-?��/??}H+?c>k�������\|ؾi�?/F?U?a�?�?�K���Ľ<��5l���y�(d���R�=���<��׽J�u�E�S=fS>Ҽ?��,�7��@��Ĉ>�s7?���>�S�>N�?���0���>���>��0>�4���4f�5���"w�>��?p����<%
>���=��_�<2r>5ʈ����=�a�<����!>;��>��=�&�W��<�?���=����f��>&+7?�s>���>�ϯ�Zz��{澺W`>S>6�[<Ne�=ɀ��8퓿}����_����n>�ւ?�%�?��>�0�=���4�������#����zs�=ig?��2?[�I?&�?1�B?Dv?��r>=������N�g��̧��	�>J!,?l��>0��ʳʾ~��3�Ϟ?[?�8a�B���:)�	�¾��Խ��>4]/��-~�����D�x�B��Np��i��?̿�?A���6��w辅���I]��Y�C?[$�>%Q�>w�>'�)���g��%��-;>���>)	R?���>=?�U?�|L?D��=ro�pT���i���X�=&E�=�j?��?��C?Y�y?�b?Md�jײ����}�z�.�q�TǤ<Z�A����<��>&��>}��>�J0>_l��%MF=}� �����j�=���;T�>�!�>��>I�=�e���G?���>=����cV���~����<�"u?�q�?�<)?� =�7��EF�~���|��>C��?!ӫ?��(?��L�!��=h*�,ȷ��q���>?|�>�h�>3��=��A=��>~�>S��>������O�7�L�5�+�?E=F?9��=\ƿ��q��!r�����p�<:!���1d�0ڗ�p�[�r>�=���L%��©���[�����d��O���A���')|����>��=��=���=�7�<��ʼ�O�<UN=�"�<�=Ҿq���l<�6�?�лKL���X��Z<��F=�����Ǿ;;~?��H?3�+?�+D?�e{>B]>��0���>xwp�cE?�M>���:W���<�$������Ohؾ#�վBpb�;L����>��c�F�>��1>��=*��<���=&}~=Z��=���o�=(|�=C�=��=r��=�>��>�6w?U�������4Q��Z罞�:?�8�>�{�=��ƾv@?��>>�2������zb��-?���?�T�?G�?Lti��d�>>��]㎽�q�=����=2>7��=��2�D��>��J>���K��m���~4�?��@��??�ዿ̢Ͽ"a/>G�9>�>�fR���1�ZX�	`��Y�]Q!?a�9��Pξ\̃>6�=���Ⱦ�+=�4>=�o=ݾ��3Z��G�=�	����0=/h=�ى>k�D>���=���O�=PO=t��=��S>1V4�7�5��.�y,F=�0�=��e><_#>�/�>�%?��6?�e?rO�>��9�yFžGx��q�N>���=͐>�S<�ڀ>��n>�?&0?6u4?E��>��=ɯ>�б>kZC���l�=L˾aϾ
)�=ڢ{?te�?��>�<WPŽK,�8�@�n��C.? �/?��?W��>�����ҿ��[�9����b�>>�>}�B>P��
�d�n��=�ą���w��r�<��8>Pt-?>1?�o>Fl�=��-�ܶ�>���=�=���=(���Q���C�㽹*�=b�c���L=Lv����=MM���E��Z�=t4c�� �.���r�at>d(?�z,>*.�>�N>�h���c8>����>N�Ѡ�=�?��irE���K�Ng�@�/�T�7�>
��>���Ə��?1��>��>Y�?wp?oR�=��Z����K��w�ݧ{���d=SD2>����V7���Q��jE��پ���>^ʩ>��>[$Y>�(��f'����=��羹�)����>啾���	ۣ�,=^����A����e�O�{=%�A?ӓ����]>H҃?=U?A��?g��>�0�yZ���L�<�����:|:� �w{�_���?S?�k�>(%ݾME�+�˾[����>�UH���O����� �0�8���˷���>󪾦�о� 3�6l��J��_B�or�&к> �O?ͮ?f�a��h���GO�ھ��숽ba?�Pg?V��>)?�:?���r��������=f�n?/��?/�?�>2�->Y{F<�h�>S;�>��?��?: Z?��Ƚ�`�>�yм�Y�=�;[���>�W⼕C�<�#�=>�?�G�>��?���%��O������1����9[O>e��>��>�~�>��i>PQ)>A��<3#�>��y>3��>�+>���>5)>�񢾀
��&?|	�=u��>�/?|	�>{=e��O.�<t!��5=�~�)�v���m����<��g�M�\=�Ǽ��>�9ǿ��?i2O>u��L]?q���8$��S[>[BZ>\���۪�>P�=>♃>�s�>��>K�>�C�>��%>(���>ݎ��&�[kM���R�S]߾��e>�����3�P���@��jN�n9���P�@`����qF�{}.��ڍ?�#F�$�e�$�>��
�-?
��>�*?%�U��h�OR�=%�>�>
f龻��LP����2Z�?A�?��l>.C�>ӰU?�?f�/��*��cR���`�:�=���f�5\�������x��	��>��EY?'m?5n;?V�o=��s>"�z?'t9�r���/�{>�?��/�>�=7&�>�,��>�M��䦾���6�:���;>��l?C�?G�?9�H�e�b�^c(>wt:?*�0?�0s?�0?Y);?U����$?�8>!h?a�
?�s4?��.?'
?�J2>ٔ�=`i(��!=��������ֽ�н�<���(=�8�=TN���:<�J"=���<P�׼��;�я��-�</^4=���=3��=�>�>�[?���>��v>�9?���6�5������1?�
<s
������8��������>�=Zb?_p�?PYP?�Q�>��<�&1J��>�΃>�d3>��`>Y�>\����I��{=�
>#�4>XR�=V@Y��V|�o��ga���� =��>�i�>��>���jG/>7����v�7X>\O\�j����K�4/E���/��f�{��>��I?��?m[�=Hv达̏��wc�˪,?��;?EnL?���?e$�=;�Ҿ_6�N�L�c��}:�>��3�����I���֡���9��]<�u>[�������؂>��[��#�j�[�3�)�:��b�=Q�����$�������X��=��=Ao(>{�f,�z��"����`?瞪=,"��\��<�/���=x�0>��i>�K��Ik/����ϘO���>�l�>��h>��Ǽz`��u\����
�>�D=?4�[?��?𣎾ރx��tD�����:��:A	�n ?뉻>G ?�m><;�=�������Kb�#C�cS�>`��>����F��H���<�R*�TX>���>FK>x	?��T?�*?@�d?�f5?�8?�"�>E� ��R��WQ&?٘}?2{=v.��&4��r6��VF����>�#?�"��̺>ɷ?�A?��3?��Q?�9 ?l�=U��+-����>��>ůT�Vz����>�S?�W�>�hQ? �^?�g>��4�X�þ�5 ��{]�Ѽ�=�(?x�?a�
?�ܝ>���>6;���=<~�>�^?��?Զl?l�&>��?NH�=�j�>r��=]A�>�:�>.?��W?�o?6�7?�?x��<|m��"�V�����<3�&=>��=�h�4ㅼ�<�:�;=��|=�����T�`<>�}���\<�����>tJx>����_3>Sþ�v��F�B>�h���;��ZჾG1����=p?r>��?�v�>�(�gg�=s��>\�>-�z0&?��?@?��&���`�{�Ѿ/%H����>z�A?=��=�p�uג���s��E"=&�l?�\?�ZM�����-[?�<?�\־m$�n澠]ľ|��3F?? �u��?�y�?<lK?��+?]#���U�����L�b�/u�qӶ=l-�>B���^����>�2?|Bw>�X��;�oʾ��o�`W���!?T�? E�?�K�?�F>�^��p�ֿ�.����^?�L�>�����#?UeϻOϾ�ԋ��̎��&��B�� ����픾[��m�$�҄�
4Խ���=Z�?Ɂs?J�p?��_?�� �F�c���]����xV����S�I�E�QBE��B�Yn� F���#O���H=��7��;���?°/?�t���?�؄�5F��5����P>,_���<Q�x^J>\���d���"Q=���~�3��yC��?�X�>#�>�J>?��y�9G3������yw��x>'.�>�j�>o�>9"�K�����0�u�VS���d���x>-c?��I?�Mn?����F�0��������3��-����F>��>/O�>�R��I��I&�d�=�Ayr����lQ��dv	��z=z�0?��y>�i�>m��?��?p	����%v�G"3���M<�ɵ>�?e?n��>z��>;ɽC� �p��>��l?D��>��>%����X!�t�{�6�ʽM�>ۭ>��>H�o>'�,��!\��j��;���
9��o�=V�h?#����`���>�R?PF�:9vH<{v�>H�v�G�!���򾬺'�w�>�?+��=x�;>��ž�'�Q�{��3��i�#?��?��(�-�'1�>G�#?���>���>g�??�>7���9��;��?.^?r�N?^�B?�N�>:~=�Խ�p��PO+�M�2=�Ju>�~P>0U�=�=�;��_\���sC/=�I�=�␼lN��dLX<�Cg�]�R<�	�<��2>տ��9�b��/�]Ҿ��{���H��勾�HL���ʾ� ��X����Q*� P=8n̽�6��vm�@-���!�?m;�?��'�M*ľM����h���:�4n�>ב$�4�d=ʍ��D��Y�p������]A�1�0��#u�l:p�;~'?}d��
�ǿi����mܾ,�?��?Kny?��T"��f8��� >���<	V���c뾁���NϿ嚾/�^?���>6�򣽝��>*o�>�HW>�xr>銇�*���,V�<p*?�-?M��>��r�u�ɿH���yͩ<��?� @�(??|�	������M�=��>���=(���'=%���]�핝>��?��c?�N�>&�9�W����?$)��3 �v)��;=�> ��={4���f[=I�>��,���нJ �� ��=�O)>��F��1��{L9�r4>d�s=��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=u6�󉤻{���&V�}��=[��>c�>,������O��I��U��=t/��ƿ_Z)�!�b�2=�gu��c�Nl���Ľ.�ǽޭ���Q�	O˽ag==�,)>�zx>�W~>Lq\>,qC>��`?B`q?�[�>0�=  �=��yzɾ>3=�P��[��b.z�_�,����WԾ�Lྂi��l�v�������S>�~��=x8K��ƒ�:N�9�[���W���,?��>�W����N��#0�dy��d���"z�8�p�m-¾i8� px�?�?�\@?;�y�a�:��V�����?�J?]����^���MH�=�$�<]��=A��>>�=��t�E�D e��0?��?<鼾q�i��>v����x<��,?���>���<�>�"?�^�鱇��J>²�=�E�>�,�>d��='����7	�"=?��??��_�����e	�>�א��_Q��{�=2�>+����7�++>��׽oc�1/�<� ��莖��V?���=C�	�"��>���-ȽY:>ߩ�?,3?�L�=Նc?>H,?OȽ�ŀ��ųe�B�о�=��?e=z?*�u>y���)����;A?�(�?�DY>"?��[�ž�iM��I(���?`�h?��>��=�D@��j����:�W?Su?�X�$���S�,�������q>���>
	�>��C�R�?E>?e�x���eT��/�9�*!�?L��?H��?;�B�����4�k>��:?��(?g@�������3����Ƚ���>VGr��w��A]�"���e?�z�?]�?]y��M�����=�������?��?�Z��s�~<\��V}k�ϱ���3�<ꋩ=1�������� 8�VRƾ�
��~��[�&�>�>@�ｉ��>�8�%⿢�ο�����ξ�q�^?���>�9ͽ����9�j�S�t�/zF��<H��ދ����>>����Z搾��{�Ʈ;��蝼J<�>93���q�>��N�2,��綠���S<dI�>V��>O��>}���<S��ja�?-�����Ϳ�S��D����W?R7�?&�?��?��><~Mt�3�{�����F?Ekr?BZ?i"��[[�I8��~j?ȫ�evt���W��,��t�>q�:?�%�>���yL==�=���>�>$�.������[�����>�?
չ?�i侓�?��?<<?�'�����b��3�R� Sl�Z?�~=w}%�^0�a���T���+�>��?��$�'�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?z'�>g�?�j�=Bf�>�d�=�����.�)q#>�)�=C�>��?��M?X@�>���=�8��/��XF��ER����C���>`�a?�|L?>Pb>�渽R�1��!��ͽ]L1�׎鼊p@��,���߽�5>��=>>��D��
Ӿ��,?߹0�`��F���HIe�=?�>xU�>���45`��hz��^?x��>�V4��󣿁��ݡs����?)Z�?��>Ozľ�ĉ�z���G��>oI>>+^~������d�>�$?��:��׏�R��9̧>��?�r�?W�?�Ǉ�-<	?�L��m��m�~�y��1<6���=q�7?�C��{>Jg�>�2�=�v�0۪��s�z2�>��?��?>��>�_l?�o�B�Ҡ7=Tݣ>U�j?�-?��g�Q?���D>��?��-���T����e?z�
@Bm@�-^?��ͺݿ�'����پ%�Ҿ�n�=u�=��->S>E�\��m5>6|=zO� �f>��>��>b��>���>6�c=>>�F����%�=a��UR���!��4$��#���+������v������U��ڨ��5b�2#��.C=T&��h�^�����=��U?1�Q?��o?{?�o�G- >�?��q�=�� �f��=4=�>��1?כL??+?7��=а��1d��%��ͦ��L���i�>�wH>��>-��>�Į>"�$;�I>G?>��>Fx�=a�%=��D�w=��O>h�>v��>�i�>�� >$iB>
�B���o����� �����?�����H��)������� �E=y�,?y�>����ؿ�ĸ�t�O?8@x�z�,�ɶ�=�r?�L?���='<���|�<G�4>�e���J����<�h��E,�Nex>�"&?��e>�v>��3��8�cQ�U���<)v>�5?|޶��j:�Wku�@FH���۾(9L>��>l:��/�?[�����
f���}=$�9?0t?�X��쟱�&7t��j��L^P>�^>-a=U�=�pK>>�p�ܱǽ��I��E'=�%�=��a>�
?�	>=�	>sr�>��ƾ I�����>[F�>Md�>�[?&5R?7�̽f*'�,m���u����>��>���>�EX=a��0�<O��>e�>B^�"��z�����u�>9����\f�g���$�=�0�ۘ��Wg�=e�h�a�޽���=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��L��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�0)#�jS�?��?��/�Zʋ�>l��6>�^%?��Ӿ�o�>�聾�q���i������w<��>#K?�!ξJϔ;Ճ��?�/?�l�zq��9�ǿ�<��eR?μ�?v,�?�R�� ���_��%?�z�?�X?[m}=���*g�;RU=�-?r�y?�xd>
���G����>���?b�z?�I>���?�s?�k�>�1x��Z/��6��Ŗ��-r=�c[;9e�>�X>i����fF��ד��h��'�j������a>j�$=�>VE�#4��=9�=�����H��Y�f�ϥ�>%-q>c�I>�V�>F� ?�a�>t��>z{=�o��ှm���m�K?�z�?�����m�5}�<=l�=^5`�Ѧ?�*4?i-K��1ξ��>3�\?��?t3[?��>���T_��}˿�����I�<K>��>�P�>�H����K>�vԾ7YC����>�h�>_T���{پ����Z�ջ~t�>�n!?.O�>鶮=�?!B�>��5>�8�>:d��2������j?�b�>c�>��?��?h��li������Ɍ�r�&�C�B>�7`?���>]�n;9Yp�ե��� �f���H��|r?5*p?�#���R?C�?X?�}v?E�^>@��_���g���&�=�"?����A��~#����Q?��?e�>A���ǘнOy���T���G�?>�Z?c!#?W����`�������<X�I������KE;���:�>��'>d�r�(h�=/�>t�=L�{��9���;�H�=���>$��=��/�f���}-?�����DPi�pAd���4��Ks>�x>��-#E?��[�su�IϿ&����Ɉ�l��?�C�?ݧ�?V㽲s\��$!?��?f�?�\�>W�h��^���Ǿ_���8x���7�#�>�_�>�p�{�۾hі�=g��U�|�-�==�^4��nA?r�)?�A=?I�K?-��>:>�(�ރi��'վ��P�v>��	���Xt �h�
�I���3�z�Y�~m~�7 �M�M���K>J�c��t>B�?.��>tU�>�!?c�>7�>��>��>]��>u�>GX>�?�<�e�=���]gR?�$���(�\�뾑���c�A?��d?%��>�)i��݄�*0�"#?s��?�'�?jm>��f���+���?X��>^���s?��j=�o�9��Q<� ��-��ʹ�*�Q��>�l�G�=�.PM���U��E?�L?��ϼ�'ƾ47�~N���rf=~j�?��-?��/���>�J6a�D�H�%
R��w��v�%������?h�[�����x�+'���X!��x�=��+?�?{��Ϳ�JQ����s�H�.�zk>�H�>���>�α>��j>���,�,�.yZ� ����#���>�t?a�>zUI?')<?�P?��L?�Y�>Nƪ>����8�>�@J<w��>��>��9?B;.?[1?l�?X�+?��b>�����I����׾E?��?G�?q?z?�����Ž����^��Px�X�{��"�=Æ�<:'Խ�?m�%mT=�RQ>ٺ?�('��!A����yGn>9?ԅ�>���>𡁾bs���_E=su�>�a? �_>ͪ���	b���k�>�у? �"����<>I>���=e���S������=�0q�Y=cA1�8/��e�~�d�=���=�Ǫ�ccU�tټ��=�I��� ?Y�?Т�>dc�>�ٍ����jY����=��U>�fQ>�a>4+Ҿ-ӊ�|���j�cp>:��?�ð?cE�=b��=�=�⭾�þ���
��־xi�<�?��*?��O?`=�?S??�??S>�������Ů��]���?#,?9��>&����ʾ騿�{3���??P?�3a�t��p7)���¾O�Խ��>'[/�*~�b��& D�{������Θ����?���?U#A���6��q�?Ƙ�l����C?r��>��>[��>��)���g��3�L;>C��>]�Q?�Q�>�E?6<-?��=?��mi��M���}]�5�Z>Ƶ)=r�c?��?�.Z?�?��??>���E��%����F���Po=�����2�=���>���>��>VTF>��P��$>�ڽb����˅=�p�=q�>Ov>�=>:�{>�=�H?ڥ�>���"�	��͠�I�u�ٕ��K�v?b�? ?R@q=���u�A�\?���
�>�V�?K¨?��"?��%�;�=&���8��xvu�8��>���>b�>X��=��k=�>f4�>`?�>k�����2��uL��I?�<C?�K�=��ſ��q� �o�Uw����_<֞���d�ft���[�ٗ�=O���N���e��b�[�޵���Y���>��ޗ��T&{�@��>�=�S�=���=5A�<�ʼḿ<�TK=*�<��="p�L�r<��8�3лo����G�uc<`�I=� �ѾmB�?�GI?9�.?OL?и�>tw0>�����>��J�`?D->�_B�f���p�#�b	���J��\ ž�߾��k�%+�����=G���9
>��!>jz�=��o=�U>�=�Ƥ=D<�=���=*A�=�E�=���=�:>d�>�6w?X�������4Q��Z罤�:?�8�>e{�=��ƾq@?��>>�2������yb��-?���?�T�?>�?@ti��d�>L���㎽�q�=J����=2>p��=x�2�S��>��J>���K��K����4�?��@��??�ዿТϿ6a/>`�9>�>�gR�̓0�:�\�hhd�h	]�_0!?<G:��X˾��>��=ܔ޾9�þ��5=�&3>�`=<�E�[�
њ=}\|�G�9=�i=��>d�B>mr�=s����|�=�P=1p�=�?K>`�ĻT�E�l�@�g)=�'�=��c>��$>J�>�:?��(?*a?t̒>�?i�W���I���$p>��>έ�>�ܒ=�g�=r?�>o?.??�9?��>���=��>�2�>�m7��U`�1��XѾ(��=�Q�?O��?Г�>&�=�-U�g5#�_1�R�R���?�5?�d
?�h>�������V�@�4�5[�=�v���8����}�g~�<0��qs콅,\=M�>8�>[�?�?ы->su�=4*>Ӡ�>�E>�	=�	�=�T<6�<k����=�J>iɔ�T轅�`=�
�"oT�׎��L2�����&>4)<��>���>�_�>a��>;q>g7x���>�pܾloy�+J*=�m ��k��o��t�1�+���,�Z��=�X>�Ed�<�����>7Դ>���>�|�?��i?�ED��!��4�߾a���VT��t�|��(F>��=�y��&�?�m��h�����O��>@^�>�֓>��R>��`��]`>k"�yYL�B��>��ž��r��C�1N�Z��M���!k��a�=Y�7?�⋿R�>1q�?* �?}[�?�ɫ>��}�=�z�|����S�T��ҟ�x�2��9?�T?���>����p<�[���5D���J�>���!A_����1/+��Y�=���5W�>�O�:���٘8�S��������M��W���F�>��G?�ߥ?����Pj�s�6��P&�b�*��#/?9��?�8�>	��>#�?��d�a��So���!��%F?���?Լ?���>Γ�;�ӻ=5v�>�"�>?��?c �?7(y?�D�I�>V=ݼ�=����lɁ>��=��>+}�>T:?5��>PA�>t�Ҽ�~�e�վ���m������<b.�=�Ű>�=>Bc{>F'>=��=q�(>{�0>�}�>���>��T><9c>�� >g�����!�*?r��=��>�;2?
��>�.j=��ɽO�=>�D��F��h!�u������ַ<F2��)G=���c��>T�Ŀa�?�Z>-�
�̞?�B�3.
���_>T�X>\ ̽+f�>�P>W�}>�k�>"�>`> ��> 
(>|��1�V>���ȋ��L�|�W����*?>[G��z�U���辸ۉ�*�B�՜߾��վ��Z�wB���N�����Ӌ?֓M�}�I��
�������>]��>�6?2�7�2��=u<�>��
?�܄=����뛿���!��Qģ?w��?��l>|��>�	\?�?��E�b�$�\OS��<m�
�@���_��_�r���|��e	�j��D[?߳q?-;=?5O=뵂>O�?k�2�*�S��>�^7��4�Wd=/��>�T����T��6ľ��Ծ�j���/>��g?Dԅ?�V?o�R�����wq�>�(#?�8?��?gf?w�]?2f���?��B>�������=ž<?Gg?�si?�;�>��>L�>�"���[�~���d���9�Rfս��3<���=8��8�{��T8>yѥ=�=<�Y�=�3>Ր=�
�=!�&>�ż!�=�8�>% \?���>��>��6?H
�+%4����Uz4?i �<��|��O��:l��%n��@>lk?!��?-U?�Q~>��;�0�E��>>e��>�,>�yh>���><!Խb�K�|��=�a>�#>0�=�Fz��]{����P���7f=�b>m	�>��|>vN/'>��Msy�Be>�OS�)����R���G��1�>v�e��>=K?&?�v�=3V辚K��s9f���)?��<?C�M?Z�?�=�BܾK:�lK�6��=�>�R�<�	�슢�&ۡ���:�8�:Vr>.���ɾ��>������o�n��aA�B��s�=Dn� X�=@���Cھ���m$!>Ely>���_��f������P?_%^=�����ٽt���KR>��>�c�>������"�Š(��T����=b�>��,>	�D��HG�c����>	DD?[�\?��?����s�7B�~���1О��Ҽx�?�/�>�M?�C>�|�=���T����c�t�D��:�>N��>�����G��ӝ�:'���#�>B?;>7g?��Q?��	?@]?�)?_�?/�>��0I��:&?�i�?� �=:Eҽ��T��9��F�:S�>t�)?eBA��q�>��?��?�R'?�YQ?�g?|�>�� ��?���>E�>D�W�M��$I`>3�J?�>��X?���?�6=>��5�c΢�}j��P��=� >�F2?�#?R:?�v�>�f?�u���n����z>�`?�m�?bic?N�{>r�?7=>���>Pg>�o�>Q�>p>?�i�?v�]?�)F?�?�<�x��F�=����f�T<�ߟ=�n<�>�=�F�aC㽸ٯ�uc,>6	�='�=��}=�N{����-AJ<;6x;�_�>�:r>����4x2>�5ž��
�=>�����ݙ��N����5�/��=��>�?l
�>��$�x�=�߻>���>F�� h'?_
?��?�L�;��a��ܾ�wM��@�>%A? ��=�l��c��'�t���n=�Zm?�X]?��U�u
��J�b?�G]?���;��qþ�4e�k��BO?&9?�F��'�>FL?�Yq?�S�>^�c��ln�O���D%b���i�1�='��>?���d�0!�>�6?��>�t\>���=lgܾ�w�R����?�%�?6�?:��?O�(>zn�C�߿�=�Ky��F*d?��>�Q��k#?7fV��ξA���΄�-Z쾨�Ѿ�����?���2���ZO�|2��i�M��-�=p�?P�j?�g^?zQi?�	���\���`�y�z�i2I�8���O
���:��o7�q�>��}f��T�5�߾�N����0=`$|��?E���?g�#?ľE�>$�>A_�����<�վ"}6>�L����Y��@=$�q�����B<��o�)&�U�� ?�5�>ޕ�>�D?�l^�g<�V�3�E�3�9�꾆�>8�>6F�>�>�}�[�>��ƽ�Ϲ�U���qF½dru>O�P?��8?�Gh?0cF�3�0�����7b(�3�VS��t5>���=|el>�?�#���� ���:��n�8N�����w4�+��=@4?U	�>�>�>�?���>?-��������M�x����Z>s8P? ��>�>A>!�5� �ΰ�>Ɯl?�/�>C%�>Y`���|#�Low�+׮�4��>�e�>�F�>��w>uE.��}[�􊏿4^��[�6��@�=I�h?D4��(�d��܄>�Q?ض�D��;`0�>�"E�G[�\����PP>�	?��=�;>Ȫľ��
�b�x�5H����)?�?����}�)�K,>��!?���>y��>$*�?��>�����n�;��?�+^?E�I?n�A?f$�>7V =���Ƚ��&�N#=M�>`OZ>�m=/��=6��bA]�)� �7?=��=�y���۷��8<׾��e/<��<[�1>/꿺�7� �Ծ�,&������l��������H�A띾w�<�[��-~���!��Y���E3=�2�G�0���r�^x���?:g�?��_�k��$��ےp�ޔ����>�]��	�G���@X3�)S꽏'̾&n�����1K�l�~�d����'?�����ǿ𳡿gbܾ�. ?�H ?xwy?���Ș"��8��!>�Y�<5&�����+����Ͽ5T���
_?���>��飽��>���>42Y>��q>���3����<��?a�-?�r�>}�q�Auɿ�t���-�<��?i�@\lA?��(����$Y=F �>��?e�>>�0����$��Ȱ�>V.�?���?e2U=*�W�[�FEe?���;�F��>ػ�j�=���=1.=��\NJ>Fr�>(_�ףA���ݽ{�2>���>+i!��%���\�Qȹ<�]>H�ֽ�ɕ�5Մ?,{\��f���/��T���T>��T?�*�>D:�=��,?S7H�^}Ͽ
�\��*a?�0�?���?)�(?,ۿ��ؚ>��ܾ��M?fD6?���>�d&��t���=7�E�������&V�b��=P��>^�>��,�܋���O�J��;��=����ƿ��$�]}��Y=:�ݺb�[�G|�k���9�T�%#��4go�m��T�h=ٞ�=��Q>Hl�>�%W>�2Z>9hW?�k?�N�>|>IH佚���ξ�I�G�����ͦ��.���ꣾwR��߾_�	�	����D�ɾK�Q���!>V�I�]����Q.��U���C�#0?��=3�{�l�@�*�6�R{���F���t�=��U���nH;��I���}�? /R?�h��6+L��}���iZ�S?�!�[���{���=D��=�c�=�޴>��=��ܾXD���p��N1?q?�o׾.�~�	>��$k�=A�*?��?H"=�A�>��4?�����#���>�$v>1ҙ>l<�>\�P>���Ǫ��u ?�VA?PA��E����T>J��鋄���=�K>b���Q%��Р>�D=EӾu"C���+�@���{O?� �>U���]�e*���zٽ��{<�Ā?>V?���>�?�SQ?LE��x�u�r�@�le��==(FG?A^?'i">w(�1���HB��Vr5?�U]?!1> ����O�"�@#�9?{u?|��>˵=�n���ꄿ�a���*?:kz?^�l�`���+���Ua��>�� ?�!�>�h+��'?��A?@X�E����r���-0����?q�@n,�?P��<kl��{>�M#?�?>+i��������i��{����?�耾��n�� ��ͽS�+?}��?�V?���ӱ�j��=V������?�9�?����b��<���z�i��I��u<>uG=�:ɽX�{�9�徦�=�:;��� ���ʼ1R�>�@0#��r�>��L��B��ǿ���Ǿd1{�3�?�+�>��ܽ������e���e���:���K�����2֦>�Z�=��#��nq��u�I�B�.����8�>aNm��zv>N��A�Ⱦ� ��/\�<ŝV>0b�>�k�>��U��vվ�z�?���Sȿ&���NZ/��7?|ҝ?���?_�B?�C>͜�-�,�����JkC?�)?͕[?��=�~�����o+m?jǾ<�l�~?��f>�.L[>�b6?���>,�(���==� >�>*+>��)�����L���gվk��?ó�?a�ݾ�r�>W�?,�/?�!�M0��Xr���ؼ�&\?Xd>�(ھ��'�X�3�`�&4?�H?�����%�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?~��>�>?��=\'�>(~�=�׿�����d
>Q>��D�@�?�R?�;�>dL>����"1���?���R����NQ@��ׁ>�9Y?�GA?�|>[S������e�'��]$���G�Q�B���d��H����2X>�N>&^�=�D��4߾�.?�V��nֿv����xg��iY?Gc�>��>UӤ�$��l����m?[H�>@�Ծ�G��9��������?"��?=��>����b�Z�>j-�>��v���7�	�;ű�����>՛Q?"��L闿;$V�xL>�V�?]T@��?nP|�&	?�=�^��t~��x�E�6�`��=��7?]%���z>c��>jƪ=Rv����}�s�dj�>�?�?�|�?���>��l?�Xo�"�B�9z3=&<�>dBk?�P?��Z�^
�
D>n�?��e���{=�f?��
@�z@x^?���ڿZO���y����Ǿ�]�=cj�=Ն>���s
=
7�=�E���b�9F>P�>Hb�>���>�.c>�1:>�<�=�����"���������D�;v��� ��=������K����0����д�酸�G�?��¢��I��&�n���]z<M�e?uqY?h�x?'�?^sH=L��=���T=C�S���<��/>0Q.?&0?��9?��{=����eO�e�x��þ^�����>hOO>���>��>�ӳ>�CW=.�l>�}>���>��>˽�=��=�̛=�Ja>)��>	�?��>@�
=�i{>�ϫ�=<���N^��:y���ž��?�׾�07���|������5�u��=un>?��8>�T&Կ����I\?��a�	�=��=E>��??�5�=�ш�)�v�d&[>F);R:� ���ZJ�eU���	8���>T�?�e>ˣu>I�3���8�A�P�����z>�6?��9� �u�u�H��ݾ�aM>��>�;��2�����F��*h�iy=�:?��?:]���s��'iv��:����Q>;'[>��=7�=nM>1ce���ƽH���*=���=�^>���>E�,=hy�=��>�����^�Mڈ>�++?]�	?��.?A�t?5`�>M
Y�`uq>��Ǿ��=sv�>�N>z>l����7�k�>t%?>���=Sb1=H0��`Y�n�>�܎�b#��%��<�����R>� �>�\?=H�Fͅ�[��~?+���1爿�a�����D?0L?�u�=�
N<Z�"������ĸ���?��@�T�?.�	���V��?�P�?���G�=�o�>���>c�;�L��?�ƽ������	���"�9I�?�?�'.������ l���>Ä%?j�ӾƱ�>�پr�������1~���^=�g�>S�"?͇������n��x?YlA?U� �n2����˿�r�����>3��?�*?�y`�믎�6�b�D�>�4�?o�?��<��r�����)���;?�d�?*(�>�Q۾���D.�>�<�?���?�I>d��?��s?�v�>��x�6b/�g(��i���T�=��R;IW�>��>����mgF�.Փ�b��n�j������a>�$=��>���2��4�=�u���(��?�e�>��>�q>*�I>2i�>�� ?�[�>[��>,�=�T��vۀ�J���>�K?.��?�� n��#�<9��=�W_��?a@4?�\���Ͼ��>�\?-À? [?O1�>h��~;��;ۿ�S���g7�<b�K>� �>���>����-�J>zվ%E�lB�>5��>𔩼�9ھj_�������_�>�=!?S�>jޭ=��?Oc&?��K>Ƚ>L�E��W����4�=$�>U��>7g?עm?R�?��Ⱦ��:�@W���噿Q�N�Ӛ9>��o?�?+��>蘿��S���3D��A���W�cP�?;Xk?�S½aC?u��?]|9?�s;?�X]>
�>�ž!윽� �>�J"?���P�A��d&�:����?��?��>�z��|�Ͻ���K�������?6Y?�!%?�<���a��>��ue�<)��=O���8<����� >�>Bǈ�ϳ=��>�Ʃ=Ǵk���,��<6<�V�=T�>/��=*$.�\E���/?S�Ƚ�U�Xv�=,�X��}-���>�"�=/�
�Y�`?���v�t��/�������ȉ�L�?�/�?�?�d	���`���0?n��?�I?��>v?(�F���V־�	��K�þ�3/�<�=v�^>l�Խ!߾�����X��[Bk�JԽ�r2�c�?
?�`?�(&?3E�>L)�>��KXM�"�(��^F�;�V�g%T�����	�/Oþb�� �-C����I�۬>���=�v#>���>�&�=���>�{?�B�<Z0�>^K>��>ᩔ>��/>a?=�B5=�=�2���oR?Sܾ�F-��� �Թ�y�K?�'k?<��>s�f��߅�����n,?�ט?㕙?��Z>@n��:���?��?�w���?�<=�6��H�=������o����s�`>Ź�3h/���M��B���?��
?�b�<?���G���ъ��wn=�f~?��5?�&1�\�B�^�Z��F�PQ�.ɰ�2���`l��G�)��o�,����u�A�l��"�I=�#?�ɖ?-���Ӿ� ��邁�!j�V��>N��>q�_>?��>�8�>̤�D�@���G�_��/hI����>ei?
Ar>AN?�0A?��S?�5T?Ҽ�>�ۤ>U��6�>?�E���>���>��9?Ņ)?�p5?OB?�a*?��p>O����5u־�?��?ݐ?.[?��?)	l�:��F����AC��^�c~�,�=���<��+bF�yLg=�a>�?n&��L:�N���B\>�*:?F�>h��>��ȅ��+Y<���>�?o�>�, �(�s�/��b��>�r�?/���:�<��)>��=K�&���<�s�=C˼I��=���*��<&��=�g�=G%;�Ⱦ��$f<3#�<��<t.�>2$?��d>���>���PZ���>�R>��>��>-���lB��V��EAm��a>ɇ?&.�?�=&��=�1>������� ��K۾�O�=��?�.?ʺK?*�?�E?}�"?��'>
��g-��u������~?p!,?늑>�����ʾ�񨿲�3�ӝ?Y[?K<a����p;)���¾R�Խ�>�[/�$/~�����D��ⅻ����~��+��?ۿ�?A�N�6�y�ܿ��\��C�C?�!�>KX�>I�>�)�K�g��%�41;>Ǌ�>"R?���>��@?��g?4�U?�?>Lf?�ǋ���Ē�]�3=�>�}=??��?O�?(?�?b�>(��="��������o�����ps~�ErC<͎u>kE�>ʯ�>�bZ>��J��w�罭k�#E|=�> l�>��>戰>��R>�h@��K?�h�>��&��꡾�����<gjJ?��?�^7?p��=nz
�qsR�J��ϥ(>���?��?��?���y*>
;`ȾA��T��>0�>{�>QA>](�=��>).�>�u�>*��H�R��|�>j��>�/?9�X>�¿!br�UY�����u��;8:��g_�ɯ��H�c�r��=�;���+�����7U�����Yt���ᶾ�+���x��U�>���=�/�=<��=���;=Jۼ��+;4�=ev�<oS�<Tb]��x+<�]&�R�$�e֕��I�?<]h=��컳ھ��?8O?�J0?YvK?��>�&>�a��̚>���n?��F>i�������7��q���Ͼ�4Ӿf�r�`����j>�\��>�`6>�? >WI=��=�Cq=W�=B�I<��&=��=K��=_i�=z;�=K>9>�6w?X�������4Q��Z罠�:?�8�>i{�=��ƾw@?��>>�2������vb��-?���?�T�?A�?<ti��d�>C��N㎽�q�=I����=2>u��=x�2�I��>��J>���K��K����4�?��@��??�ዿ͢Ͽ,a/>v�z>4�=�N��s1��e��@���<3���?0-������U>�6�=���+۾�a��V�>v�>������@���=Y���h��1�*=&£>�I�>YS�=ج佋 �=
j/=���<ņJ>�S�=yݽ�[=jP�=�@�=���>�?�>��>�??J�,?"�f?���>�"��aԾ3̶�K
>%ʩ;8I�>�2��˚�=ge�>c�+?)�-?��1?E��>�<C���>R�e>ec&���x�ڒ*�'�þ?>��?�!�?��>=' >u�	�#��PI"��?1�:?��?�>�U����9Y&���.�$����y4��+=�mr��QU�L���Hm�2�㽱�=�p�>���>��>9Ty>�9>��N>��>��>�6�<zp�=$ጻ���<� �����=$�����<�vżė���u&�:�+�2�����;q��;@�]<]��;9��=<}�>'�[>���>p76>�$��B�%>X^���]�.b+�c4˾�^�r�P�6�k�?����^��>�Z>>5u��D�����?y�>D�>���?&d?��=\�� �	�����ؾ�<��q�|�g�۽� ��>�k�h���_�Gľ���>Wَ>�>;�l>�,��$?��9w=V⾏Q5����>s_��%v�{#�� q�5��W�Fi��Oֺ5�D?�B��k��=� ~?t�I?�?<��>�t����ؾ�/>�S����=+�*[q�Yn��u�?�'?&u�>��~�D���Ⱦje��<��>��>���N�s[��&>/�����^��I`�>�����ҾFm3�����!��
A���q���>--L?xǭ?�Gb��}���:Q��T�?���n�?Xch?Uߨ>��?�?������gy����=��n?���?�E�?�|>Q]��d��>��D?P?�V�?]�?��^?]�s����>y[�i�@��t	�l"I>B;�=���>�?�>@�"?���>��>P%�D���K�������������~�>藤>|�l>QG~>UP(=��=Ɓ�<-x4>�8Q>^�>.�>�֝=Ehp>�x�����`B+?�y�=H��>11?���>��D=�(��u�=Y���:AM���#������/Ͻ+ �<TV <�g�=`�μ[(�>؂ÿ��?�7:>u����?�����v=�RS>��_>ńȽ5:�>9�:>Z]�>���>*ݚ>A>dք>��>Q���<��<�e��-����F�#�V���;��ˏ>u��ٖ����6f�=�l&�l	Ӿ�����Dh�M����-�Z��l��?=�׾e�>�!����c����>{�?�?���ڻ��/>�>�>� 	>�n�e���H�����X��?b`@b>���>$�W?�?(4��03���Y�˰t�֕A���d��`�H����m���
���ʽ�]?bw?b�??��<|P{>( �?h'�j������>��0�J�8�y�W=���>p���\�#�;��þ��~�A>;�n?ᕃ?J?_�R�����᧕>�.W?��#?'�?��C?&�+?"'O���)?� _>��>v�>�b/?��2?�+?��>�׊>N�P���<�Fj�3 ���ֽ#Fx��K\��1�<�.��_㛼�AB<�Y>>��R�'CD��k;�-��=30��rK�<���=���=�
�=0�>u�]?�6�>!��>��8?o��{�7�S2���/?v>=Q���抾ue��V��m�>F0k?۫?`�Y?R�b>�kA���C�^�>��>�%>��[>6��>G���D�{��=2>�A>q)�=!jE�:I�����r��ْ�<��>���>�7�>
���c>�C��T����=���h���HDC�eu#�&S!�w���%�>�mH?��	?vá<�!���ν��j���6?��Y?��S?=��?՝�=�,Ѿ;�V����ޱ���8�=P���f�R4���犿�-O�l2����=>L���B�����d>��Y߾��m�C�I��d�N�@=�G��E=^��	]Ѿ2�w�i��=p�>z��i�!�藿߫�,�K?�т=��FW�����g�>Sa�>��>��H�rZx���=������=#�>��6>���ԘF�O��G�>�SE?�I_?o�?�悾?�r���B����N@���	ʼ��?^7�>oA?F
B>>�=ː�����1�d�!�F����>KQ�>�����G��^��"����$���>�?>�>��?Q�R?��
?�{`?�)?.P?�/�>+)��M0���U&?�H�?Ge�=�ս�T���8��3E�2��>��)?�x@��-�>*�?�?�'?u�P?�!?��>�% �s�?�ꈕ>@�>��W��;����_>$EK?��>�wW?�ă?4wA>_�5����h4��{s�=�c!>(*2?��"?,�?�ٸ>ʥ?�Γ��Ea;��_>�O?}��?��z?F���br"?䌱>���>���<�>�? �?�hQ?��l?��g?���>�<��ҽ-���ɲ���k=&�=�e�<y �=��o���轟�V�8�Z=2H�=)쫽h~�<�X�������KV=���>�d>a���3>����zy�$v9>98=�֍��w���齦7>3�{>��>^�>j�
���=G��>+�>� �C�9?�c�>�$%?���=��Z�y}�^.���)�>+5!?w�G���o�d��:�q���>9�K?�KT?������J�b?��]?h��=��þ��b����|�O?D�
?��G�0�>��~?O�q?h��>-�e�:n����Cb���j�Ѷ=�r�>OX�6�d��?�>s�7?N�>��b>Y%�=hu۾/�w��q��\?r�?"�?���?.+*>|�n�C4࿴yھ1≿?
Q?}��>�����K ?\ӣ�j�ɾ[蝾l���DؾWzz��#��m]���Z��f������ݽM�=-:�>q�|?�!{?��j?��߾Khf���k�f����C[�� �����Z��R�$�;�x[�64��s�e�ƾk�,<D�v�.�@��@�?{)?�7:���>=���b��zվ_g>>`6��NJ�i8�=����r�=�m=�f��t+�G���?��>���>w'=?![\�ە;�7�-�j�5�GB��j�>�6�>�ӓ>"��>�j<>�-�D��!ɾ�ń�K�ɽGy>��c?��I?Ip?�<���0�Ԋ��c@����p����:>���=��>�rR�?���$��:��tr�h��k��������n=$�,?��j>�ٗ>��?�?S�	�1���b�x0��d�<��>�%a?Z��>㌇>�Խ�F$�}��>*�l?��>2�>-����T!�^�{��ʽL�>��>��>ʢo>B�,��\��^��|����8�6�=��h?����~�`��݅>�R?-�n:�)H<d�>�v�ӱ!������'���>At?#�=�|;>Tvž1���{�&���t0?���>�+��.G���>�C?��?��r=�:�?�z?lC��~?xfo?�&?X�J?]r�>�/�>��=k����>����:��6>��>r�>4F�=A'�<Ka��_����'=�]>}Q>Pw�<�=����~��o����->�9׿�
V�w鳾�4Ǿ9�������ξ�;]���q��ڽ���Q���G�+�@�C��;��$���V����_����[�?�W�?�kf�X��;錿�o����{�>��ȽŐ8�^���Fɽ�q�����xuy��N���;��偿�%d���'?O;��W ȿ�������r_$?�M$?[or?���"%�[�>��J>MM�=��������i��(�ҿ𛖾o�g?��>p+�{Ĕ��u�>�>�>�Gp>�4>���+���3ﺆ�?�/?2�>�EL���Ŀdc�����<k��?�;@l�A?�e'�:��}]&=�R�>W�?�J>�'�;Q��g��8d�>Į�?�$�?6GF=4�T�&���Xa?VV�<�BB���7�L�=_��=9I=�����?>M^�>B����V�d���>�&>�ԋ>,�)�ET��	V��C^<\	T>]�+Т�5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=s6�����{���&V�}��=[��>c�>,������O��I��U��=>�8	ɿ
��s������<��<����R6�0*I��o����{�k��{��q=s1>��%>>�I>9�h>^s%>p�d?��_?'��>n�S>��+X��]ھ�=d��z8߽�8��7�`��\���<��u��*J��4��Y�0þ��?�:��=�7��
|���'�"�Q���}���>BC>����]����=P���X����>d�<H��@Kj������Q�?�m?��9pg����H!���N?L ��~�;n�Wm�>m�(��,�=��>A�@=������F�M^��F0?��?%�߾zn���=�-����=��*?��?s!>�Ŀ>�u%?'�� &��s+>8�<�q�>g��>�:/>Aۯ���;?iY?ڱ�`���Kj3>�W�������.> {�=��3���z=vʶ>�m�=�2�J�l�U��Ȓ�<}RV?ҡz>�+�����~�oQ�ږ>mk?�?�Ұ>~j?�D?�;�_¾+�H��QǾx�=�O? �b?�>��<�_ Ѿ�Ŗ�>)?�[d?J�C>=#����ݾb���+�B4?�yk?x?� �=��q�@����;�o2?1�s?��Y�fl��������{S>��>�l?�04��l�>�S;?�������`Ź�&-+�h'�?̬�?$��?U���WѺ����=}�"?&E?�<���L�/�7�]qɾ2�U�n��>�{���ˍ�ʛC�Ur@��S?`�~?��?qyǾ�(����=�ʕ��S�?��?�x����d<s����k�;D���<e�=z����"����/�7���ƾI�
������"�����>�W@����:�>R�7�8!��UϿ���GGо>�q�d�?sj�>��Ƚް����j��Fu�2�G���H��v��t1�>��>�����|��*p���<�<!+���>��׻�>E�'`¾�Ϋ��P�<��>��>G2�>��Ož���?&���`ƿ�f���S���L?_)�?8��?m�?��l=���k�j�����$"<?F�S?�Va?s!�HU����8�j?�9���g�51B�F�9�
q>�0?��>R����m=�%>д
?a	>��4��K��B���%�zP�?g��?�!�� ?w^�?��0?���פ�>���C�!�5�Q�gfO?v�i>�%���$8�T=@��	����?Y{F?�|⽋�1�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>iH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?n?�>��?o�=ޫ�>g��=�����0=���#>b|�=�->��?M?���>p��=dp8��/��F�.0R�>���C�l�>�a?yL?�
c>7︽*�7�.!�w`ν�2�:1��;A�;�.���ཞ�5>V�=>>^jE�%�Ҿy)?*;J��|տ8��o�c��A^?��>��>A�Ͼ�� ;�>^�?�_?zK�pͨ�4��F�޾{��?>��?��>�#2�lf7;I�W>a�?�N�=UZW���1>�e�P�>�o?1O�T��ѝe�'��>�L�?�3@���?��x��y	?�R��p��V�~��u�3�ߍ�=2/8? ��g�y>���>L�=�yu�������r�y1�>c��?��?�%�>1�k?��m��A��:@=� �>��g?I�	?��s�Ґ��H>EQ	?49�9���P���me?q�
@�t@	^?Q����߿���gպ��A�=���=�D>'*7��!l;D�<2�`�x�r<�>�ɴ>�ƍ>�KX>��?>>l>�4�=֞��,��뗟��O��А@���/���a{�Kk���b��z�k����y��U�����{�}���2L�����O�?����?*�?��?�e?�!�>�.7=�'�>� ���վ��)� �>�L?��%?)�H?��*>�^��9�]�L�I�/���9V�x��>8��=t#�>���>(+�>��>Y�>�>`��>��R>
��=c�>���=���>�J�>}?qT�>��>�G>�t������Q�^�%����Nf�&;�?e唾��F�2ԑ�;9A��ў��2�=>L1?D�>
_���Կ���o�T?��k� �x-
�M;>�?�E?�+ >*´�
��$g?>��G���Li= lP�Mɔ��&��`>�� ?��f><u>P�3��d8�1�P��~��	g|>46?�趾�?9���u�вH�5eݾ�GM>J¾>�8D�Yj�������5vi���{=px:?��?I8���᰾=�u��A��6LR>�8\>�X=^g�=XM>�ec���ƽ�H��a.=ɹ�=w�^>��?�`���=���>{��e���U>9�??���>J|U?P~?��;�:}��3
>����`�B�Ƥ�>�($>��>��6����=�?��>��=��T=�2���h��T��=��b������<�=B*�=�S�<g��=�$�>�"ҽ2��x�x=�~?���'䈿��
e���lD?U+?^ �=��F<��"�C ���H��G�?q�@m�?��	��V�B�?�@�?��A��=}�>׫>�ξ�L��?��Ž@Ǣ�͔	�0)#�kS�?��?��/�Xʋ�<l�w6>�^%?��Ӿ���>s̾�b��C��.��q��<S�>վ#?�Ї�ux�o���U
1?~�?O0��E��-Ϳ`��ZhH>��?��{?v%��oS���Xo� t�>���?���?�ݴ����s��"���Q�8?�t?�4�>+�̾�V��*qj=��?�n�?�;I>���?��s?���>�Hv�oY/��=��ـ���t�=E�S;=5�>a
>���PIF�l���J]����j�����*b>��#=� �>�k�`-��yյ=����I��V#g�	d�>��p>�sI>[�>"� ?�-�>�}�>�=�A��򀾽Ζ���K?���?,���2n�O�<R��=/�^��&?�I4?k[�z�Ͼ�ը>�\?j?�[?d�>;��O>��E迿7~����<��K>*4�>�H�>�$���FK>��Ծ�4D�_p�>�ϗ>�����?ھ�,���R��EB�>�e!?���>�Ү=�� ?[u#?p�i>x��>ybE��5���E�K��>���>hU?��~?��?�#��R73������ۡ��>[��&N>��x?f!?i��>�l���K��`�B��DH����1t�?�qg?X����?6�?e�??}�A?�6g>U��L�׾ ���,&�>��!?�,��A��&�4V�/?2?�?�>ܐ��kӽk�ɼ���ۺ����?մ[?�&?C�'a�$�¾���<oN*�[P�q��;3�G���>��>�W���b�=��>zܰ=uel��L6�oDk<۟�=�̒>�K�=N�6�t`��g�/?�����aD�{Ǹ��Fc�SD��a5>�@g>��)�Ź>?��*�ܸ~��ͮ�z����s���d�?EI�?��?��Z+T��?Ob�?	S3?�>gl{�E���ʾ���ZmB�����=��?�	����@߁��=��Dt����=p���x�?Vc?+�(?z� ?C�>
8>�����Q��C+���)�l+e�r|��9G�� �=	���ؾ�;��A��;�E���2�D<n>�">�xz>e�>�@>�~>�A�>��%����>�_�>�r�>6�>Λ>]�*>�Ĥ=�:���ؽ0�R?ſ�.�&�����ª��C?�&d?�w�>�����&�����&)&?���?�+�?v>�b��J+�m\?` �>8����P?S�m=�\�<=��<���_~-�L���P̆�Vƃ>MV�ҽ8���N��o���?�}
?�l��H4ؾ�F��������n=�M�??�(?��)���Q�;�o�ҶW� S���d8h�ki��@�$�ěp��쏿�]���$��Y�(��*=��*?��?[��E���"��q&k��?��bf>��>��>�>�tI>S�	�X�1��^�,L'�÷���Q�>BZ{?@��=�bj?a�V?S�`?��?8�>�>Vו����>vƼV�/>���>�<?KS7?|�J?� ?)�?��2>kt�W��ff̾�.?Ă?x��>���>��?K�2��d��^;M��<�������j�=Û.=��筻�<��>?F�(/:�p���v�=�:�>#6�>�2�>�J�T_�<��+>�Ώ>��>o��>";羧����bپF��>
/�?0��73���(>$��={Y:7�p��]Z=S!�<���=~H����� $�l�a=
��=������"=����ݼjf=�?
�?5�g==Vk>i]�����]��G(>O;%>�d}=�=>����"��������^�5�>���?@x�?bq#��0=<!=آ��3�6&�-���k2��� ?��Q?�h?��?Y�-?OG ?��>n����-��tY����վ�p?v!,?ℑ>j��=�ʾe���3�+�?�\?�<a�\��68)���¾H�Խ��>�\/��)~�����D��脻�������ݛ�?$��?�MA�D�6��s�弘��\���C?�>�X�>e�>�)���g��#�n;>9��>�
R?�*�>.�O?k,{?6�[?ښT>�8�,5������/�s�!>@?}��?Cێ?y?9s�>.�>{)��"�����,���₾ZV=]�Y>-|�>��>ש>�Q�=S-Ƚ�e��2+?�V/�=�Xb>?i�>X��>��>�Iw>+�<��D?@۬>�u��a@��H��*�����=�8`?�3�?>12?[��>���e�R�����>Xʤ?̷�?��
?�j~���>z
׽�lϾ�ľ	{>6��>Ƭ�>��M�>y��>P�>���>������}����<*��>��T?��>��Ϳ���� a+�>7�J�ټ��}���S�cu�zʅ���=�ʲ�.�1���y�3�Y�&9q�W��y&Ⱦy��������?J~�=?��=-J�=æa��켧��(	�͆�=eCc=YfL�x���06�=�B��/������<�"=W�<�/�q[ľx~}?�F?��.?I�D?�cl>�H�=98�+�>�����r?ϚI>�'��).��]v.��ħ��J���gھ��̾��f��ޜ�,� >��V���	>e�,>	��=B3<�t�=�CM= Hp=/���S=���=@�=@��=�H�=>>�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=J����=2>r��=x�2�T��>��J>���K��B����4�?��@��??�ዿТϿ6a/>�XD>#�=�N�{9/���`��_v���R�Q�"?.:�Xž�l�>���=��6nȾ��<�I>�0�=���[����=��`��TV=�bm=���>�P>���=bd½zĭ=b�3=�L�=Ci[>#�*:fK�f?���f=��=E�_>��<>�E�>\?�((?��g?���>�
������ɗ>Ƀ�=D�>B�<\�=�ٵ>��,?�8?�%K?ת�>��=u�>�_>��%��s�M5�K���?9�=�Z�?�*r?mY�>H��=E�M��~���7��?�f�?��-?}f�>�"9>�5����S[%����&ڶ�P�:sӛ=	���Dn������#�V<�W�=�R�>��>Aw>��C>��}>PC>��>"��=��=5>z�<9C|=�FI<�X�=O6v��V��/���m��M+����`������jּ��=���<��>��?�|�>e��>�]>7����< wо�mP���P�̗���[J�0_`���j�y���Dn>�@��=ĸ<�����0��z�+?���>���>���?�be?���;I���^Ҿ���T�ᾢ�Ѿ$b��L=����?8�WT�ĞZ�Z�����>@�>�>�hn>��)���=��Zm=����5�_�>h���v��v��w�o�/᣿{О��g�24���B?�s�����=>a~?/�J?B�?k�>2R��ڹ޾�*>3H��췶<G���y�5����?�|$?_��>=�ﾌC�0�˾{$���)�>gG��P������F0�>�qW���İ>.Ϊ�b�о��2�pS�������B��q�˯�>�O?ᴮ?�*a��|���%O�@���r����?g?�e�>��?�h?J����O�<U���=�==�n?���?<�?%	>�G�����=k?,��>�ݘ?�O�?�t?�Α� y�>�o�$*{=H���x5>�2>�ɇ>��U>��?g?-�>��X�ӷ�D���L2�l�0�'���$��5 @>���>7��>pd�=���'A=*��>�.�>��=�73>�L�>'R>>@���p	�2[(?���=tF�>8.2?�>�E=�6��a��<*]���D���#�~Q����Խ~��<ާ��$\=�WӼ���>�xƿon�?"K>���V?H�����-�;Z>Y�X>��ֽ��>"hI>��>4�>���>��>��>��(>˰��`�;>��6�Z��pH:�$rq�A�j�W> �;���ý��۾��>�G���߾{[
���|�s}�Ӛ]�����?F^�;�G�����v��lt�>$��>�hB?Z���|ֽv�M>'��>)u>Z���ۺ�K>���.���ڇ?���?�-�>�9�>}�A?�n,?b#���6�'���YG���R���i���?��<~�b�}�9���M��f?�.{?��<?�=�[>�z? `o����E6�>�NN�<
$��́�^��>	������?��B�&�����a!�>8i?�a�?�**?yUȾ� ���μ>(�f?���>�}?;%?�06?�U��&6�>�%A>(t�>O>��6?,,??{O?��>��X>��W={TU���̽튾��2�MH ��)4���}�;;��r�738<��=o�}=��I������	=-��<`�8=��=��5>�><�W�>5�^?B4�>뷒>��:?�;)���>�����Գ2?���=��rG���ȭ��$˾(+6>h�Y?��?�xL?}V>KtK��$8�5��=^�>�>�iP>�~�>̇���b�=�\=H�=ƍ�=�څ=�3�
��F�҆��S<Ű�=j�>Ú�>Q1g�6�1>�V��hl�H�G>�_��-þ��Y���A�I�(�ܷs�k�>�IH?k?$_y=$��$U��5�l�<�5?6�E?��R?螁?k�e=����~�G���J���C���w>���ߊ�&읿7���;�
e����(>)(���̠�Bb>����p޾�n���I�Z��,�L=����W=��־kI�~l�=B#
>(���f� �V��s֪��"J?ȕi=�N��fU��h��5>;��>�Ӯ>)H;��v��}@�!���C�=ï�>��:>7䙼H��yG��-��ۄ>\H?*a`?$��?�.����p�k5G��F��`���π���?�6�>ԙ
?��D>���=������f��K�܋�>&�>�{�'E��n��s����"�&9�>ː?�O>d�?�4T?�?D�a?��+?�x?�G�>Ⱦ��U��B&?��?�='�Խ��T�{ 9��F� �>��)?ҶB�~��>��?��?��&?څQ?��?+�>�� �ZC@����>�X�>��W��b����_>d�J?���>�=Y?&Ճ?��=>Y�5��ꢾ}թ��W�=|>��2?�5#?�?��>o��><k���g�=���>��b?�?c#n?n��=�?��>y��>�,�=i?�>b��>�?�O?��t?�5L?���>/E�<����鳽t���'C��N~;V%�<��=��`ev��C�z߼<%D�9ːo��H���J��P�2Ƽ��;�6�>��w>:Ǟ��k0>A�Ѿ���_�>ݱ`���������G�َ�=.n�>���>>��>a�5��?P=Z��>Ǿ�>���?�k? �?ű�:�_���ž��e���>w�G?���=�hn������/r��i=z�q?$a?NOC�&c����b?/�]?�}�=�\�þ1�b�K���O?��
?��G��۳>o�~?7�q?^��>C*f�$Bn�^���>b�0�j�`��=am�>�D�a�d��3�>��7?I�>��b>(�=�[۾t�w��r���?��?���?���?%;*>��n�.��׮����b? �>���%+?Oem���׾�X��,Be�X��K��~����S��\)�����᭒�����0�=��?�q?ĩb?�i?�}��"g��tU�
�{��kJ����N�<�;�A�9��IC�"t������پ��Y���>��\��1?��w�?z�?
9�! ?͓�����+���ʆ>������5�D�-=`薽�2=M�[=0��b�b�v��Ӭ?� �>W��>p;C?�R��h<���+���4� ��]f�=�*�>�s�>�n�>�Nh��fo�:�˽`巾��A�6�; �k>ʠh?�;N?�Lq?
���.��,��x$���[���a�c>�>9��>�D>����n�,���C��t���畑����ݘ=�(-?�q�>���>;�?��?�8��̰�v�j��#�+�<��>��j?Y�>��>�����.��>&�l?�>�>Y�>pG�����4��aɽ8 �>���>���>Z"j>_���[�?Y��n�����:����=��g?ߌ����V� ��>�O?Ks(�gl[<#̠>�v��z���h�B�
�>sc?��=	�1>��ž���\y�g��p�+?���>��&�+�z�K>�?��>���>M�?��p>E�b(�?�+_?p N?+�H?�P�>�WA<�8=*�ʽ�"�Eo���l>��=>S�A=!ۦ==Z�����/4���=d��=W��ke��H�<���r�g�Km�<�0>Ȇҿ6�E������ב��T`�IM��\�����d�x1潩A���oY��W�
♽�@���C���7p�����A�N�?���?z��!�� ���z�/�k�	?��\����0�¾����1���"	��)ھ �G�N�[���J�/h#��~'?�t��4�ǿU���ϯܾ�?��?��y?�����"���8��!>0$�<����g��꬚�[�οנ���)_?��>����M���5�>2�>
�X>��p>E>�������3�<��?�q-?J��>f$s�H�ɿ�d����<8��?x�@U{A?p")�}��f:N=�:�>l�
?.�@>��1�����:��*��>?8�?vy�?�>=#lW�=���}e?�|8<��E�/m軜5�=t$�=��=��
���N>D��>���B�ݻٽ��6>�>�!����>Z�k��<�V]>I�ֽ-���2�?q�Q��sE� 4�0s�zg>0]a?m�>"6m=S=?˩7���Կ�}O��$l?�=�?ô�?��?�����o�>�Ý�\]?��;?�!�>}�G�x���­�>:Z�=t��<���f�}� �k�2)?7�>�gu���	����@�=?��=! ��Vÿ��5�<h!�ZĄ=5�;����0M�^匽�R��V�������o��=`'�=P)1>4E�>��<>�-E>k<c?sMo?�qW>���=�'½�M��U�Ⱦ�Ik=Zހ��\��g4��'bm�����nže�������d����&=�{ƍ=	?R�Ζ��ܺ ���b���F��.?�v$>��ʾy�M���/<�dʾM���J�������m'̾>�1��n�П?��A?����9�V�,��Ρ�������W?{Q����t笾C�=~f���6=��>K�=��3��qS�َ1?;?hS�����>���=�.?�		?H䚼�x�>v�?�s[�Lʽ�jN>��V>�յ>���>��>Kէ���ӽ5?��O?�J	�͙���>p.���?��*X=���=8�?�V�)���u>�}�=�؁��qw�(3�;BU<�W?���>ֹ)�"��ك��@Z"�c�:=rx?�[?��>bk?)�B?I2�<���iT�X�
�@{=8�W?�i?`�>[.���Ͼ*�����5?�e?eN>�ai�X꾍�.��P��?˾n?�D?v�f1}�3 ������#6?�uo?x�l��Y��L�������*?�X�>ڴ> ^��*.>�v?�4�<^4���B¿�sR�?32�?&��?j��=� y���<��?O��>���<ф�+���j���m7/<ڙ?C8��Bb��%�Sߖ<Aja?��?��>m=��0_:�\�=c��ZS�?��?#<���Ym<��9l�ڕ��Y��<"��=�����"� ���7��ǾC�
�򒜾����S�>2C@����>^�8���)<Ͽ�����Ͼ>qq�U�?=T�>ZKǽ�D����j�`u�=�G��qH��.��W�>�G>����+n��D�j��4���=��?�_=&��>�P����������?��#�>x=�>��>S�=Ȫ���?�?l@�}	Ͽv硿�#3���+?,��?�N�?�u?h�|>�ʙ��p辆��=�\Q?�;?z�V?\�ɼe��鍅=�pc?���*f��/�xN��D>��?�V�>R#�Qod<V��=^��>�aI>��0�)Ŀ��@�b�?�N�?��پ���>.��?60?1��!�������x5���J;�7F?1�#>Bpƾ�y$��<�6ቾH�?��2?6a�V��y\? �G��kE���{j���/>'��=,��=Í>괔��j������.O���?8��?�^�?be��7:��9?q6�>,c����ʾ��&<ǥ�>r�>E+;>� >�_>sw���<��!�>�e�?J�?�*?н}��l���2=6�?_��>�+�?��=)��>��=3԰��?�5�">^B�=�y?��?��M?���>R�=��8�HB/���F�Y\R�E�Q�C���>��a?cL?��b>4��\%/�O� ���̽�}0���ǣ?���,���߽55>��>>i�>�D�&rҾg�?�}���տ۔��2w��2&?X�J>��>%X뾤�G�������T?f��>0��%=�������<�䑦?�?b�?�m�!�&���=cG�>��>jk�ۚ�zs����->mF?�7������n�),�>5~�?�k@�r�?��`�X3?i������+��;����}���=�5
?���Z�+>�G?8�=U {�;*��`�}��#�>�z�?���?J!?��J?��������<6;?oj�??���;�G�I����4?��j�~Lx�aG�QBs?���?� @BvT?4D����ۿ�&��5D��N���ـ>��A�{�N>��A<��
>���=�Vh<�r�sV>��>H>Q��=o=q>��n>D�#>�a��qb!�����q����%3���m�Ծ�$�F�	���Y���;㟾�g����ϽA�)�����%'۽�d��P�������?�v�?)b?���>���~�S�~4�Ҭ�>tM~�Z��>��Q?��?�{H?�#+?k>@�_��������� ;��?ǚ�M&�>�w�<%s�>E;�>w��>�>�_Q>���=$���ȩ0>�*�=�q�R�^=Q�>,ŧ>_a�>��>�C<>��>?ϴ��1��l�h��
w��̽8�?Y���L�J��1���9������{i�=Tb.?0|>���?пU����2H?&���l)�Ź+���>n�0?�cW?�>B����T�v:>�����j�m`>�+ ��l���)��%Q>Ul?Eh>��p>&l1�u�7��{O�����Wu}>5?ո�6�.�g{u�a�H��(ݾ*�M>��>�'�Xa�.�����~��g���k=;?a�?A�������t��Ğ�gM>hWY>[=��=$;L>�[��ѽo�F���/=P��=�`>�?��+>���=���>e��PYU����>c�D>Җ,>Ǣ=?v�"?Q��޴�F���0m5��_|>��>W�>�e>�H����=�#�>��c>3t����o�;p��hD��P>(́��a��Jk�az=���w��=�ԓ=BJ
�1=�B� =��}?m(�������W��LʽLR@?�~?��=@��<x�!����{��B�?�a@VS�?S���W�z�?(�?������=��>j�> �;�8P��U?�ѽ�K���:�iR�$��?�b�?�������_Ll��l!>e�$?�|ݾ���>���������Ϸ�OL/<�z>�ZR?�޾�>��(�M��3?Lj?�8��	|��2R˿cm{����>Z��?Z�?6�Y����o&���>К�?��E?� >�:ɾ�B���o>��7?�ES?�j�>�����
?�&�?%-�?L
'>ݝ?jփ?�/?ޥ��_��Q���H�}����<ݧ�=���>!0<�Q)��� �{����'���\��-���\��Ž�)�>�����8���'������&&��hv��:�>P
�> �
?�r�>�5?#T�>�s>��
��z��پi1�q�K?��?����2n�Q<�<㜜=�^��'?�I4?�a[�#�Ͼ	Ԩ>�\?�?-[?�d�>a��9>���翿�}��2��<5�K>5�>-H�>X(��3HK>��Ծ�8D�cq�>�ї>���@ھD+�������@�>2f!?ܓ�>�Ǯ=�� ?�#?�|j>6"�>LdE��8����E����>Q��>�B?��~?��?xȹ�3Z3�&	���硿�[�A5N>�x?�V?�ʕ><��� �����E��&I�����x��? rg?�B�l?M0�?�??��A?[f>�|�sؾ����K�>�$?P,&�lQ6��$��+G��>��?�L?�g�==���r#�������)"?��n?=�.?�U�{�a�V@Y���#<W���\!<0A-=��)���=:6C>����l��=>x�>������v�=�aH=�D>&�> �7�0��,?�Q�s����ϓ=�nq�VSE�+�w>]&I>�����{Z?C?�OAx��뭿ᑜ��oa���?e��?�Ԗ?�ꪽ�{f�U\:?t�?o�?�>.1���ܾ��s~�ƴy���>n�>��3�Ӓ۾�:���ʪ��	��]˽:L�����>��>��?�;�>g͌>B��>�r���52��S���?�{X��J���4������!���`CM���a`־UG�����>��"����>�!?,fB>�\Q>r:�>��=���>A�t>�R}>AKR>Cg�=��=|*<���)��R?�"���A'���辅���N7@?4�d?��>F�H�����Jr���?싒?ȷ�?Y>H�e���+��?� ?,k�!	?^bE=������m<�᷾)��0���r:�'�>!�½��;���L��]���?��?4����ɾ�U�_���Gg�=�y�?-?��%�"�L��er��9X��R�܏_������ڤ���!���m�y$��o ��i`��� %���4=�$?�m�?	;�����ܰ�U�c�"t@���[>�T�>��>�[�>	)D>n����6�E�`���+��牾1��>�w?���>AMI?t�;?��P?��L?Ʈ�>a�>�@�����>�>K;\�>[�>o�8?�-?q�/?�s?n+?��e>9��ѿ���Iؾ\3?��?T�?�h?<�?�F��7ƽ�,����N�Q�x���|�1݂=Y��<.%ؽ �p��fX=V�R>�S?�x�N�8�u�����j>tn7?�:�>��>�폾�K�����<��>=�
?v/�>c ��}r��n�S2�>f��?���F5=�*>�m�=N셼�6Ϻ���=�ļ|��=���t�;��V<��=�Ô=�s���h8S;��;�e�<�=?`l$?��n>5��>����� D��H\=\�=����Ի<�n���1���@��,W��4��>$Ĭ?wc�?��=��>�Ho�4�]��v	���0��uݾ�ٛ�Mc?��?�)2?���?	12?nEO>���=ˀ�,�~�d�{���z�V?#+?���>� ���˾e����2�a�	?� ?Cf]������(��D��^ί�o�>��0����/د�9�B��<b	��吽V�?m��?O T�X�3�.�������z���C?��>lޡ>��>��)��f��%���=>f�>i�N?��>s�l?_�?��k?N��=�)��������d3=�Q8>�W?��?M��?N�u?�w�>��w�{���P��#�1��b�������"����<x��>�u�>��?��>B�=Ȑ�C�i�m$<��=���>SI?U@�>m4�>�u>O&�<�zH?��>��q'���¾��h˽=���?�2�?�b4?�s�<�'�am2�]tƾ�1�>${�?�?��%?㆐����=��!�����x_�����>���>�$�=�K-=�A�=��ܻ�>�0o>ɯ��_F���-$��~	=�B?ֻ$?Z��=c�ſ�r� C�˜���<Pˊ�KBd�ċ���V�T��=s�������@��<�J�@Ξ��V�������ǜ��G�r	?�׋=B��=-r�=ى�<[�ּƫ�<��Z=B�p<��=��[��!<��g�2Ɠ��s��o�����;'�U=a@;r5˾�?�M?R�+?P�B?�v>�	>{=\��>�e���?Dq>�#��������+�M�������"�ྗ�޾�$f����3�
>%tV�}l>^�4>�_�=�ɡ<Ed�=�=�f=hb:Ɂ+=�=�˲=v�=t��=��>��>��d?����Ur��@Z���P>k�?K��>	G<�J㾈3Y?�?�Kh��j��R%׾PK�?w��?n�?ψ�>B���Av>A�^����A��=X�p�i����=1�����>t��>��B�ź�������W�?њ�?��??8����ܿ���=K8>�S>vrR��t1� �\�B�c�
�Z�>�!?�;��y̾h�>�(�=ME�'	Ǿ�s'=�`7>4h=^��[�h��=�7}��==0�m=[��>dD>ܸ�=�ر���=�3I=ic�= P>�ʕ�J[5�՝'�<�3=K�=]0b>��%>���>�?h�4?�4`?���>H�؉��x�˾Ӂ*><b,��G�>���=@��=�ɀ>��3?,_>?�KO?�b�>�B4=xK�>[5�>i�1����q����ƾܠ=�k�?Ub�?C��>&��4y��k�������w?�� ?��>;��>��
��7ȿ��K� bH�܂f=�_��.>��j���:L�x����;��>륹>��>w�
�@N�<3��>���=�&�Q�>��=j����=�=��-��=�I�\\�ݧ��8����Ǽ�>�i:��= �#=�)�<>� �������;��%>��>n�->�t�>�C�=y���H�=�4�N�Gh�7����+�&�k�9�~��O(�h7߽|�R>^>�������|�>��g>���>]��?�K�?��8>��~�B���쓿�LB�Q� �X1<>M\�=A ���*7��`V���8�<�U��>5�>�5�>�Lj> I.���=���'=��ݾ��2�M�>֎�:��E��M0q��U���+���yi����g�F?N������=��~?��I?d}�?���>�:��c2޾-|/>Ft�mL=����|�����~?��)?^I�>���D�:q��!��p�>=]^�{v��E����5�9��U��(�>��������o:���ܒ��U>��{� �>zm?f�?uھ�gU�`9g�����Ւ�w�/?�$?�ԓ>p>&?lU'?�fF�AbD��׌��*=�6�?�e�?0��?5�>��=������>�i?8ԛ?�ޏ?Xq?63f�Gd�>��v���">[oI�x��=���=RI�=�8 >z?Yl?�5?^��=B��{�E���X�a���<�$�=���>aŐ>Nev>���=#5Z=�<�=�6_>��>��>9k>M�>�>�t��h3��$(?D�=z|�>i�B?��~>c�<S�0�P�>�SԽ�~^��D�Ҟɽ(�ý�<*E<��U�Z���N[�>q�ĿfA�?�L>#] �!? ��ˮN��o>��D>x�ܽ���>��J>"��>b��>a�>�Y�=��}>>fV>��ƾ��>IT4�c�(�kgG��P�����;�>�y�������C�LQ����%������z#��G����t,���<>��?�uD=�F����&��<�>��>�e??:�_��J�II(=�t�>���>�������)<��S����Du?��?��>��>�:?��=?�>�=*���g�$���<.X�)���On�m�t��k���!�Xc��`N?U�q?FG?��=0C>�?�c\��疽���>�[>����3\�<���>���͂8������þ�����q�=��?Z��?�xl?���(F|�3Q.>"�<?�$1?��t?�0?>;?�{���%?�\/>��?*�?%�7?�.?.:?
D.>S+�==�M�a6=3ڐ��C���aȽ�ؽ5�ؼ1�F=�o�=�\;8*<��=�xq<�� ���ۼ�L�9q3�����<��==>�=�z�=H�>�G?e	�>�ǿ>
�I?�.�+�����ӻ>��h�}���EZ ��C �3���i<��c?;G�?+�?^�6>�Q)���C���l>�`�>��>��>\ٹ>_�!��3f�Ɉ�<%�%>:�">B�3>�_,�\!ҼK�9.��0@D=���=�?�3B> �=к�>�6���׾�	�>pz=D����!���n9�?{`�ܹ8���8?�C?c��>�=�=�Hվҽ��E��O?D':?�fc?�_?G�c>hW���G��mR��U>q+>��zx��إ������q��;eG�>��Ⱦ�ޠ��sb>V��dp޾��n�fJ����t)M=�u��	V=C�v�վ���R�=��	>>���� �U���ͪ��8J?�
k=x��fU�9f��:�>'��>ٮ>m:�0�v��@��������=���>c�:>:��d���yG��*�?L�>�HE?kO_?�f�?�܂��s�;�B��k����� ;ɼ��?n��>�a?4�A>!=�=O�������d�'�F���>���>����G��f��`����$���>A?w/ >��?ٸR?��
?�`?�*?AM?�M�>������A&?߃�?A�=�Խ��T�M�8�E�E����>J�)?/OB����>��?.�?��&?4wQ?�?�1><� �wF@�Y��>�O�>��W��^��\ `>��J?g��>�,Y?HЃ?��=>^�5�f��E�����=�b>��2?3#?}�?.��>��>����=y��>s6b?��?^p?�O�=��?�I4>��>��=y��>a��>[�?_�O?�[t?H�J?m��>D��<���r���{�5�C��9�;��<f�u=�	������Rc�<Ov;፼ϝ,���μ�+M�-���w�<x�>O�s>lx��J\1>f�ľ�U��j0A>'���*����h���9�ڕ�=�n�>��?h�>]U#��d�=r�>1��> ��(?_�?Y�?��:E]b�sھ��K���>d,B?6*�=-�l�mf���xu��d=s�m?��^?.IV�8���&�b?��]?Dg�7=��þ^�b�*�龚�O?��
?��G�6�>��~?��q??��>��e��9n����ACb���j��Ѷ=�q�>BX�:�d��=�>!�7?�O�>.�b>1'�=�r۾{�w�mq���?]�?��?���?B-*>��n�:4���╏�Wd?*�>�L��ʇ#?rO�;ҴѾH뒾~���3�β��TǢ���q���E'�}�����A�=�?�#u?�Md?hr_?�����b�&�Z�bp�v>R��8��l�@�D���B�M3A�n���	��yᾉy��`E`=<{a�)�/���?sd2?�:�P&�>l��K"��e{��A>�%��-�p�=na���� =#�<6X���9�Ӫ��
?�>[�>�#:?�T���:��P(��A4�:��>�E�>'��>*g�>�6��0�b�$���ʦ���D�I��I;v>�sc?�K?�n?<`��$1�Z�����!��0�F^����B>9^>w��>��W�=��99&�Z>�D�r�����u����	��:= �2?D-�>���>tM�?@?2w	��`��onx�
{1��G�<�-�>�i?C5�>�ن>н�� ���>��^?@�?��>TTH�7-��2Y�A���&=�>�F>�e�>�.�>����)Z�����3���6��D>�e?�T~���6�鱛>V�[?��s>F��=`�.>V����$ �	��DN���#>�=�>�+>;�o>Vͨ�����d� 3��?f&?$��>�.c�z�4��zh>?~K�>���>yA�?7�@>����{�U�NO�>�r?��a?`m?:ɭ>5��t���׽u�$�cP��Jf>WS>�*�<5JM=	��Cqz�*k,��Γ<��=2t=H~u��s�=d�6��h���ʽ��u>�Կ3%<��V��:龛��H}�������V��e$��j�|g��|as�{J���ֽk����p��7	��&���U�[��?��?�����o��)H��3�o�v+/�\�>��O�T����Ѿ��F���������gھ�(1�}�F���Q�m�:�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >`C�<-����뾭����οA�����^?���>��/��o��>ޥ�>�X>�Hq>����螾|1�<��?7�-?��>Ǝr�1�ɿc����¤<���?0�@�kA?W(�6���<T=S��>�@	?LB>�5/�]��Ʈ���>� �?��?��I=t�W�@����e?�5<g�F���ۻz��=�1�=��=[��b*L>8ߓ>���;@���ڽ,�3>q4�>�d$��r��[��(�<*�_>�4Խ�ʛ�{}?WW�Zb�!�?�F9^��JH>�g?���>]�<`#?��T��̿d�/�١{?���?�f�?<�?���X�l>�ɾ:�B?��?�-�>�fJ��~��ĭ4>g��\����8�V�k�*Bk=��?3��>m~� I
��h|��=�K>-���!ſ�%����I��<�w=;�O��˽D����;��Ւ�`]�����D��=T��=hIB>`�u>K2L>Q>�J[?/|j?,�>z>On�_I����о3����*x���$�=R����#�����w��W��.�	����<���xþ��<�[�=PTR�.����!�^'b�ϐH��?.?(&>�I˾�*M���3<��ȾRz���褼����AξVe1�8�l�f-�?܊B?�ƅ���V�`��F���Ľ�V?�Z�J�^���n�=��Ǽ�k�<X��>�Ơ=�Ᾱ�2���Q�[C0?3?���~ŀ���>�r����=�4?�o? �=��>�-?��"��߽��>	 >Pա>o��>?�<>{ ������?�??��7������>�����c���>c)J>�%C��6�Y�z>J09.�N�1=#f��k��O?�(y>+-��+����)CD��Z�=�E}?{��>C�>�Sz?�N:?�F=o��lJh����@h�=c4W?��`?��=�%���Q���i��mC?�XX?�wP>`|T�������ב��[=?9�w?"�'?H�0;T�l�6�����f�0?��h?{�m��������P�
?T-?�˼>�)T��*>�4V?m�������\����,!����?1 @/�?��>��J��<��>*��>v̔�%�{��d�nSо�E]=��?�s��r���)1��k���Z?���?��
?�^���*����=W���ˉ�?�/�?~ة�59}<ٱ��k����� �<"Z�=�[D�d���7�#/Ǿ�
�Oz���ü��>�)@�s��>e!9����	ϿC腿��Ͼ��q���?�l�>>!Ƚh�����j�6	u�UG�iNH�)��t3�>��>O ��j����z�"�9�+�-�w��>�FƼ^�>rER�ޑ���C��yZ4<���>���>/�>,/���E����?���DJͿHs���G�.�X?Uj�?�|�?�3?Q�;��{������[�!H?ǥt?Q[?�����a�_G���j?,^���S`�׍4�zHE�-U>�"3?JE�>�-���|=�#>��>�f>�#/�W�Ŀ�ض�]������?l��?on����>���?#r+?2i�
7���W����*���)�z=A?�2>�����!�.=��ђ��
?�}0?Lx��.�:X?��P��`�q�7����<��>�F��FcѽS�9�/ǽ��N������\���Q�?���?/��?)����D��?3!�>�v���þ�U=��N>��>���>�S�=�Ç>�e�8!V����=̼�?t��?��>,��ٝ��E�=�sv?Jf�>��?���=7P�>MP�=Ib������^&>��=URK�EF?�N?dv�>��=��?��j/���E�1�O����C�B���>qCb?��M?5�o>=���6F�k� �nȽ��;�y�+�R;���2��-սrC8>>�=>��>1D�vξ�t?r4)���ӿ-���� g��C?M!�>���>�^��˾�s�=�#n?Nń>�A,����4X���𦽶��?i��?��>�!��i8�;�+�=���>�C�>d���otٽ������=DyE?�̱���|��ST���>��?)�@YT�?@3X�#�?B���_�����݀�i�X�>\�1?*	��.�&>�N?�/>Fm�����o�p�Pհ>�{�?+m�?�w?��b?e�o�՘8�}�Z=*b�>8v?��?��鼫h� b=>�Z?����֋��]�xFl?�Y	@!�@`[?zt��3߿�!���0¾+�����m=�w�'g�=�?�]L;�c�>ֻ>�4>G*�>6��>\^H>�v�=㤩=�>�Z!>~��l�"�~Ű������wH�~ND�fE��;�u���s-�/D־��"��䗾Zϫ�����G�LX��=��q��>��Z?�g?��?�6?|g=��%>����|˽_\$�8B'��9>#V"?"SD?��)?g=桾[U���y�cw����(�~�> �>�'�>t�>�B�>��߻U5>3	/>�y>�u%>6��=x4�0���z�=~%�>3�?��>�C<>đ>9ϴ��1��Y�h��
w��̽2�?.���L�J��1���9������i�=Fb.?6|>���?пG����2H?���s)���+���>^�0?�cW?	�>��U�T�:>����j��_>�+ �~l���)��%Q>]l?��g>�2s>̀3�)8�I�P�)���
U>��5?纶���9��v���H��0۾1Q>�Z�>ި�s<�l�Z~���i�US�=,:?j�?|���Qb��m�v�N����VN>��X>@�=� �=�xM>-�b�h�ǽ�H�4�-=���=��\>|0
?i>>8��=G��>p�þ;��=* ?���>�U�>`t?)A?X�>3~��X��� ���Բ/>�R�>>��>���=�L2�햡=�*�>�=���<>`>�Ϙ<BD���xY>���;館�{(�3}�=|�<�v�>F�w>��=���:5�f�;{~?@`��OՈ��^뾂����:D?lt?�-�=�9<{"��	���蹾���?��@'x�?o	��oV�VG?`�?���N�=�q�>�L�>�Rξ'wM�qC?�	˽\8��-�	��#�l�?��?}�/�X�����k���>ރ%?!�Ӿ���>��=��������#��� q=�Z�>��3?������k���uk?��>���^���y컿�~\���>�D�?�ފ?����$��nqj����>�,�?0z?Z�]><8��Qɾ�Q�>WuW?�sT?I%�>2��]�3���?���?��q?�_O>��?n��?%J
?b��=)
���F�h��q�=r����=�S>ϊ���:������v���x��G辛I�>�N=2��>6�-�Է�V^=��>�����������>;[�>7&D>(�>���>$ۚ>t�e>M�¼A:ý�r�����k�K?7&�?v��b�m�jp�<-��=�T[��G?e�4?��S��о_i�>�>\?���?c�[?�-�>K<��F��6(��7 ��ma�<,�K>�q�>3E�>K���Z(I>\�׾�K��>�>�±�`|۾�7���>����>�!?m��>�i�=�?��?�w>v�>5g�����iA���>�7?x��>�b?Gj'?F�Q�1��玿�򙿣�K���N>���?��?;w>{���Zϖ���%�S#�w��=��y? Dd?���=��C?�q~?7�%?�=?l31>��G���w��Q���p�=t�?.������p2�[\���?3�?�h?c M>*��Q�ٽKg1��1־��3?Cxt?~^Y?�b��i���o��jݺڼ��d�)@=l��<�3�=_�=U���FC����=	Ԃ=��!�o�սЈ|<9y4>R�h>9�L��
��Z��;*<,?�G�d׃��ۘ=�r�L|D�(�>�UL>����Z�^?�R=���{�0��Hy��~#U���?˝�?�j�?� ���h�<!=?	�?�?%&�>3G��v޾���Cw�Zqx�ls���>���>��k�z
�K���d����E����Ž8�>��g?]�@?�-?_)�>.8�>�%I>�N߾��@�� ����&��fS���L���6���ھli�Y9-�n�����q�0x?��¼9x>�c?4*�>��>j�>�>�_>���>��>���=��t�p&���]�PC���IR?����9�'��������f-B?nsd?^'�>�=i�̈������r?���?�t�?�ev>�ph�L++�sb?�7�>���s
?y:=C�9�<�Z�����Ƈ������>�?׽7:��M�pf��a
?�'??ō�5u̾ab׽�����'�= 3v?# ?a�0���I��l��+EN�iHC�Gv}�yGe��	������tm��u���d��]���-�%�59a=�/8?�?�����򾀮��`�j�TgG��\T>���>�ǔ>���>��G>�v�[�:�`�^�jb"��i���>Y�x?�׊>��W?K:@?׬`?	�S?)��>g3�>V���s�>Ea���>���>�l3?:/?	�0?&?�$?�g>��|����þe�?	�?�?$T?�"�>��w�*���aI;PZ�:��Y��IJ�d�<�+K��
4������=�DY>`X?R�Ж8�+���Ȋj>V7?U��>��>�ُ�����<t�>��
?��>R �\sr�)S�Z�>U��?u��p�=��)>��=��� L�����=\D¼��=Ty~���:���<rٿ=̃�=�s��kָ���:��;�5�<�=�> �?�1�=[�7>�G��� �~��к�=A?>��=��#>,�������}���[o�e�>U�?��?�ɳ�ߊ>1�&�+0�k����[=�T2��W,>nGA?�N?=�S?�J�?�J?�K6?����E�{5��u$������a7?G!,?"��>D��2�ʾ���3�{�?�Y?R<a����<)��¾��Խ!�>	Y/�-~�����D��������t��a��?꿝?[A���6�J{�^����]��`�C?��>�X�>��>��)���g�%�/;>��>�
R?��>{�O?lJ{?�[?��T>}�8��$��Nș��E5�K�!>��??w��?��?Ny?�V�>&t>'�)���߾_4��Q*�N�򽎼����V=��Y>���>���>�>;�=ߵǽ�2����>�2��=fAb>_H�>�g�>p��>axw>�<�\F?]��>q�����M��2�{���� ]o? ��?��5?��B=���x ?�[���Kw�>�Ȥ?Z��?�3?p�i���=�����n��ov�� �>�F�>zT�>�5v=p;�=��>��>Ӫ>7����v(�(1���?+VC?�M=Ĺ�Eۓ��Mپ>���a=Ҧ�b���s>�3�ǫ>¼�=�ƪ>ې>kF��B]�H��)F�������˖���>��=2+,>!W�=\G�=��D>x$�=Z/>/��=�4�V3��,^���3���5�����8ǔ=Ğ4<Ȑ��&H=�Ⱦ�L{?(jL?I�+?�oC?��~>Mr>�C�i�>��r��f?�mS>orM��Z���8��ਾt{��+ھ7)ؾ��c�=���=	>U�)���>�03>���=>�<z3�=Bk=���=	"�:�8=f$�=:1�=�
�=���=>�>�>zY`?��q�ʏ��u�m��z >Io?֔�>N��;��|�]<?��>%g��|���Ⱦs2u?���?���?A��>&Ӿ/]�>��#� �y�*�=xrC=/9۬w��A�c��>~�>�/�����6W�LI�?���?�M?=W���K��a�д7>� >��R�O�1�y�\�x�b�QmZ���!?mD;��?̾]?�>� �=*߾��ƾ)>.=��6>]ub=V^�VQ\����=v�z�T<=�l=&݉>�C>�v�=^*��E�=O�I=���=.�O>����V}7��,�e�3=���=h�b>�&>�C�>��"?�2?q;d?���>��v��ξ�����jM>-�*=��l>���h�=ę�>�/?�K?<)d?Om�>_戽��>�fr>+�.�����cF�����g:+��?&��?\U�>'=�<S�޽{��|�U��AA�S�>�<5?�k?�F�>����Iٿ o)�`="�F���x��;u�<�!��Լ7��:�F���]�ҳ;>�U�>ƴ�>8��>i?/>��>�).>���>k��=��;V�='�>�C֘=��>;��F=��<�"�<IwT����/h��O�]���<����<6�_��#�9�.'<���=���>� >���>��=�߷��1>c���nJ�v�=E⣾~�>���a��~��P0�H�<���=>Z\>F)}����Kj?Mf>��J>�W�?�Du?�I>��s4Ҿi���g�u�3mH����=�8>��5��a9��p`��8L�� ;A��>���>o@�>�0j>j�+��\C�L+�=�о�-�~�>�Nz���>�<����q�Ң���Ş�!^d�m��<��A?�����=�5�?dO?�ؔ?^�>���eo۾"�4>���}��	�kp�
p>�D?�B$?x��>=���2:�>7��"|=�>@G�ٌX�pI����r�f�R�}����>�}i��8��5�,��c��<^���O�l��-�y>R�]?��?�8ɾ
�h���N�����|w��a8?F?���>���>�V?�=Y;r��(����a=d�m?2��?�?�=�>�[�=`հ�ȇ�>C�?O�?�V�?z�s?�u=����>��<% >>!���{�=�u>�K�=H�=��?�
?�	?�眽O	��C�4o�O]�N=1�=QƑ>P��>�p>�D�=�Q=���=�B_>(ٟ>FW�>�Oe>�><և>hC��C��$(?���=��>m=2?21�>�M=D!�����<^C\�x�@��r,�<A��l#����<����1�D=�ܼT�>ǿqK�?�vU>��	T?��񾃽'�o�R>T>V>��޽�Q�>�1I>}}>J�>�>cr>>fn(>O�վE�?>z�����.�L�s�I�����dl>C���H@�U��ٽ&.�� ������s������9��O9=^Ζ?,��tg�V�)�����%�>�yh>�')?��q���>�4��=���>�]>z����h���ľ�y�?0�?$uZ>���>�G?��K?`��<���̐��?��f`��[�o�d��D��piy�o��Տ��V�Y?'iv?�C0?Y;C��>,�?��v�����Z�><�7�Z�4��콶F�>m1�����ھ	���z��K�>dX~?���?�?��ƾ.�m��'>�:?Z�1?�Mt?��1?��;?U����$?�x3>y9?�l?ZJ5?z�.?�
?��1>���=\���R�'=>���ꊾ�ѽ�Fʽ���3=9�{=+R���<�u=+�<E.��ؼ U;g����Z�<�.:=��=�/�=jK�>>G_?$��>4��>c�8?4�د7�7��j�,?kY2=,�������z���W��>��h?���?ǙY?R�]>u"C�@��o#>�·>�7">�}\>^S�>����A�i%�=��>��>��=Ub�H慾k(�&���O*�<�P >���>y�>�K���O[>ԲB�^.��H>aGᾬ%��[���b�X�V��E��$?��e?MT#?q��<����S�P�E��!I?VTN?�،?@"Y?=��<b��z�q���f��-���~>�{����.�&���! ��F�8�*>5��>��ʾ%����b>,8��༾�0k�<�Y�i���ۀ=!�
��X�<&'
������@�J�J=/[�=Eپ�R&�V~��z���U?h[\=�˰����S_��r�>��>���>��S�b=���C�@|���s�= ʶ>M�>>v�(�60쾽�9����xs&>��\?��t?Ⱦ�?�o���Ub�ԩF���wΟ�Z�;��7?�u�>Tg?��X>���<����&�G�j�.^U���>���>.�}�5�� Y� �Ǐ��q>�a�>)�>ԁ?tQ?��"?Ơo?��3?l?ܖ�>)� ����h5&?�|�?뾄=��Խ]TT�G�8�( F��n�>e)?��B��#�> W?o�?��&?#lQ?��?1x>͊ ��M@���>.~�>��W��W��R}_>�J?��>YY?5�?n>>�|5�*΢������-�=f>��2?�^#?��? l�>��>$-��OP@=N��>��Y?E3~?�#p?[>D�
?L">{�>�|4=pE�>�>TW?��N?�(v?�TJ?S�>-/-<%����ֶ���N�:]���d�9X��<r�J=��'��Q������FP�;�� �xT�<��=& Z�X���m�)����:���>�s>򕕾W	/>X���o��2�A>�6��w���	�7q<��5�=�I�>;�?��>Q� ���=e�>���>�&��)?�}?�8?=a%;��a���ܾ�yR��ӭ>�A?���=)'m��f��lQu�n�_=��l?�^?�NT�����+�b?D�]?�h�=��þM�b���O?��
?��G���>��~?��q?��>��e�w9n�J��5Db���j��Ѷ=�r�>�W���d�A�>)�7?]M�>q�b>��=�t۾��w�jp���?i�?��?L��?�+*>�n�4����>����%X?4�>�w����(?���)!ݾ5I��J�����r`���߽��\���㡾�>�Ň����98=�
?j�c?;�x?U?���jf�"�b�4����J�>�
�Ŧ$�M�6��bB��D���e��:��վ�\]�,��=g�~�k�@��0�?�'?V�0�^.�>�Ù��$񾹦;h�A>�v��������=�����9=��N=�j���.�s���T?k��>^��>QW<?[��/>���1��38��2��Fg2>v�>��>A_�>�C��*/����_ɾɃ�^нA	Q>)k?�gT?\�s?���?�,��,��7�#��3I��:��Z-�>�>>�)�>��C�I�+���0��E��Nt����j"�������F=��,?)T�>"~�>��?Ǡ�>�h窾�e���#��j�=�G�>�j?�+�>㿆>���r�(��>��y?`~?Y�>�������jo��-��5��>�!�>�?2��>V/�oG�&I��h���A�}��=�pd?�B��U6��K�>b�U?0�f�\]�8XX>y�	�q
�8���=�2�>Bz�>���=��	>��9!�|�w�)����&?���>�����+���F>�c
?�r?�Y�> %�?�up>�O̾X�<��?da?��W?��A?|>�̀�!�=h����^�oZ�;6�>��>}O^=��=��½;�������<�R>�݈=�[�� ً=Q���R�T�T���F>oJ��6�5�B�þ�m��>����0;�8�ξ���=GpA�'��J���S��D���qQ���I�Fe��S8��4����_ѽx4�?f��?�YƾxG���6������D�5�ކ>ٿ��E["�+�Ͼ}�˽.�0��}���˾8�@���\�I�.��a1�B�'?躑�ͽǿడ��:ܾ�  ?CB ?��y?��&�"���8�^� >KM�<H#��s��\����ο����<�^?j��>��0�����>Ŧ�>ۡX>�Gq>��鞾#/�<w�?��-?s��>7�r��ɿO������<���?��@�fA?��(���SU=�q�>Lh	?S+?>�J1�x'��[�����>%.�?%Ɗ?��F=� X�����e?1�<�F�f��"��=9Ʀ=#9=�	��J>d@�>�2��hB�޽o�4>���>�%��f�Ac]�>�<Ld\>��սWY���2~?y�|�A�m��jI��d��y=>��S?��>&+8�th:?A��@�ѿU�Y�{�\?���?�:�?�'?��)�s=ᨾR�O?J0?���>�PY�д����>��n��}���D�}������?g��>hlo��l��֎@�,�=~@Z>��,Lƿ��#��!��v=�Aϻ.W���ٽk���!uJ�w���y�k�C�ݽ�}b=d�=�qL>��> �R>~X>^�X?mm?ռ>�>w�����.}о陻������Ջ��B�@������<�ᾍ!�ѧ��_�lV����>���==�Q��D��u� �I�d��MH���.?��">d)˾�M���R<�gƾ�����I��.���H�;��0��m�<�?�HA?�ⅿhOS����V&�%D���WV?��ʯ�Zή�*��=؅��;}�<VΜ>�H�=��⾢�1�D�S��0?.?���в����=i�V<�=o+?q�?�9�4-�>�?}����C޽oX�=4L>H��>���>&9>X���%���`?�cU?�Y��"K���Ĥ>Ze���蘾*��9�8>����G��Ɲ>i�B>�`��7��G�`i9=>�V?��>�(�I]�w����k"���]=	ky?��?B��>�6i?&�A?W�<���]S��A	�:Ԁ=;�V?�i?��>#l���Ͼ䛥�c�5?1Vd?�/I>�Gc��:��.�����?�(m?��?'�����|��l�����{5?�w?�ii�v���+�G�Y �>�D�>�.�>%;��̰>�DB?�ٽup��p���m�(�_u�?l�@�h�?nI���[+�̼?=�/�>���>�gĽyj����M��_9R=L� ?��{�ݽ��1a�=WP?x��?B��>+������=�'��0Q�?p�?�p���k<#��;�k�IX���q�<t �=����"�Y����7��eǾ��
�ux�� ﹼ�H�>\B@���)�>�8��⿃CϿ%���:�Ͼ�=p�>�?��>�Qǽ������j�S�u�#�G���H�����lZ�>�8�=�%�*cm��x���5����=���>���<�݁>��ؽ�������f[,��I>���>/�>U	a=��s�?�?r� �y
������.-���8?h�?���?VyZ?���>�t�������>5JS?�pY?Inc?��=�ᙾ8)�=j�j?)^��R`�̎4�\HE�U>�3?OC�>�-��|=K>3��>�b>�$/�؎Ŀaض�A�����?���?[p���>���? u+?�f��6��JX��D�*��L:��8A?X2>'����!�2.=��˒�o�
?�y0?n{��*�=vR?N+P���[���B��]���{>�=�8��5>�`�"[���"|N�֩?���?�J�?�ކ�&E'�5�H?�j>��Ҿͤ辶+�;5��>��>�Ad>;�>���>ږ��	;�2�>I��?���?�6�>T���۳���O=;�?]h�>���?�*>hA?�ͥ=r���Gv.��	>U��=d$�	 ?�O?-�>l��=paR��
=�D�M�n�Q��:��EE�+y�>u�_?}�H?��Q>�>Խ��P��s!�\�н��!�x��<����)�ꮽ�P8>�@>,�> �f�f���?Tp�9�ؿ�i��Op'��54?%��>�?��{�t�����;_?:z�>7��+���%��|B�`��?�G�?E�?ǻ׾�T̼�>h�>J�>,�Խ����n�����7>*�B?W��D��j�o���>���?	�@�ծ?ni��?�x!��>����x�(�@�x��"�=M�A?Qb��M>�?+�[>?�g��W��f�v��s�>�?1�?���>+�q?���z�Z���R���?�|�?��>�U۽/p
����=���>sB��タ��ܾ��?9�@��@neW?e��Nhֿ�����N��֗����=���=/�2>��ٽy\�=��7=��8��H�����=`�>�d>q>�'O>`;>��)>���3�!��q��H���+�C������Z�#���Wv�0z��3�������?��U4ý�y��#	Q��2&��C`��]�/�?�ԅ?��t?u�?��½<~f����9܌=���E�>��?4�?��n?�
?~#l�$|��o�}��懿ξ��y���M�>�0����>�Ӳ>�O�>���=�I>�;_>0E�=&f�="=2o�:�n�=O>˼�>h>�>Y>�>D<>��>*ϴ��1���h�
w��̽@�?����J��1��U9��#���-k�=�b.?/}>����>п����s2H?	���r)�m�+��>��0?RcW?�>�����T�f9>@��Ӥj��`>�+ �o�l�|�)��$Q>l?�T>�Y>[�/��O-�.C�Ex���n_>h�)?��ǾX&���k���N�O�߾��Q>@/�>󲪻F��^ŗ�x���Z_m�@� <0D?��>�@
�j��y���<��4[>�<>0�껣n�=x�3>�������JL���#=Ϫ>��_>��?Ke>���=���>�|��Z]��K�>�k�>(ك>\�M?dR?7k��cA�1�t���=��h�>��>,�>%4>%�E���k=do�>w"4>.ጼ��<����*�i��>�g#��k|��Ž[l�=2A%�d�=�˞=zսZ:_��>�<��}?(榿b���[U�롰���B?��?ՙ�=ߘ�<~%"�g���9������?�e@q��?ކ�pX���?_��?��~��=�m�>�>�Ǿw/J�,?9�Ľ����4���"���?��?�"��Ê�X�k�0�>�+$?Ӿ�d�>ڀ�Z������u��*"=|��>�?H?XD���O��=�{
?�	?\n򾃪����ȿ|uv�s��>J�?$ �?�m��B�� '@�2{�>��?�gY?�hi>.f۾�sZ�M��>Ȳ@?�Q?*�>7��'���?�ݶ?-��?+O->���?�#{?gb�>숹���*������{����p=�*k<�^�>*�'>����\{@��璿�R��x
p�����M>��4<P�>�{ӽX���3в=�����Τ�Jj�����>�>m>�Hj>!2�>'L?*�>NP�>��=�|�~ԍ�=�~�K?|��?/���2n�CT�<9��=i�^��&?�I4?�m[���Ͼ�ը>��\?q?�[?d�>]��N>��迿%~��`��<��K>4�>�H�>�$���EK>�Ծ�5D�Vp�>�ϗ>����?ھ�,���S��!B�>�e!?���>�Ү= ?ou#?%�j>Y/�>�VE��'��Y�E�g��>(��>�?��~?��?޹�KX3�,����š�B@[��/O>��x?�H?$��>�|�������W�EIJ�\��ǂ?��g?r�߽�V?��?k�??��A?f>�f��׾>��V��>��"?n���� 8�<?���O=��4?0n?1��>��k=w��=��
>&L*�B��ؙ?ȿw?4@?þ��V���������`ٽ�d���=�Ž�8�_�)>�7��=2Y>�X=�����W����=�0>sU>��/u��f����!,?�I��)��3,�=Ǡr�&"C�mx>��M>�Խ�l�\?[�=���x����m�����a��Ռ?;l�?Q_�?�\�g�{;?ޗ�?x?@��>�����xܾ0Sܾۛ��N}�W/�́>!a�>S�C�:�߾Yw��]���ռ��n䳽<���<?V֣>��,?��?�Ck>q�>ľ��J�(!�R���7_6��E!�'���G�m������h���1�{<��ܾ��&��T�>T� ���
>��>���=j�>Ju�>��=W��>9Y2=d�d>��=8����D1�roh�%eK<:b;���M?�U��?a#���澿���-?Wlh?y�?_T�<&�u�.&��%?3�?���?���>�A���?�r��>�"?�J��M�'?��3>`��<���=�`������,s�*k��m�>z���/�:�>L9�z���g�>.��>*I�=!��H]��~	��a�{=S΄?Da)?S�)�7R��p��V���R����g�I����#�?kp����������)����'�p�+=g�*?���? {�Y�������{j��>���e>�.�>YP�>fx�>*�K>'��4�1�Q�]�Y�'�<ބ���>c�y?w,�>&�I?S�;?x�P?vL?vt�>'�>b�����>niq;E	�>W��>9?*�-?�<0?�0?�+?=qb>����SK��r׾��?~�?��?��?G�?F�����Žˆ��1�\�Auy�Y腽{=ү<GHܽ�r�lj[=S>�X?M���8�5����Lk>sI7?+�>S��>�!���K��bz�<�9�>��
?᥏>�����r����΋�>���?;���>=�)>��=�.n������_�=֙¼�\�=�!;�5/<%u�=T�=�_���W��;`1�;G��<gI?��>��i>v>�g��nԼ�3]��B޽�e>�x'�ؕ�����_�T�0p��9Ć�6�w>?�?�w�?��[���>����5$�d⾾GD�=��������N6?�6%?�>?�M�?5JX?�$�>��e>�\�����[qW�4��I�4?,?ܸ�>�����ʾ_樿�v3���?5R?�0a����^*)� �¾8ս\�>�Y/�s;~����#D���y����B����?Z��?D(B���6�8��n���%����C?
G�>0o�>/#�>۷)�/�g�A��:>�Q�>��Q?�$�>�JP?�|{?�[?�S>cp8�����ƙ�p:�> ">0�@?{Ӂ?�?�	y?���>�e>K�+�ǿ�6��4R$��'���#W=�7[>�?�>���>bǩ>Rl�=�Ƚj���z>�]�=͘d>*
�>-h�>d��>�@v>
��<RY=?䮚>ʞ���"��q�L���c>m�h?4��?�*B?���������b�;��=값?�_�?b�7?W�ܽ�J�=�(�����1DǾX��>�ո>�>�O<���=�An�Ǒc>�s<>Ç��wD�!!�m"�N?7�0?C��%'̿�q�
+o�� �����<����R�k���x��"M��ڳ=^���xZ�򷘾�wY��y���蔾���Jw����΍ ?��v=5��=�%�=��<�Jüiz�</4d=��k<�}=zt��6Z<D�Y�2��,����Q���;�JE=US<+Z��OM�?��l?��?{8O?��r>���=�h�-~>�P=��&?��>ל�=2����v(��7ʾ%.��~Ծ�|þ��a��Qx>3�w���>G�K>!��=�,D=�C�=h��=hfI=����i����M<tr6=��=w>�i>��M>�~q?Ӛ������XJw�p_i>Mq�?��F>�=pw۾�.M?{�>�5b������D��?q��?��?���>�}���R>�'����(>Y{=#wQ<�>��=�d���>YY�>���ܫ�����?���?�8@?����6�ۿ��=a8>2S>0�R�?1���Z���`���X��:!?�:���˾;��>��=�߾��ž[v/=t#7>{Yg={��"\�zy�=I�~�C�;=I@h=�ڈ>(�C>"�=		��&F�=ޜB=£�=]�N>?���
2�sK'���4=��=��a>m$>��>�??�R?���>�6=���޾�v�ݵy>��=>���b�.>9��>b�%?�L?g�Y?/��>���Z�>G޹>M�9�g/k����VY���3>���?շ�?��>³���+�� ��\�[�{��8?�H?��/?;�u>����4޿� �"�*�ԯh�?tּZa='Z��o	�L�&�3#�C���%�>T��>pҺ>oi�>O"|>D�!>(��=���>��>7,�<��e=Q5<;��<^�\�2��=� ���s�<EK��n ��s��G��'�	��;��;��� <�=d >=��>AX>r��>K�=t��EE->����R�v}�R�����u�a�:���-�	�I�~oH>�b�>z����|��u��>�x4>�ǎ>!G�?٥\?�)R>d	d��\� ���۞�Z�����E=z~=_���^/��*W�H�-��H����>�y�>���>/@�>0!��9�I�u=��޾��8��2�>�Ή�C�<2�*���t��4��C���(^��ZS=��C?	����=��t?�oO?�:�?�]�>;�#���X��=8��I�޼8f�o�p�Q���� ?ǜ ?�Q�>DҾ;+I�Цվl+��
%>��<=��z�A����2��/>~o�����>y]���0P�����ۊ�����w`�.$���H�>mI?W\�?X�@��Ht�����~@=�#?Z?DG�>na�>-9?�G����WV�$�p�-4�?���?��?w)�>SԽ=ﳽf7�>/b	?���?�g�?/ s?��@�z��>)���&>L������=��	>9	�=r|�=�_?F�
?f�
?�ߝ�p�	�t񾴍�K^��~�<K��=��>�8�>�q>�:�=7�^=��=�<[>�>�>zU�>�Rd>� �>W��>8��0a	��[?��=�>LJ5?l N>���<V�z�=��u�����xG�ϕ�������<�'���8�Ж�����>��¿Zf�?h->qE�sY? C��X��ݒc>4U#>u�1�d(�>n�>�\H>���>/}�>�)>� �>��9>52��j�>4b��V��XC�jXe��5��P�>f����%'�W���x���p���3־HP
��t�m���Z2�����㔘?�a�`j����_�%��1�>�"�>�3?�#���8�r��=���>��q>�<��W���43���Hξy�?�T�?@>�N>�[E?�?�?��9�0�m�u8��Y�Y��$|�qc��򙃿O�y� |��?>���bH?�N?Y?�p���bt>g?�v+���f�8�>��&�d���R��*J�>
�������찾�/>�U�4�F^>�v?s\�?��?l�\�񌃽q7.>�m<?�0?d�t?n1?0v:?-��l$?��7>(?��?�6?��.?Z:
?"�,>@��=w�û��(=�����$нi�ɽ�F�D):=�5}=�{�:� �;38=�G�<u��0{�?�*�Bʬ�Hյ<� B=t��=f��=(x�>-q[?��>���>/�2?zV�c�4�iE���,?�J=�󉾮R��G硾���'�=��h?z�?��\?��\>j�@�VH��� >,9�>��>a�S>H��>�ܽ�D��
s=ۖ>�U">���=ɞ�������;I���t�<�V&>���>~v>>��5k�>�6�����Q>���nS龪q��<b8�c �|<R���?�V?c�?�/��O���/W>-w�|\?�U?Yu?��P?�%>��㾈�=��;M��Zk�P4�>�o��
\<��������003�<"�=�FE>� ;Tݠ��Wb>$��h޾k�n��J�W��`?M=	���V=��־�9� ��=�
>����� �A��yת��+J?�aj=qm��	WU�q��	�>S��>]֮>�:�'3w�o�@������,�=���>~�:>�|��"�{G��7���>^�G?�l_?�v�?�Z��C�p�>C�~� �����#ϼ��?�]�>��
?4�D>Oy�=�d��e�o�d��CH��$�>���>�U�\4H�mɛ�o��i[$�@�>|M?��">�C?�P?w�?z�`?J�*?"U?�Ԑ>���	۽��A&?e��?��=(�ԽڳT�� 9��F����>�})?[�B�ݲ�>��?��?��&?�Q?$�?��>�� ��@@����>mS�>}�W��b��`�_>­J?H��>�=Y?^ԃ?c�=>�~5��ꢾ�ʩ�>C�=�>��2?H7#?]�?*��>P��>v�����=��>~c?�,�?��o?x�=�?�2>���>�i�=cm�>���>�?;^O?I�s?�J?�{�>���<����D���*s�v�O��;�wI<�}y=t��m�t�s�Ֆ�<;|�;�۵�3�y���'�E���&��;y#�>wgo> 뒾V�:>/���U����7>������s$���\5���=F}>t� ?��>+u#�(��=F�>x��>E���}(?7?e?��<a`�d�۾XzZ��C�>W�>?�ǵ=�k�U�����s��|}="�k?��]?�DK�]���8�b?��]?�g�=� �þ۷b���龟�O?;�
?�G���>��~?D�q?��>��e�:n����Cb���j�Ѷ=�r�>�W���d�l@�>g�7?	N�><�b>%�=�u۾%�w�Wq��,?l�?�?���?�**>7�n�"4��y��� ���]?���>��"?����ϾΟ�����c�ᾆ�����WL��Ux����$��ȃ���ֽ㊼=b�?��r?�<q?�_?�� �f�c��$^�O���/V�W0�m(�3�E��E��C��n��g����%���LG=�~��@��G�?�L(?�0���>����5B�K1ϾOj@>$���J�X'�=K���"68=�4U=��g�^�,�Z��q�?PE�>S1�>�<?�=[�yX=��1�p*8�\t��s	0>�w�>6`�>)��>� {:8�-�w��ɾ|����ѽ1�i>��g?L L?�n?�K	�u�-�����28#����&��?�V>"m>�Ԕ>Q�K�����7)���A���r�p��u������؁=�),?5�>ש�>	b�?3?�1��t��@�q���/�=��<ݛ�>�i?���>u��>R7ܽU�#��½>��p?�P�>���>����Ɋ��y�4����A�>�O�>B�?��>�+�|�R�5�������&�;�5]
>W�`?d���|�$��}>�TK?��,�c�痒>g��M<��W�LN��9�O>�?�֦=��>��Ѿt���z�����(?��>�־�� ��>b�.?k�?$� ?҉?�!>�����t+<��1?r�z?)��?NZF?��=2�c���=G罀Y"��a�<�3�>��>����x��D�Y=O�Ⱦ��ͽt ;�8�v><I����5��P:���!�f�D">KDῒ�9��W��꾶����N��Ҧ����ZI��P��;I��GZ��,vC��D@�|���ʪ���̀��$��N
����?L+�?l$��&_�7���k��|��>e�:�˼���̾0`$�c���L�ؾv餾��+��U���]��G�P�'?�����ǿ򰡿�:ܾ3! ?�A ?8�y?��6�"���8�� >]C�<-����뾭����οA�����^?���>��/��n��>ݥ�>�X>�Hq>����螾n1�<��?7�-?��>Ȏr�1�ɿb����¤<���?0�@�XA?5�(�[��*�a=�,�>~?��>>'.�k������s�>�-�?c��?n�==�4W��N���d?��^<�>E�X�޻z�= Ơ=ܘ=����O>�ה>���T�B�$߽\�4>��>d�%�����[�%W�<Va>m@ҽ�M����?��b�k�R�Z)#�����
����U?�S	?�q	�LR)?�6��'׿yuI�,g?$��?���?��(?�P����H>��ʾ�`Y?��W?J0�>5���{�&>���� =w"^��w�=&�?�Ԟ>^�F�e��r���D���V>����ƿ�$�mR��=����]��=轪���M�S��
��Gfo����T�f=���=��P>3�>�V>��Y>-�W?� l?�?�>�>��L]���GξS)� %����� q�I0���M�~߾�	��������ɾ4=���=�2R�򗐿	� �r�b�Z�F�I�.?�$>��ʾ��M�)�+<�rʾ»��7a��Q���v̾&�1��n�<̟?l�A?���a�V����Y@�½��̤W?�R�s���款f��=���
=�.�>Et�=���� 3�7zS��\0?�<?6鼾>䌾.>��� ~�<�",?��?�l8<3`�>��%?�z,��潦!X>�80>բ>FA�>�>X��7�Խb�?u�T?T��΃���b�>(H���}��9R=[��=j_5��t�� Y>YU�<7Ë��7-�b���v�<$pO?�V;>\�����پ�
��&�=�g�?��?W��>���?t@?/=�����e�)��A�~=�LL?bf?>� >�R9�^Dt������??�B?�ٴ=�E��.�ľ�fX��/���_?�S_?Zu?-)��{R�"�����p7?�i?��s�yZ���eA����g?ɒ�>%�>�W,�ҷ<f�\?Ҕ��b���gF��~*�=��?��@�E�?5���j��=���>��>�%��`ﾱ����ѻ���޽P?����܁��5/C�YG���F?�{�?�}?E��&�#��c�=�E�-��?3C�?�奾�Lr=�?�_3j�*��,鱼���=�F�Js��R�澳#5��ܾ1�	�%�����f<(�h>��@� �8��> We�3�ԿTȿ:&��9.��&�e��(?]��>�p��ë��Ks��ل���Z��gG�����9�>��=�l ��]��`�m6�SF>��?�:6<تu>��޽�敾Q����dԼ@<x> �>~[�>^�<&;���)�?��9�¿���R����V?@A�?>�?$
P?PX�>q$���8�ʜ�=�>?�|I?wv?�O�=�u�������j?�o���C`��4�SeE��T>(!3?x�>.s-��׀=w�><��>$]>�$/��Ŀ5ն� ����?{�?�U꾓��>�~�?�~+?�M��3���k���*����@?��2>�f��V�!�$=��֒�g�
?;U0?&'�a�C�V?r(N�ah��<��c��>qR�=�{\��z>�}�5�V�h���霾h�?}� @���?�S��#;���?��>d����4��/�=�+�>/$�>�Q>��+=�S>�0쾖a'�Q��>��?K*�?��?�X��mɧ���w=2o�?�1�><�?M10>��?��=B�Ⱦ�˽�(>��">v|���7?w�U?���>�.�=h�W�Go5�6mE��?���E8��ˎ>ƶV?l�E?	�>�P���z����*����Q[7��zｼx;�J@��������{>i�E>�!(>��E4��%?E++�55տ⚿�뾾L$?J��>�?
揾���}�9>�o?f�G>M9E�()���s�l�D�?�;�?��>NB�۪ݽ��ټ��	?��(?��7>���H��֠��|HL?�����M���@���>L.�?���?��?h|�}�?����&��נ��\����ŽIJ-> 9?R��f,>�?�>��g�~}���:s��٫>BS�?
��?��>^?��q���8��`��h=�>�&{?v?��"�BI���s�=
�?�j��Ĉ����sc?+�@�~@��]?�����߿	T��q`��1i��H1�=
�O=��>�����=�SI=N鍻 K!=��6>�[�>�R>��A>e�3>4i)>�u&>�����$����8���&9�*���<�P�J�����.~�ӫ��F������S�Oɩ�R��b{O�v+�G �S��J�?!�v?aR?���>�=�Yὅ�!��.E=��!��c�>:Q�>��u?rU?G=?��T�P	��Zx�eq��vŹ�Lj���/	?A�=��?���>�H�>�wK<�>֧g>qG�=���=�g�����d�=$��>�C�>���>�r�>�C<>�>Bϴ��1��E�h��
w�G̽5�?^���N�J��1���9�������i�=^b.?J|>���?пQ����2H?���o)���+���>^�0?�cW?�>`����T�7:>&���j�/`>�+ �Tl���)�j%Q>ml?N�f>čt>�x3��!8�q�P��r����|>;6?F���8���u���H��BݾRM>7��>=�$W�
閿��~���i��i{=�|:?ͦ?�#��Ԥ����u�އ��bQ>b�[>#.=�ͫ=e�L>��b�3�ǽDH��-=^R�=��^>�y?2��=s��=F:�>��Y�Ͼw�>��>��O>��3?�I4?XH�=���.W������i�>T��>��>s>�,�-�>(�>Qr�>��>�xl��jR��n�g�>ف�䮐���������K�/�L>��=�b㽨����&=E~?����ሿ|��\��g�D?��?���=l/�<c"�K���8��>��?`�@�ٚ?����V���?�4�?q���8�=0^�>(�>�̾��M�ݗ?}���+���	��v$�O?�?�%�?��6�`O��e�k�J>�$?�IҾ�7�>��'�����r��^�������k>kLE?ëȾ����U-�-j?���>���-u��˿�2p���>�>�?c��?!�o��V����E���>ig�?�c?�5M>Iɫ�-k�<��>��<?�Y7??Sl>����S���?���?5G�?��=ڡ?��m?g�
?�`?��<������V���w3>x����.�>�6�>�.�-="�����ڗ�����{��"�=Ah�e3�>�WV�/L���r�<�r����U��)��>܊>��>���>B>/?FB�>z��>�QT=�-�e�ϾW���K?�?>���$n����<���=۔^��C?DE4?�^�S�Ͼۨ>��\?�ŀ?
[?��>���A��T̿�Wx���͗<�K>!`�>V�>�Љ�
	K>�վ`�D�.��>6Η>�ͣ�L{ھ����請�E�>Vp!?�k�>}®=t ?s?�w_>��> qK��k��3�<�d��>���>�5?T�?[�?�+���G3�v��<��a�T�w�Y>��v?�Y?�͎>�i���Օ��;�����[�����?0�b?0� ���?5�?��>?�A?�`Z>�a�\�۾�S��Nb�>�#?(���5��,�����b~?|�?J
�>��>�D2�������/�^;���$?��s?D�<?��۾Y6a��0���t<�r��m�%��=M�8�S$>�D'>�k���Q<��>Fظ=/�$��B��=�Ę>���>!鬽=��2�r;�2,?�R�[>@�=��r��D��3�>��L>�}���I_?J^<�+�{��⬿�i���QV���?�v�?Mb�?�)��
Yh��<?q�?e?l��>�ů���޾�6߾�v�Sy�ذ�q�>o�>K^W���Rj������W\���Ľ62�}��>���>�=?��>�cD>��>l�����G���ɾC��c�\����Bo5���)���1K��A�ڞ���������S�>(\]�B�S>��?��6>_>�Z�>�5׽���>�Ua>X�I>
Yc>c�=��p=/��<�G�<V����Q?�b��E(��[��S���QA?�\c?�
�>;�Q����c;�}#?�?샜?�)�>�Je���,�<�?���>e��X�	?�X:=`�a��[�<�C��C���슽)�J��ߏ>m�ս�T8��NN��fe��Y?��?:=��̾u2ֽ�>����=��?N�)?��(�smO�� o�}W���R�æ*���g�z�����$��[o�@R���B������f�&�*s<=�(?�?�S����Fu���!i���>���a>Ÿ�>� �>s_�>8Q>�� 2�c_�fN*�r
����>��x?-\�>v�I?O�;? �P?j�L?Zm�>���>|N���J�>�Զ;4�>ah�>`A9?�.?5K0?_?H/+?o�b>�������>r׾~$?�]?�?W�?�{?�(Ľ`��$�h���y��(��#|=�<ڽ�o��]=��S>:Y?g��`�8�M���N?k>�q7?�}�>���>L現�?�� W�<��>�
?�T�>?���sbr�h�84�>���?���0=��)>��=�O���o��6�=�濼5+�=Ղ���;�:K"<�{�=���=��s��=k���:��;X��<Cz?U��>I�=���<4��+����g�Ү�w0>�6?�+�<����ۊ��ۧ��l���5> ݉?X��?w~=7w�=��!��o��Q����)�N(��>nn-?�,?H�z?�N�?�J-?��?s�=r��#����������c�?N!,?���>����ʾC�2�3�C�?V]?�:a�̲�9)���¾y�Խү>�[/��.~����"D�G>�����Iy�����?-��?��@�m�6�7z������[���C?� �>�Y�>��>��)���g��#�0;>[��>�R?Ԛ�> �P?֐y?N�^?/�U>��8�G^��T?��A*����>J@?B��?���?h�p?�{�>���=��=���־w���	�>����(O��y��<�f_>ݓ>���>�Ο>y�s=~�˽l߰��"A����=�d>���>�ܦ>��>m�q>�tW��<?�v>.��:4��J���hM��I�=�wM?kU�?��>?,���u&� .�����D�6>o��?n�?В/?֛m�)��=��ȼ�C۾�ݾMBc>=D�>�c>��>��>�L>�O>�bC>O�r��	�ڴ3�EzP=F�?��&?�P�;%ƿ�xq���o��\����<u?���f�S)��zZ��+�=Y���������b}\�:x��v����~��B���]xx�#�>ߢ�=�-�=���=���<8T�����<��H= C�<b�=1�p��`<��?�Q5󻨊��ȭ���h<��K=�I���%��m�?["�?���>�y?��>���>�T��uF>���=��?>���>&펽��v�d�f��;(���ƾs j��(���>W�"��TN>�>$�b>Ћ�=$[ػJ5�<����'�7o
��c=܂�<�e�=w�&>�A>�x�>�i?����s����o�vѽ��"?��A> �->����pr�>l�=�ב��6����ܾ��Z?��?B�?�T�>����>���3/>3��>+4��F��99>��%=U�V>�$>�|�2;���,���?=��?�E+?4a��<�˿%��=��7>A>��R��01��{\�f�b��3Z���!?Xz;�P�˾��>��=�V߾��ƾ�Q,=>G6>��a=QH�a`\���=i�|���<=,vl=�p�>��D>���=����%�=4�F=���=�O>�٠�޺8���,���2=��=�Kb>�=%>c��>ݏ?��?ԭ_?���>��u�����ʾXJ%>�`���K>���=b�=��>N�$?�F3?�JH?J:�>�&=ƨ>?��>��,���{�(
��79�L(^>�i�?P��?��>�¿=3YS���e�F��4l��M?��6?��?�T�>��HLٿt'"�5%�R��=H�Y&:�u#�Ļ�<W^�~%ݽտ�=��>�S�>�ӥ>'Rq>��->*��=�۝>
#�>���=������=z�=�i��ܤ�TH�=�:�L_=���;�+��㽽����[�2�:I=��:i:|�=�+�=|�>��>���>+S=�����.>�S����_�n�%>�Ʀ���K��\���x���.��p+���C>ېH>RO����]5�>+�M>-9=>%˰?�q?��>����u����[����1;�\�==��<ZAn�(?�o0j�A�I�Y������>5�>��>�{y>�?)���E��L=%�ƾ�G-����>�o��� �~i�hn��)��-����(d��9�;*�G?�ӄ����=N�}?bP?�a�? 	�>c�ͽ���S�,>���6���,.�����m����?��$?1s�>jR޾��>���Ⱦ��ý3��>�M�BUR�v ��%�1�����lt��u�>؝��_�˾�+2��Z��B��t\D��4u�\9�>�PR?u�?bh�b��;�O��!�{Er��?��e?�D�>��?S�?cP��+��e��<��=_o?���?���?�>�/�=٨���>��
?�!�?͎?O�p?�J9�j��>�h�t|!>�����4�=�>��=x��=�?6�?��
?s���i
�MO��$��yg��-=J��=�O�>���>"8t>���=��@=n	�=m�\>�ӝ>���>c�j>�f�>N��>fȞ�7����&?�@>�S>1?L�v>Ï�<�}�}Gu<�I̽%0��r�R�}��v+�E!;z��{�=��`b�>�[ſ���?N�o>�V��-a?i"��i���L>���=KN=����>!�<>��>S��>�,�>�c;>���>�{G>�ᾞ1�=���o�	�w]Y���b�t����>|������^�$6��%ž����&�����=P0�/��=´�?��E��8����>��᾽�>`0\>�*>?�}�����1>��?�/b>�����������."ƾ|ۃ?g�@��i>��>ZXE?�)?��ǽ�'���x���2��lv�"v�����K���4r��F�A���Y?��b?�4?��[��Y�>�S?Z�A��w�|��>���T�>�Ch�v?�N��D�����M��s��u��PC�>Xzn?Ↄ?/�?>�)��1����4>�@?��-?mHw?��3?�4<?Il��!?r�9>Ǟ?t�
?K�7?��.?d	?�@%>T��=(5��� #=!���3\��x<ɽj׽�ü��@=�_�=L?�;��n;w@&=�Ny<�4���{/�:�����S�<~{U=���=+�=�)�>0eY?�c�>r�>9�8?��:�j6�^짾{!?�i�<h�Da������[�����=�3]?�0�?��Y?��>��>�{#��>�}l>2>_5k>&3�>$����K�-1=�3>Z�>	�K=�,½����HB��D��8�{=��>���>y!R>=fw�K�?���=yx@��X>Np��������|�b��U2���&?3+Y?Ƕ1??U=�� ����=�V�&R�?��J?U�M?b=?�}R>�J־�`_�=�U� ��%yg>}�h� y�󷑿z��-S9�ɲ/>��>���ゞ�it`>�J���ھm�+�J����Æ
=�����==֑��Yھ=傾|5�==>ͤ���W����7�����I?zHf=����4[�σ���f>%�>��>1�d�A�$O��A��=���>xy6>�>�R��>G��g��N�>��H?�`?�{�?KH��b~p���E����?���ȇ��Z?�ή>z�	?`J>���=����:��e�"UJ�R��>��>,3�D�G�!��0���!��N�>��?(>��?d�R?�?!nb?U�+?�?�ː>H���𕹾�A&?���?i�=1�Խ��T�~9�5F����>�})?L�B�7��>��?Ÿ?��&?�Q?�?��>Z� ��B@�ʖ�>Y�>E�W��b��*�_>��J?x��>V?Y?�Ճ?�=>�5�7墾�ϩ�,8�=�>��2?�5#?�?)��>4��>C���K �=���>�
c?%0�?��o?$��=^�?392>��>�=5��>i��>�?XXO?N�s??�J?���>���<�3���9���;s�H�O���;{DH<��y=��HGt�y:����<̢�;�<��m��}��x�D�0����;�>g�h>cp����2>����Ϗ���L>�Ë<|M�����FeN��=�܂>�`?��>�C�yCR=�w�>'�>4��N�+?>h?�?xi<A�a�Uھ^O����>�B?�x�=?�h�.哿j�q��z5=k?N�^?�#S�H���J�b?�]?0h��=��þw�b�ĉ�_�O?>�
?#�G� �>��~?f�q?Z��>
�e�.:n�*��Db��j�Ѷ=`r�>IX�R�d��?�>m�7?�N�>)�b> %�=iu۾�w��q��i?��?�?���?+*>��n�V4��f�)�����Z?]�>&���r?�*���о���ۿ��*#վ�N���5������`b���)��u��l��k�='�?h�v?�s?��g?\;���a���_��A{�E`Q�ט���MJ��LD���D��&h���������>���Q$=F�g�o�>����?�*?�	7���>骔�X?�on�i�I>�!���1���^=����W�<_2/=�%g���8��=¾TK?�o�>���>�:?�W�(�:�G�(�.`5�D+��E,>w�>"S�>��>�w<v,����\��6i\�ǻ����u>��c?s�K?�n?£��0�!���ŭ!�0�0���n�C>��>�ω>�GW�����T&�-j>��r��#�F�����	����=�v2?�.�>���>09�?G�?�f	��:��V�w�~:1�#2�<,��>�i?:�>�ǆ>I�нS� �&��>6H|?��>�@�>Q���>��������+��>� �>��>�L>ˬ��0T��֏�b��l�G�{��=�`\?*����q��>�I?v
&�4"<jkS>��߽A����u���$=�0d>bc?�m�=�x�=���N�\~�\���,?�?������"����>��,?�U�>���>O��?��>t��ن�%?��n?.�]?^�>?�ت>J������aSƽ3�"�d��<��>zw<>��=/�=Δ���S�`9R��L��m�=yf��{ʋ���<T�~��:J��|�<�R>Uҿbi:����������� ��]
������i��,^��2�4�(����֮�;~������6]��g��ƞ�������ų�G�?���?�0��Kh3=+��;[|�Hw!����>�I�Ay��w��-DQ�؝/�g뾦e���5�F�Z��N��_:�O�'?�����ǿ�9;ܾ! ?�A ?<�y?��A�"���8��� >�E�<�/���뾵����ο?����^?���>��'0�����>⥂>h�X>#Iq>���b螾q-�<��?E�-?��>�r�-�ɿO���R¤<���?-�@uA?�w(����|�]=�7�>��?�@>5]2�&h��?���q�>�?��? �<=�\W����e?��h<��F��B ���=�?�=̏!=��^G>"��>���BF����]2>"!�>�0���x"[�/��<0�Y>FRѽ�o��h��?�t_�~zU�Ȃ��\�@��d�3?:�?j����#?4�#��RֿQ�\�V�\?��?���?��3?�2�#>aZ��j�.?��F??�>'�H�)&���>(>U�@�`z]�KҾ3o��I:��1?�_�>��~����#���q�=j0y>o� �=¿)��>� �ȥ�<�{»Vx�������SL�>�e��L�3齞��<Z�h=��=>��>T@:>0�>ӈY?�s?ta�>�Nu>1��6�����׾Wy#��s�C.%�Vॾ'.{����A.��n�ӾZW����)��Ͼ��<����=I�Q������ �plb��xF���.?׻&>jfʾ��M�~�< ʾ�u��Z��W���˾*G1�on�l��?�B?ㅿ��V�b����a�THW?����<�*#�����=v����=�5�>�&�=�|��T3��S�ܾ4?�8
?�ӓ�n����04>kY���c=�7 ?f"?�c�1�>s2 ?�q��X�O��=�Y>�>�?I!�=z��Z{����+?8uf?��
����u>m�ƾl�꾎b�	\>�0���{MT>/>�ķ�������+p4=��V?<�>~~'�Ҏ�⊾����=wy?�9?��>�b?�u4?\�<y7쾭�R�:���>��=��S?A ]?6>�ϼ`�Ͼ����8?�c?�<>Mp�=���.:��L�)0?�	_?�M"?ԋ=I�u�v�����01?�&p?P�c�(���^-�1�F�q�?���>�L�>[,��x%>g�J?�����ę�4���4)�C��?�@���?wh3���2��>=W��>��>_�<�����u��b =;?�ƾ������%��9���U?�?�W�>ϯ��e$�Ʊ�=��{�i��?!d�?�f���w<B}�n�d�����[��;��g=p{R����˿�T7��վ.�����{��!y>)$@OQȽ.��>LsJ���ۿ�@ο�3���s��8GQ��?���>����Ҧ���q��{���O��G�&荾A��>� �=ws��/���hw�0}X��0�=O�>@MZ���X>�~)�uA���Ⱦr�ٽ�a>B��>ey�>Ф5=�յ��l�??S ��Pɿ�Ȧ�(G3�<<?h��?�ܓ?��m?��>���z8Ծ�I�>NTI?�:?�fb?x�3=߯��n��=$�j?�_��tU`��4�tHE��U>�"3?�B�>S�-�P�|=�>���>g>�#/�x�Ŀ�ٶ�5���Z��?��?�o���>q��?ts+?�i�8���[����*�?�+��<A?�2>���I�!�B0=�RҒ���
?Q~0?{�f.��j_?]C��d�]x��-�=>��>�s%���$���>
�H<g,�����   �+,�?z @Vέ?�Q���?�W�?z�>T]�+`��*E>F��>�I ?d}�>� Z=x�S>�f���<���>!%�?���?p^!?����"奔e��<nlj?�}�>�`�?<��=k��>���=#g����`�q�!>{�=�8=�S?гM?E��>���=5�9��/��F��7R��@���C�_�>��a?��K? c>�ĸ�W*0�� �r˽�0��=ۼ�=��*�;�޽�m5>ɱ>>��>k�E�k�Ҿ~)(?�L!�HRܿ�)��](Ⱦ�.?0]n>η?n���"2��><�?$��>�D�$i凿���?�?s^�?���>إ��jS�2�����>�,?�0�=[������^�=��Y?��#���-A]����>�h�?�D	@��?�����?�$��q������[���c=��>�.;?<Uܾ�Wp=�?pC>Ȏh����r� �>�L�?�E�?XF�>��T?t��/,�8��	B�>�E}?�/�>� 佹p
��D@>=6	?�5%�2����̾�n?da	@C�@oy_?�f����ٿh����Ⱦ��Ӿ^�s<,��<ss�>�U��r>�i>gC�6��=�#{>}}�>��>KU�=j�9>,�7> A�=.-���)&�j�����kRN���
�خ쾻NY��⾪,m�������������xb1�;t���i��B�T��g�轁�<���?�qr?w<n?Jq�>-���m$�;��4�>�Z��fA�>��>��F?6�S?kO?�:f�*�龰�l��g~��ٺ�'ք��q�>B#6=�v?��>���>��5=i'">S*j>U�=b�= h�n�=���=o�>C�>���>	%�>TE<>�>	ϴ��1��Λh�:
w�P̽	�?v���J��1��G;��馷��l�=}b.?�~>j���>п����22H?r���p)�շ+�D�>�0?�cW?L�>���(�T��:>���צj��b>�% �V}l���)��!Q>�l?p�h>C�r>��3�3�7��O��v����~>�k7?%(��|�9��v�E�G��۾�P>�>�- �����薿��}���h��/�=O~:?  ?�:��\�����u�z��eM>T�^>j�=�:�=�I>�0c�A9ʽ}GF�1�8=��=Yz\>��?��$>D-�=l�>IV��3H�hP�>}L>lL>�'>?g?��B���ǅ�d=��v�>�y�>_��>���=%�@�@��=��>�Wd>?ʟ�� _�|�+�dO?���?>�/̽�aG�Ɉ���B=|zP��O>��=s��W:L�1l=Ħw?<ŕ��ل��`߾L�<~)R?O- ?>�j>vS>g�)�����'վ�R�?YB@­�?��Ѿ�g���>J�?�i���Aq���v>lN�>���d�޾I��>"»uX��_"�������?�y?Oef��
}���N����=��?#������>�n�G���~T��В�����7>��T?�E����=��$�0�)?��?f��:���̿��z��d�>!�?HD�?Ln�R`��I�f���>9:�?�k?t�$>��s�;�����>�R?[�*?.�\>��,�j���#?���?�*�?�>�ʣ?��?f2?�tg�,��+q��Dρ��>��=ҏ ?7R>�,b�ߦ"�������@������W�o<c]����>�ۼ]����Au=zv�������F�uQ�>���>Y�>F��>�?�??��>3��=������E�]�K?r��?j��"-n����<�r�=��^��/?�I4?��[�D�ϾSԨ>l�\?�?�	[?Kh�>����=���῿E{����<��K>�<�>�K�>�B��k;K>.�ԾPD��w�>]ӗ>壼�Dھ�)�������B�>Ug!?h��>)��=�� ?�#?��j>H6�>'aE�A6����E�e��>���>�A?P�~?��?͹��X3����&衿o�[��?N>O�x?bO?ѕ>W������ɼF�.'I��/��ۗ�?�vg?��?�1�?
�??0�A?��e>���ؾѭ�N�>j�(?w��CWB�g~!�g̵�̼�>�>ҙ?���=}X��ީ��+���;.H ?bWn?�j0?\��'�`��ㇾ@M�<���v�0��Z�=�x�<L!�=�
I>Z�����$�B>�=�Z&�7B�L�=���>l �>0ֽ������{�-?�����`�=7�c��:��>	NA>2��HZK?�5��f�����/m���Co����?��?}��?$ؽkEa�b�2?n��?;�?j�>D׹�<�־���MQ��n0��!F�D>B��>�@���D������F��D9y��Jƽ�HG�>H|?z�"?U��> ��>j5Z>�ǚ��<_�$���"���\����;@2�J� ���	�������C��7����Y��i��>�{;V�>S��>[�d>q#�>��>���= (�>��'>cWx>�.�>�đ�	���߿ =Ƿ:=��&�v�Q?o;ľ^G+�rG⾡8���9?�e?�Y? ���ț��9��|�?���?<��?��>��]���0���> �?`	{��G?k�5=ș<]��<h�˾�����2�/���큓>޽-���N��}���?Sc?~+ֻ/�þn��ύ���R�=)˄?kN-?�#)�Q�L��}m��R��QQ��,J��L{�9ɤ�!� �m��A���;��0&����"�r�L=]�$?{Ј?������������d���A�EO^>���>M��>Px�>0R>�6���0�(~c�B�-��Д�,�>eqt?t��>S�I?|�;?��P?�mL?W��>�R�>1���#�>���;y��>���>4�9?�-?�>0?#a?da+?�.c>,�����*Nؾ�?�?u ?�?�?KŅ�
�ý�Й��zj���y�b遽���=Q<�<ߥؽ��t���V=�
T>�^?Ƥ�	�8������[k>È7?���>�>ɏ��-��>�<$��>��
?���>�t���Vr�x����>T��?��(c=r�)>��=�1�����DD�=}����=]�����<��f$<#|�=\֔=�{�S4�Q �:Hu�;!��<�B	?�o�>�l�>�c�>��C��^���ӾW��&>e���=����T��b���:QR�K��>p��?���?U���(�>~�=Ъ�P۸����(	��c?���;+?�U+?BeM?'�?��?�2?��6>=��Ʉ��o�Y�ᾏ��>{!,?���>���*�ʾ�憎R�3�ʝ?)^?{9a�c��9=)�ݏ¾��Խ��>�V/��+~�.���D��݄����g�����?���?�	A���6�0y�ھ���^����C?Z"�>Y�>��>K�)���g�*$��1;>���>�	R?���>��p?�v�?�rk?v >�$�[���?e����=��:>&u`?�)�?F%�?��|?r�>�B��}���7�������ٰ�"d�	b\�^c��>�֐>'I�> ��>*B�=��n�۽a락�+>�Ί>4��>�]�>y�>� B>`W=KD?�*~>�]���������b��?/�?��~?�jV?������t[�d)���g����?�ַ?�@Q?v�мe�>��S=f��礱���>QS	?Gy>"#>���>0��=�#�>T�>��|�Cƾww��`��@/?�0O?ٜ����Ŀ��q�!
h�Ѭ���;�;Qe���b�Yۗ��3c��Ƴ=/f�����9���Y�jʢ�l����rV������~��>�v�=��=i��=�&�<gO�ӆ�<��9=n0�<Zh=-�n�U�v<}vG�ί��p�ˆ�:�V�<�c=�����⾡��?5�f?H(?��\?�c�>��>!ν���>+(�=� ?Mm�>���=�K=����1÷�����X��lҾ^�p��Bھə�=�	���O>�BX>,�>>㨨=U��=�ma=�>���+ν�<��=oI�=C��=�$>��>W�6>��s?�6x��q��;�\�0�=;'d?�[(=hj>>�&��`e ?�ڑ>Ꝃ�5��0���\^�?.l�?#��?��>�<��R"�>�8�[�=�|>�j>��J콨��=��b=o%�>ⱬ>����棿B:ҽ.M�?5A�?
JC?����u��R\/>�8>'>1�R���1�T\��hb���Z���!?U�:��L̾� �>Sl�=6/߾)hƾ�n.=�7>��d=j,��G\�B�=Gz���:=^�l=�ۉ>=�C>��=߁��b��=�ZG=y��=�_O>z
����4�<�&��4=�h�=��a>�J&>ա�>��?$�?}W?JK�>T�lB��U��WM>�HS=V�>�����u�=Z�>�,?�iX?cJ?M{|>��=��>T&�>��l�w�4���|�S��>�	�?���?���>��a=I���3����N�I���z
?)�8?s1?���>u0
��\Ϳu�5� �]��]�������s=�ca�<(=)�1>�s��54i>�>�>��>�G=�ꀽ�N1�?>��>���>�a>b-f=q�=�Ln=B��<9׽ʟ=.�����?�@�J=T1a�
�t��}���
��:��=]���S$>�T�<�>���>?�(>+��>.�=�Ԭ��>󿟾Z�R��o=������<�C*g�?��in*��> �T�G>^)e>
i��#����>�z>FX>hN�?fcp?��>�C�՟�ѱ���TJ��D�y�{=���=��>�f|@�sb�0�D�#+���>���>��>��l>H,�j ?�Z�w=��Nc5�p��>�r��Ay��E��:q��<��󟿬	i�hU��j�D?�D����=�~?��I?&ߏ?}}�>�$����ؾ�0>�X��o�=H�;@q�с����?�'?�~�>_���D�"!ƾ�������>�H�5TO�7G����/�gռ�������>8Ǳ��$־�
4��ꅿ,�1�;�՞d��Ŷ>��N?xĭ?׬Z��~��sP����[/W�$�?�]i?I�>�]?,�	?)�_���s�����="�k?���?Ux�?s�>Sν=�W���3�>�	?�Ŗ?0��?uxs?��>�j��>��;ģ >bB��J��=�>�*�=��=v9?&[
?.�
?S���'�	�������O^���<�ء=�{�>�e�>��q>Y��=zh=q��=��[>���>���>��d>��>�v�>쬜�{1�fT,?�)>�"�>��3?J@q>��=1����<����Y�B�4��Nֽ���ð<�{���<�����9�>&ƿ4��?w%^>�R	���?�q�,h��"Z>W�\>Q�ν,�>��B>�H�>6B�>�Q�>H�>���>1>Aa���w>���\"޾��m��{i�>��t�>�ĕ�ۅ/�����U���l���ھ]s�L�u��ހ�MV3����=7J�?4��S��`8V�p:��Ν�>�"T>��C?�9�����q2>�y6?��>��ؾ�/���z��=MԾd�x?&{@�0�>�V_> CB?�5?|ԕ���2�'�f�m➿7a����U���j��h���҆�����BM�JR?Ob?�?���eSm>��]?��l�y���7q>"�:��C�ӏ��B�>H�˾Q�p����X+˾�@��0^�>�͊?�g?�U�>����zξ��>�	c?��>��?SA�>��5?3����>W��>L�?��?�N?�L.?���>�2�YD��H:Ž�No>~�|�F�辘�R�S�5��ݜ�;½`>k�=/t�xoI=�&=�����d9X�｛��A%=��7> �H>�j%>:�>(�A?߁?���>�:?��S�Q�X*��zs ?l>N��3T��|(������(�=j�T?��?�	�?\��=?~I�/w]�q>t�>��0>ј�=��>j|%�L6���2��>�V=x��=�Ǳ��Ӯ�W#�������a��=J�=�]?�Me>�{s�;� ?����?��&��=�!�ʄ
��?���儿J�'��ֽ��?��_?1?�}��\��kC+>�(J���}?�W?˖/?"�(?Ҹ>��ﾃwW�6`\�5�d� ��=K�=�I�;H��EJ���oM�Xe�=$О>����!���b>Ȟ�`޾�mn��0J����zO=*o��U=0���վ���:!�=�	>������ ���ֶ����J?p�k=������U�괺�4�>�>|Ϯ>͉=���w�{�@���g�=���>��;>h���g�B;G�.��9�>�8E?_?Є�?�?��,Qs���B�0���o���Լ��?��>/P?��B>xȯ=�������Ee��F����>���>:��G�G��&��$�$�#�>�=?�%>��?IQR?��
?K�_?�	*?�{?�W�>.8������ߍ?�-�?.��������ZaL�R(?���?wU�>'���쾛>�t�>��?�d?p\?�9?L�N>��l-����>��>ڊY�ͦ��z�>��h?0��>�q?\0�?,;�>t'��z��.J��zx�\)G>!q.?�??� ?��>>|��>L�����=ƞ�>�c?�0�?"�o?��=<�?�:2>N��>'��=���>c��>�?SXO?>�s?��J?��>R��<�7���8��#Ds���O��ǂ;]uH<��y=��3t��J�4��<��;�g��<I������D�;������;v��>�8>����!.�>t?P��iԾI�A>�@{�7# ��*��)O��ˣ=�Z�> �?���>��L����=�+�>e� ?���?W7?���>Q�?��H>�e��$�wI����_=b� ?.��>��c�߀���t�Ȳ�<�H�?\ew?[�߾���O�b?��]?@h��=��þz�b����g�O?=�
?3�G���>��~?f�q?U��>�e�+:n�*��Db���j�&Ѷ=\r�>LX�S�d��?�>o�7?�N�>/�b>'%�=iu۾�w��q��h?��?�?���?+*>��n�Z4�>���F쑿o]]?��>M���J�!?�o��!ξ	����� ��&��奬� ���a���n�$�`����׽���=�?πs?��p?�j_?� �-�c��]�����<V�I]�I��'�E�KCE�.�C�3n�;��1���1��oqK=�l,��G���?�'?"ꊾ���>�r;d��'����>�h��@���X>χ7�i �=f�v=���F�ս{t��ϩ#?�C#>惠>K�X?ԋ]�5=�<�0���5��X���,>�,�>N6�>�?�j�=�
�3<����t�����/�u>��c?�(L?��n?�K���0� �����!�>�*�m��ܮD><@
>�>�>��Z�R� ���&�A>�7>s�
��i�����	����=A3?}��>�>��?��?�o	�����ȿv��?1�΅<|��>$�h?A��>�X�>;�ҽ �ԫ�>e�??��>�vo�Ɂ�3U��#=K��� ?s�>��?��}>J���jx�Y���Hؑ��N���h�/�3?mM��e�Z�$8?&b~?�ؼ�'B��=�>�橽�P$��Ӿ����y��i.�>���=$�I>"��N}$�sk���X�
P)?�K?�蒾��*��4~>�$"?��>�-�>S1�?�*�>hqþ�LE�ұ?)�^?RBJ?lTA?@J�>�=� ��Y=Ƚ�&���,=��>]�Z>�m=�~�=m��#s\��w��D=*t�=��μ1P��2�<����Y�J<N��<��3>�ڿ�C���Ծ�B���C�y���5�D�[o|������g��,�������b��2V���Y����i�x�_:�?=B�?2B��f/~�<����~}�<������>4�~��}�������x�p����侺z�����tRD�im[�W�W�T�'?Һ���ǿ����;ܾ9! ?�A ?�y?��5�"�ے8�l� >G�<5'��^�뾠�����ο9�����^?���>��z/��}��>ƥ�>��X>�Hq>����螾/�<��?[�-?@��>��r� �ɿa���7��<���?+�@MhA?��.���ݾ�:�=���>k��>��>ɞZ�eI��׾�b>�>��?In�?��=v�N���ż:�O?�§=rD��"�:��>�!���z�<�	��M>�O�>e�t�)����j��(>0�l>ᡅ��ҽtK�L-¼��J>����rP<Մ?h{\��f�ڤ/�U���U>��T?@*�>+5�=��,?78H��}Ͽ�\��+a?�0�?Y��?��(?�ۿ�Bښ> �ܾֈM?mC6?W��><d&���t����=2[��������'V�m��=	��>F�>�,�����O�s3�����=y���¿��"���JL=Y��n|a���i�3����y�����E�R� � ��<?=ؿ=��N>�Á>�3C>�=>u�X?��q?���>�%>7��r|��\$Ҿ8_��D|�N�B�����7'�85���,�h�ݾ������Q{�ǉ���T=�8��=L�P��/�����ƻc��F���.?�,!>l�ʾ��L�p�F<�5;d'��@F�������Lʾx70���l�`��?*A?�����W�������c��ԙV?3�'[�@H��M��=Y��b=1@�>Ӏ�=�$޾�:1�:�P��W0?��?#�����r
*>�_��>�	=�L+?}�?~�s<�Q�>�p%?9�+�I�齏mW>��1>�ۣ>ڼ�>1�>7;��@�ڽ��?��T?���������>ƽ��I{��H_=�"	>Ι5�[�缗�[>T�<ہ���V���+�<j$W?s�>��)�������g����<=�x?�?p͟>�uk?�C?1�<�3����S���Nv=F�W?!i?Υ>����+о���)�5?C�e?^�O>o)g������.��R��?˘n?$b?eF����}�b��@��b�6?��v?�r^�vs�����.�V�=�>�[�>���>��9��k�>�>?�#��G�� ���}Y4�%Þ?��@���?��;< �f��=�;?c\�>��O��>ƾ�z�������q=�"�>���sev����R,�S�8?ՠ�?���>������Š�=�ٕ��Z�?��?o����?g<Y���l��n���~�<�Ϋ=H��D"������7���ƾ��
����ῼ���>>Z@[V�w*�>�C8�T6�TϿ!��\о�Sq���?;��>/�Ƚ����5�j�~Pu�L�G�.�H�֥��y��>h� >���l��N�����G���%=Fj?za׽o\;>�6g�:D��qӾ����X �>3��>�f�>�s9������?�����̿����'|��YT?��?�~?m&?t���I����۾��-1i? �?<fk?��={p� �="�j?�_��tU`��4�sHE��U>�"3?�B�>U�-���|=�>���>9g>�#/�m�Ŀ�ٶ�=���T��?��?�o�3��>p��?vs+?~i�8���[����*���+��<A?�2>���O�!�L0=�cҒ���
?N~0?{�h.��i^?�g�`@w���T���u�A�> �n��K��ݤ���f?u��޴���g�e��?c�?�K�?D���9�&���'?Ճ�>b��W����'����>8��>o�2>�AN�2�4>X��:�c��#>^u�?���?Ga�>x����p����C>�/�?T�>k�?7�=bY�>eC�=�߰��-3�]#>r��=!>�ԥ?ޗM?��>0E�="�9�t-/��KF��GR�����C�/��>7 b?�L?yAb>¹�gc2�� !���ͽZ`1�-���@���,��c߽05>�|=>�>�NE���Ҿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?y��P��a~�3��)7����=��7?�0�h�z>E��>+�="ov������s����>�B�?c{�?���>��l?��o���B���1=ZL�>��k?,t?4o���"�B>)�?}������`K�- f?�
@nu@��^?������;���F���.��w�G>;>��>a0�|g�=�>5�>��={��=lHa>3�7>�R`>`;O>a�>��pz� ��(���ۿ���I@�����R��
����O�o�6���K��D��	4��XC��{����G���V��E��=i�U?�R?p?�� ?��x�ؚ>����'=d�#�8=�,�>�g2?��L?ݢ*?ԓ=A�����d��_��6B���ȇ�k��>�pI>N~�>0K�>�"�>�]T9(�I>�4?>���>�� >�a'=u��c_=��N>%M�>���>hz�>�C<>��>Fϴ��1��i�h��
w�m̽2�?|���Q�J��1���9��֦���h�=Ib.?|>���?пe����2H?'���z)� �+���>��0?�cW?�>��C�T�/:><����j�3`>�+ �zl���)��%Q>tl?ѹf>	*u>A�3�Sf8���P��y��(w|>�+6?�EZ9���u�۴H�x^ݾ>JM>|��>3E��m�8���*�|i���{=y:?�?�K��.԰���u��>��l]R>�S\>ٶ=�X�=�OM>tc�I�ƽV	H�R.=	��=c�^>�V?  ,>j��=2ԣ>�Y���4P�/p�>KjB>:-,>@?8(%?nA���Ñ��.��w>�S�>�
�>�Y>�cJ���=u�>@�a>h�T��{����?�>`W>i$~�"V_��u�7�x=1�� ��=���=�� ��8=���%=��u?�o���{��5���ܬ�(}<?�/?���� �%��b���ؾa2�?Z�@���?L��U��?5{�?Ύ���e#>���>}��>�������(�?�=�Y���Y�/��F�?ғ�?�kE�:�u�a�f��=>#?ш�Sh�>�x��Z�������u�X�#=M��>�8H?�V���O�R>��v
?�?�^�ݩ����ȿ5|v����>T�?���?b�m��A���@����>8��?�gY?�oi>�g۾``Z����>̻@?�R?�>�9���'���?�޶?د�?z�>@G�?9��?z?�[��'
�񧘿�߁���C>=��>r��>&��=��׾��^�������?�o�7JH��>n<�:�]>΁�=#Z��͆=Qd=�~ٽ���<� �>��>�-n>i�>�h�>��>���>��=�Z-����UgO���K?���?-���2n�
O�<Z��=)�^��&?�I4?k[�|�Ͼ�ը>�\?j?�[?d�><��P>��G迿6~��H��<��K>&4�>�H�>�$���FK>��Ծ�4D�fp�>�ϗ>�����?ھ�,���S��GB�>�e!?���>�Ү=L� ?��#?��j>�/�>YeE��8���E���>H��>�B?U�~?� ?
ù�oU3�����䡿ߒ[�0PN>P�x?tT?̕>t�������0E��*I�:���k��?tg?���?�/�?<�??u�A?�,f>{���ؾ�������>?�!?#�ںA�N&���~?�P?���>�<��w�ս�eּL��/����?�(\?�@&?���+a���¾�1�<~�"�jaU���;T�D�f�>{�>���đ�=>}۰=TOm�fF6���f<�i�=��>Q�=�-7��w��&=,?��G�yۃ�K�=4�r��wD�y�>'IL>*����^?l=���{�����x���
U�� �?��?Uk�?����h��$=?�?Q	?�!�>lK���}޾��Pw��}x�$w�x�>���>��l���W���𙪿�F����Ž�r���?+�>�>�>��"?�$>؂�>4ޭ��4��s��U$�%�e�!T�3��b#�b��"�ľ� ����<pl˾�/g�r��>�н�P�>˕?Sˎ=�i>�N�>Gk>��>Q>��J>J\�>�S >��>���=졢<sY�$�N?Z��H��)�O����g�?]D�?lC?v ¼P�����\�&? S�?�:�?]��>i�P�q=��xG?�� ?�j���?p������3��>Y�����=c��=s콓N>�ʟ�PE2��_�Ё/�$�?��>1��=%
Ҿ��=����y
o=�L�?��(?;�)�y�Q�սo�<�W�^S�&���0h��f����$�1�p�쏿^���#����(�T]*=K�*?w�?����"��~%k��?�Z_f>��>n�>�׾>@nI>y�	���1�n ^��K'�3����R�>�Y{?���>I�I?'<?xP?�kL?I��>�c�>�3���l�>��;� �>5�>%�9?z�-?80?�z?�t+?�3c>�~������ؾ�
?\�?�J?�?�?Gޅ��sý�g��_g�`�y��~����=$�<��׽�Eu��T=G
T>�U?0����8������k>�}7?=��>���>����3��a�<1 �>�
?6H�>�����|r�%e�S�>��?���c=��)>X��=#����˺�)�=?�����=_f��;�ƃ<�y�=)�=��t��z�4��:��;�3�<-L?
�8?9�?>�ʗ=M��N��U�{h�	I�>_A�>�T�=`����兿c����8��c�S>���?�M�?7���(�=:6#>��>�zޣ�������mE�=-U?�~?B�9?'��?F;?��!?�=����u���!��p�ľ5?x!,?���>�����ʾ�񨿶�3��?5[?�<a�����;)���¾?�Խ~�>�[/�[/~����D�!Ņ�����}��!��?翝?�A�d�6��x�ǿ���[��B�C?I"�>^Y�>(�>~�)�t�g�Y%��1;>��>7R?��>1�?^�v?\�i?�F=�\6�r䭿j/���O�Be8>H�A?��?���?�br?��> �8>�j�M��d)���w���E�Ͷ�=1G>Wzv>w��>�C�>�ū=\X�����A��>�؃>zx�>Zώ>r�>Bӯ>wPl=V�B?�C?��� %�'�̽UlQ=GW7��v?��?�c5?�%@=2!��|X�w�
�P�>�^�?��?�'�>�,�[��=+��;ڙ��ʹ����>�[-?�F>E+s���>]<m>��p>e��>�^^�U�-��W}�����B? �}?G.���˿��i���w��s��Ҹ=#1����:����=�+��V>��$�A�������ea�.D���ȅ�0����� q��;?[;>��=S>
�G�R���
�'Q=:��:�6��5�Z��=�L�r�����n仇[*=s�#=�ځ<��žz}?��Y?�-?�z:?��>>)Wr��>�69;�?��]>������ž�_��=��"��KO�&�;	�a�G����
>~Ae�	>F<>���=�]�<
��=N��=1�=]԰;�,=Ր�=���=> �=-�=�w�=��=��r?�d|�@���W���3��F'?��>�Q>VHʾ�<3?��>i���?繿�~���ހ?!��?���?���>�V�w�>�qþ�m�T휼<����q>%��=��F��Z�>	N>��86���֙�tG�?�o@�2>?�Ń��ɿߕE>�7>#&>��R�>�1�g�\�;�b�;yZ�]�!?�I;��K̾�4�>���=,߾4�ƾ��.=��6>Xb=qh��U\���=�z�G�;= l=�։>�C>�l�=�0��e�=[�I=���=��O>:����7�)1,�_�3=���=��b>|&>��>̓?Xs?�s?p��>1��q�羵������=v���C��>��<�-C>f�>h=;?b�Q?�}K?�p>Ii�=z#�>K�>PF0�!n���о����x�;��?�~�?��>>�D=�d�d��*G���R�%r?��,?1��>]�K>���	�ֿ z�2��&�=8�T=U��=v�-�Dm!��	�='5�;0�;=D�=B��>;ץ>�:�>�fQ>jV>/.�<e1�>��>�*%���=�⮽P��p���> ��<,��;��{�{�O���`���M��cüϪ7=Ey=ۼ�51�<P�=\|�>��>l��>��=d��8�8>C���͹M���=۫���A��Ub���{��m-�k�7�cw<>��V>��j����}?�Y[>k=:>K�?�;t?�>�b
���Ӿ���D�e�u�\���=4>�A�#t:��_�p�L���վo��>�>���>��l>��+��!?�~�x=�⾻h5����>�������p��*q�7���🿽i���Ѻ=�D?�E��C�=�~?;�I?v�?���>�H���wؾ�-0>�D��˱=Y�-Mq�=�����?0'?F��>�쾶�D�)W׾�i�I�>*(�@~G�go��Zl-�-��<�涾�1�>�Hs��ޕ9�8Q��n3��n>�Œ^����>�FB?���?�	J�X���vQ�$������*
?�)_?Wp�>CG�>�G�>4<��%���h��	>ώm?���?�s�?8y$>%��=9��9�>�'	?���?w��?,�s?^�?�1s�>�i�;�� >ؘ��F�=$�>%��=�=�o?��
?%�
?�m��8�	��������^���<��=���>p�>��r>��=R�g=v�=�*\>؞>��>1�d>-�>�L�>������I*?��<`�{>l)?��K>��¼y�����<��ڽxh�x�������f�����ؽz�n=X=�Q�>�ɿ�n�?&��>#R5��x?���b���`�>q��>�x>/�?���>�cw>nH�>Y��>[�">�+�>a�F=�@Ӿ�n>���[!�"0C�ĂR���Ѿ�oz>Ȝ��!&�E��	B���"I��f���e�-j�c-���2=�S��<�F�?���w�k���)�J���H�?�i�>�6?�Ԍ�s]��t�>���>��>{A������}Ǎ�\cᾒ�?I��?�|c>��>�ZV?h-?�*���;���Z�]Su��,C��Be�f_��`�����������@`?�x?�X??`(�<E�v>p��?��%�b]��Ĩ�>X/�p�;�BQE=�{�>?豾�Y�N�ԾRľ?*���F>�Sp?3�?;�?��\��m�u'>��:?��1?�Ot?��1?i�;?�����$?co3>F?�q?0N5?��.?"�
?=2>�	�=�����'=�6���7�ѽo~ʽ��C�3=p^{=�͸�<��=T��<ʙ�£ټ��;I%��F%�<!:=z�=��=�*�>�a?��>�->C_>?�K=�5C�0�˾E�C?�	�=҂��V����ƾ�1�61<L{n?�S�?�:h?>�r=SE�n��q>I�`>H>Eg:>�E�>�  ��,c��=j�=7Dc>�R�=��Խ1о
Q#�w)����=�KB>a&�>Qz>�x��=��=��n�/��y��>��������]��ԢX�"� ���9��\�>dEA?8�?�jG<-ξ�J=�Kg��$A?>7?�4?��?�z=�/ܾ�A"�E�;���+���>q�ؽ���w%���ѝ��(�Nm����O>��Ҿ�렾
Zb>���"a޾F�n�J�K�羋NM=�}���U=����վJ@�h�=0
>/����� �A���Ϫ��2J?�}j=uj���MU��q���>���>��>�k:�2w���@�������=���>Q�:>	������+zG��1����>SQE?�i_?�c�?�$����r���B�.����⡾'f����?�Ϋ>�(?�fA>�G�=Ẕ�f �Ne��G�f��>X]�>;��*�G�xמ�JB���$�Qh�>�'?w� >�?�}R?X�
?B�`?t*?:C?�C�>[F��B���1&?�S�?�F�=f�ѽ~�R���8���E��R�>��(?�C��k�>��?db?]�&?#�Q?�?Gj>���:@�ڸ�>�)�>�OX�3���Wj^> �J?�&�>_�Y?�#�?R?> �5�⢾%᪽�a�=�s >ߟ2?��"?w?t[�>&��>����g�=���>O�a?wʂ?�"p? ��=�?��3>;O�>]��=*�>b��>��?;O?��r?\=K?���>v�<����:e��.�j��a����;WVi<���=�'�����~�qm�<���:�ޭ�R9b��D�<�����u�.<���>�>�J\�UX�>W4��;�����>hS���'�T���:��ɪ2=�$�>n�?��>��)�p�;>Gu�>���>��E��<?���>�|?ݖQ>4XK���X�1�3�->�?�����p��J����f���d= H? DU?�M���L �O�b?��]?@h��=��þz�b����g�O?=�
?3�G���>��~?f�q?U��>�e�+:n�*��Db���j�&Ѷ=\r�>LX�S�d��?�>o�7?�N�>/�b>'%�=iu۾�w��q��h?��?�?���?+*>��n�Z4�a����ۑ��]?>��>����V�!?����>Ͼ��������Kt� ����j���,���禾u�&�媄���ս)�=(�?;s?�q?�`?�,� �c��H^��~��U��������JE��"E���C���n�$��=���I}����N=��:Ch����?m�?Z���v2�>�ö�^�������>"2�������>�7=���=lݽ=s0������f����*?9K�=i�h>�LB?��y��F��?
��H2������N>Sg�>���>��#?�=��g���N�UԽ�"�J��C�\Hu>�}c? �K?Q�n?_��h�0�����]�!��v,������<C>��>4A�>�kX����YJ&��c>��r���������	���~=!�2?��>�u�>"�?��?�P	�fR����w�AX1��˄<#�>�h?Q;�>���>��ϽU� ��>�Tl?>��>zw>����Q�`wg���G���>�~�>u5?ʈ�>ϝ@�/�`�0I��膑���+��x�=�Pj?^ɩ�ٸV����>�FV?�g�%�
���{>)J&��p�L�پ��X���=�0�>���=��>{qľ���yO��b)2��)?b?%���ܡ)�80{>:�!?f`�>Zȣ>��?���>+������;?�^?Q�I?$GA?6I�>��)=O$���Pɽe$�B�$=4�>��]>��r=͹�=��AX\��c!��HC=��=Wg�l�����$<�Ų�.c<L|�<�7>�)��9����=����Ӿ]O(�|u�-�,�=m����Y��䄾�Ą��s��=h�hҽ��}��3����}������?(t�?�)�E�9�"����7��$�ߗ>�<���W���Ҿ{����1оU-�n�Ծ��<�#9M���&��'/�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >kC�<�,����뾭����ο@�����^?���>��/��p��>ݥ�>�X>�Hq>����螾a1�<��?7�-?��>Îr�1�ɿc���l¤<���?0�@k�G?�E�@X̾��=`Ô>"b�>��(>aʉ�]6�=��e��>�ה?�ژ?>��==�F���=��E?�e�=�*�||=c�> R����=}����^>W��>��T��ʖ�jK��i>&�>��_�!���2v��/!=�Y>�Ti�L�<=8Մ?8{\�Gf��/��T���U>��T?L+�>�;�=p�,?�6H�)}ϿS�\��*a?�0�?Ȧ�?��(?�ڿ�jښ>��ܾi�M?�C6?��>�c&�R�t�Q��=:�����T�㾒&V����=���>?�>΁,�a��;�O��T����=����ſ��*�$��tm`=�[ļY���ͽ� ��Gw�����T�c��һ�RO=���=(GM>b�{>_�5>\�_>��b?�cr? ��>��">�_�?����˾NTK��犾f�E��ˤ�ĥ'�c�����������bP��|��U¾8!=���=/7R������ �"�b�\�F���.?Zu$>g�ʾz�M��|-<�qʾu���uބ�~好�-̾9�1��n��͟?��A?=�����V� �9M�F�����W?�F�}���ꬾ��=�ϱ��=S#�>���=}��d3�|S�%�.?��$?�hľ������>�θ��.=#�0?�}?��=?h�>��'?�0��jD�ߖ�=Ay�=�@�>�4�>��>�D�����/)&?h W?|�D���ѾwHo>�l��"�o��A>O�>��L�-ϼ��>N�7�~��d���_�C;>B-W?�p�>^�)�Q���O�� _�A}@=�ox?��?*��>�pk?9�B?,j�<������S�G�
�,Ny=0�W?Ji?�>81��B�Ͼ���]5?��d?M�N>sgf�͘��l.������?@@n?\H?���s�}�X���:���6?��v?��]��V��@��eT���>:;�>��>j$9��o�>xk>?�"�v1��)����x4��?0�@a��?a<�"���=1?��>?P�2�ƾ�)�������l=rT�>]%��Ju�v��{-�\�7?@�?�l�>���������=�ٕ��Z�?��?z���cDg<R���l��n��S�<�Ϋ=���E"������7���ƾ��
�����࿼ʥ�>DZ@�U�u*�>�C8�\6�TϿ(���[оSq���?J��>Z�Ƚ����?�j��Pu�_�G�3�H�ɥ���z�>��>a㏾��v�<�F�DbB�G�H=y�"?�=�/�=2�����"�X5�`�X=(��>M?*?^�����V��?�'���߿���������G�?v�?K��?zYA?��>	�ݾZ��N��<��7?<G�?#m?|���c����H<һj?FJ���P`�i�4��DE�KU>m3?�L�>��-�tQ}= 9>{��>mY>r'/���Ŀٶ��������?L��?Ev꾊��>���?=w+??l�;8��O\��n�*��.��<A? 2>����9�!�E$=��Ԓ�ΰ
?�o0?�����[?�*V�e[���?���>����>�m�<������� k�)x��}��{k��%�?r��?Hr�?�~H�	���1?{��>j��9Ӿ�m��f3t>h�>jd�>��=�\�=X9,�"[��kj>��?C�?�'?-����x{>��?/7�>��?W�>>�&�>��<S
����W��w=d0>g'�=\R?��:?�ۭ>�����֫��4@�*�;���V�o����P�.�>�u?I?o,=>�n���򽽧)?����4Ώ�T���qZ�D�� ���z>j�A>݊�=�Mj��Vվ��?Mp�9�ؿ j��"p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?[��D��u�o�y�>���?
�@�ծ?ji�)J?ڄ����s
}������<����==�7?9ﾙ�w>��>�O�=��v��i��96s�u7�>NQ�?�
�?�m�>�'m?tn���C��=Y�>J�k?`[?+�B��D�aE>.?���O����� �	Ag?�@�v@�Y^?�͢��hֿ����_N��P�����=���=Ն2>�ٽ*_�=��7=��8�B=�����=t�>��d>"q><(O>a;>��)>���Q�!�r��\���S�C�������Z�C��Xv�Xz��3�������?���3ýy���Q�2&�(?`�R�=9.Y?��S?�Om?���>�މ�SP >�J�{�G=��)I�=Jw�>
/?�G?2D'?�k�=�J��}gg�����dP��~=���j�>�M3>b�>���>�8�>�;��9>�z@>���>���=��Q=�Ȓ<��A=fMM>lj�>^��>���>��=>��>xʹ�JJ��l�g���s���ǽ@^�?�0���7J�l��8���Aҷ���=+6/?xz>����Eп����F�G?:��HY��(0�jr>��1?#�V?iB>�9���=M��$>���OCl�-�=�#��μj��\)���Q>�?�f>�u>��3��e8�Q�P��{���j|>46?�趾E9���u�ŲH�Ucݾ�GM>_ž>.�C��k�8������vi�1�{=x:?c�?�7��D᰾Q�u��C���RR>=\>b=�f�=gVM>�lc�R�ƽ:H�mg.=|��=+�^>��?|��=�l�=Ҷ>�H��8M�<{�>X�5>�9">Ě>?�Q&?���@��:��R�����L�>��>3�>Q�l>�\��f�=L��>�f>�^'=f� �0ν���1>�n��V:a�Cߥ��h��(�M��>�c�=����)_���=l�~?tg��G��j��G����,?�Vq?L��>ګ�zWW����Y�t����?9
@�+�?�o��;�:�1?��?+V������?@D�>;Ye� �����>�r��)"ʾc��[:<�d�?��?�=��� �{�l�=H�$?�y#�Lh�>{x��Z�������u�J�#=N��>�8H?�V����O�c>��v
?�?�^�੤���ȿ5|v����>W�?���?g�m��A���@����>:��?�gY?voi>�g۾>`Z����>л@?�R?�>�9�~�'���?�޶?֯�?�ȃ=Ϭ�?3��?���>�I����b�������-1>���=O�> ��>+r�B�I��吿� ��x1z�9� ��q>�, =㏁>��a��ݠ��>�`�Do�<�Y�2�>��>�h�>�ڇ>6v?A�>�~�>���=tr�<�K��2+����K?���?B��3n�P�<顜=в^��&?�I4?�h[�u�Ͼ[ը>��\?U?�[?^d�>,��U>��8迿~��e��<�K>�3�>�H�>%#��%FK>�Ծ04D�zp�>*З>�����?ھD-���\��_B�>�e!?ד�>�Ѯ=ۙ ?��#?j�j>�(�>:aE��9��O�E�ɲ�>ޢ�>�H?�~?��?�Թ��Z3�����桿��[��;N>��x?V?jʕ>X���惝�SnE��CI�V���\��?�tg?�R�0?42�?�??_�A?b)f>��Bؾ����> �"?V'�gAC��5*�Ь
��V?�c?���>�//���ʽK�������.�?��_?�/)?���Uc��`þk��<���f,�ޓ�:����/>Ӹ>qi��M��=��>H��=�n� }A����O2�=�"�>̓�=W&��Н�Y?,?�D�t��=��r��?D�G�>�+L>����ۢ^??9=���{�
��z��,KU���?���?�r�?˯���h��#=?��?��?q��>�q��g޾�t�~bw��wx�h��<>m��>�qo��'�㘤�[����:���bŽ��.�F�?���>���>��?*~!>�m�>6r��+J2�Ϟ�����tVY�j�A` ���)��<�����M���a�W'ؾyYm�>�-@��>҄?�pP=_�D>P�>2u>��>Tq>� >2H>^�[>/�(>�K=Dz<����Uc?���Z&��ߩ�G���_�?,7s?K��>��d���m�|���$~*?�+�?Zh�?�>�1-�"���#?��>R���1?�I>��=J�>�����U���3���=�N��E:�AT[�V����_�>Y?=��=v�ž�v�<S���=Aw?��+?��0��]�U�n�kM��M��鰽�@X�p���U`%���r�?돿�W������n ��S�=�0?ł?:�辿Aо�T��	�d���>���i>�+�>p�s>*U�>�B>�
�d�(���\�oJ(�־}��0�>d�w?���>t�I?�;?�wP?�tL?���>�c�>�0��7E�>r|�;C�>s��>S�9?��-?�30?9w?Iu+?t9c>�m�����yؾ�?U�?F?�?�?�ׅ��Wý-����d�>�y�����с=�b�<�׽�)u��oT=��S>�x?"{�Ռ8�iD���-j>�Y7?E��>��>y쏾�̀�`m�<���>@�
?(l�>`����4r�EZ���>췂?�����=T-)>���=��z��꡺�~�=�׻��c�=h݇���;���<%�=�W�=��V�x2��;^�p;�J�<�{?��&?�w�=�W�<j�彴�(�n�׾���=�֙>8�r>��[>�Ht�G�|�}����Ap�7�y>��?��?�A��|`�<��0>Rxi�����������1;��?�Y�>s�B?�	�?��<?�-$?���=���'���}���I!̾�3?A!,?>'����ʾq�Y�3�L�?�[?[;a�]��j:)�t�¾>�Խ"�>i\/��/~�B���D�y��#�����A��?׿�?�A�3�6��x�忘�v[���C?, �>�W�>L�>w�)��g�:%��.;>��>kR?�
�>�I?��y?H#[?�C>)9�%���/���s����'>\�??�	�?���?�x?��>4N>�^.�p�پ~���lS�뽿چ���h=�T>�,�>��>\�>̴�=!Eν�蜽�F���=��^>�%�>�ץ>��>?�y>�l=��Q?
�>�3���Y������>�9�<�|x?���?ø?efY=[�+�]����?X��?a��?i��><pؾ�{Z=*�=�g���;�.ɣ>�v ?Y>s��
[�;�	)>���>^#�>�.)�MN<�����Zf���r4?�؎?n���7Ŀ,`��+��d�_�Ҁ�Ɛ������3d��_Z�U��W������+o��ˆ�>�������C�о�9��>z3�7u?7�=�$>ӏ>��2;����vI�Ԙ=1�=߷��4*��	`�����b|�<���B�׻��R=��2=T��<���?qB�?]5?�T�>��Z>츺��+۾��>L��>��D?J��>�;㽆	Ⱦzޏ�A�۾F���-0��|�
���ʭz���=�����t\>���=���=�" >;^��7\�G|�=��=���='�
>hAf>��>i3=�6>��uw?�y��㹝��/Q�>��#b:?�V�>��=�Eƾ��??��=>Y��ѓ���:��0?���?`�?�?�ai��Ԡ> [���S��,x�=�Ɯ�	�3>!X�=�2�%'�>�QJ>~��[@��/S���T�?E�@Ǫ??lߋ���Ͽt0>Z�7>('>��R�Y�1�^�\�m�b�ivZ���!?�J;�mM̾n.�>�=�)߾�ƾ�w.=q�6>�tb=�[�T\��י=��z���;=�k=,҉>��C>�Y�=52�����=L�I=���=R�O>[�����7�,,�޵3=\��=�b>�&>��>���>��?�S|?���>���2������5ή=�Q�<���>�$��>��>|�B?7�S?�_?�Y>����?�>!�>��D����klھ�^���=���?�%�?��>gʽ�Hf����5�a �<�
?P�?(�>�+>�U����:Y&���.����о4��+=�mr��QU�a���Cm�/�㽶�=�p�>���>��>6Ty>�9>��N>��>��>�6�<�p�=⌻���<� �����=K���U�<wż]���w&�Y�+�S���B�;#��;��]<Z��;:�=6J�>�{>}s�>zޔ=o���.>�i��@RL�8�=J���>�A���c�43~��P/���7���A>nV>]��]4��H�?F�[>rH@>�:�?�0u?de>����վM��aUf�2�S�a��=��>�<��
;��`��M���ҾK�>�6�>�ç>��g>I,�=6:���X={���.�1;�>�煾�������q�*륿����Ff����lF?ɩ��MR�=XÀ?�/I?1�?H?�>Q���]��ʎ'>�����5<F��
t��I���O?0�$?��>�Z�C����V���=�>B���Z�
g��7�=�o�=����>Ѡ���Ǿ�yA�}E��,����M��hi�R�>S?�?�?�[�:�h�]�F������N��<�>4v\?Q�>:R?]*�>z�u��g��;���e>o��? t�?�|�?��0=�q�=/���("�>	?Ɩ?l��?�ds?�^?�'��>Թ|;Z�>���]z�=a�>�K�=���=�b?�
?��
?
�����	�-�����Z^���<#$�=�[�>O��>`�s>�{�=)Mg=J��=Ȯ[>|�>�ۏ>Qzd>Yѣ>�B�>D���w���#?r.=�x�>h�?\:
>����
)l��<���>6_�C��Gh|��'���;��2��#>��� ?��ҿ~��?�;I>q6���?AY
�?D�c�i>o_�>�>"V?�>��>���>���>��F=��v>AI>ԍ޾Zs>r�	��j"D��aW���Ӿ0�v>(����/5�Z� ����R�_G���
��k��[��ej8�K�=&��?#��c��] �ʷ�n�?&p�>��2?9,�����&�	>G�>�B�>�_��<��Bh���c㾃��?�$�?�Wc>0��>u�W?M
?,�/�83�uLZ��u��iA�Ie��e`��ɍ�%w���/
������_?(y?t A?d��<�=y>+��?��%�ُ��e�>\&/�* ;��>=ݦ>�����a��Ӿ�ľ�r���F>�yo?��?��?�X�H�o�S|'>��:?,t1?mat?��1?�s;?V����$?�3>�`?&�?�G5?��.?T�
?F�1>��=����'�$=�ޑ�����fѽ�3˽�[���4=��|=W�9c<r�=7��<���#4ټ�3;�������<�@:=`ޢ=N��=T��>��\?��>y|>��8?z(��_5��d��8�/?�FH=l�}�y���Q����7���d�=�k?���?��]?��R>�&F��+8��3>�ڈ>�v>6M>�հ>;@�}�I���{=T/>�&'>���=GAp��_���+��J����=�X%>{ ?ߡ5>��{�pWp>�c�,r����>�]L�	�ݾ������>��
+��1,���>1D?�t?{��=��ž$7/=�Gr���.?�<1?=N?��?b>=�_����3�bR�Sz�Lu>�\��i���7�������%�l��=��>p���ޠ��Zb>޼��q޾j�n��J����ABM=��(bV=e���վ�4����=� 
>����	� �G���֪��0J?-�j=~x���dU�Ko����>���> ߮>��:���v���@�%���c7�=ض�>T;>l[����[~G��8��\t>=SM?��c?5�?���U�p�(�=��W��檛���j;�7?���>a�?`2>Qo=�z����sm���P�[��>��>%X�1sK��@��:Y�U���Et>=k?9��=��?4`S?�	?�`?��0?f�?��>�:��/�Ծ�@&?��?���=_kԽ�T��9��(F�p��>�g)?j�B����>�?d�?�&?N�Q?��?�>ͯ �N,@����>VX�>��W��i����_>̩J?�>�OY?�׃?��=>َ5��Ң� Ω��:�=>�2?�!#?߮?�˸>B�>�����=�=�>Ͳe?�ق?�m?��>�?	�<>�{�>���=���>rE�>}�?/cJ?Rs?1xL?���>���<>f����ɽ�iY���:�&%<]Hj;�C=�o２Ev�R3�K�<V<x�����!О��q �����q�<�(�>���=�s���$�>���k;qY<�/\�^���Ѿm���O�<�?�>�S)?h�>L��3#<>�8�>j ?�Q!��� ?���>v?~"�>�g��b��;ٽ$� >:�1?%�e>ե�� ��0Z���=�t?t�o?�$ľ�l�W�b?��]?�h��=��þi�b�C����O?=�
?��G��>j�~?V�q?���>��e��9n����Cb���j�&Ѷ=�q�>XX�|�d�?�>ݜ7?8P�>��b>�*�=�t۾�w�>r��D?V�?�?���?K**>*�n�K4�=��������]?+��>gj��}�"?u����ξ����`��ӧ�����ά�Z���u<���&�m����/׽Q��=,�?B�r?ftq?�&`?�� ��d��h^�u��&U�f�!�dkE��D���C��n�������9���S=��ʃb��ۭ?��?/Ǥ��v�>����T����KN�>����~�齍��>D�=|>[��=e���u˔���F�b
0?%�;#s�=I�l?C�P�3<����O`�}G��\�=;�>.l�>�pJ?��>�K�o@
��ʾɏ�Fn��g>�Qg?��N?��o? �	A1��m�����w�*������:\>��$>���>��X��6�|�(�,7?�GKw��s�ߔ�8��I?=b (?� �>�s�>~A�?���>m-��߲���q���(��b�<��>$�j?�2�>�O�>7Ž��'�#��>�G�?�C#?m9�>�o��;Jܾ�RW��<:�>��>~��>b�6>)��Sd���G���*�����UhԾK�t?��Ǿ7�M����>~;?����ؽ2Q�>h���^M����>U>�ڱ>Qw�>�+�=�W��%��a4�M�W�P�r�)?��?�����+�z�|>�E#?&�>��>���?B_�>W[¾_R�V?Z�^?JK?�,B?w*�>�G!=�����*Ƚ+<#�KT1=�ć>A�[>��b=���=8~�`s^��!��fV=�W�=�r���CĽ�U<�l��#��<���<A/>��ܿ_�I�F��)��s	��bU���|n�R$�WI@�����
ľ�7������Q+�i������c�=n�ۀW���?Zn�?YcD����*ڛ�H��qN�D�?�|ɾ�Ͻ�i��l@��I�����|�����<��I�aBR�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >_C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾s1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@�B?�/4����v�=���>�!�>���=��~����-�����>.�?��?*�=w4O�bž�_gQ?��o=x*9�]U��_>���;hkV=ͧ���L>{u�>����F�UgU���>�Q�>��Z�Nw��sT�����;�q>>��JKG��օ?�.U�s�n���O�U2��{K>�P?��>_>�G?�fV�I�ӿY^���X?���?��?&�#?�����k>r=ؾs"8?Ae0?�>M4� ���(���Hl�݁վ	nU���.>��>��>���� �\���Z4Y���=ym�9ǿ  .��r���=Q:Y=Fb��H�?�.Z���<:���]���潟��=�N	>�T>��Y>���>f�R>^�^?�v?d+�>�}>� �p���`�վ�<�,{�c����֑&�ɼ���V�
e��	��=��-��2��y=��ҍ=�6R�ꇐ�v� �(�b��yF���.?�#>�rʾ��M��C*<ȤʾHת��n��F5���˾�B1�q�m���?��A?�煿�V�S$�*�
�$���t�W?�����嬾j��=�����=�G�>J��=�����2�kS���0?�?a.��A����*>L���7g=mm+?[� ?��A<|X�>o�#?��.����o�W>t�1>��>ڤ�>��	>.���@ս�,?��T?Dy�@Н�鱎>���-�w�Y_=s>��3��Ѽ��U>�W<7菾r����W��F�< (W?v��>h�)����`�����wZ==��x?ђ?.�>|{k?��B?`�<�g��[�S����dw=�W?�)i?��>򄁽�	о����4�5?��e?��N>ch���� �.�1U�f$?��n?�^?+����v}�<��2���n6?��u?R�\�
��E;��a�Tˠ>c��>X��>Ŵ=���>��4? �;�ߕ�!l��c�7�~�?�U@���?��������<��>��>^c�*j���^����̾�.�=�T�>(���d����B���F?�c�?� ?_���?6����={ٕ��Z�?c�?����<g<����l�~n���z�<�̫=�lA"������7���ƾ{�
�����yٿ�7��>Z@V� +�>�D8�6��SϿ��4[о=Uq�7�?v��>ǞȽ����+�j��Pu�g�G�V�H�礌���>�f.=��z�<�����O���Q��`��b?}��HR/�)��� ٓ�H?���g>���>���>"@^>xp��D�<�p�?�M����˿���L,�Ɂ}?$˷?��?&9u?<q&����aZ� U=��!?�h?aC?ik��]<���=�j?_��.U`�ώ4�CHE��U>�"3?�B�>6�-���|=�>��>Sf>�#/�i�Ŀ�ٶ�����5��?ǉ�?�o���>n��?�s+?�i�
8���[����*�m+��<A?R2>�����!�`0=��Ғ�X�
?�}0?�|�.�� `?�b��'r�v�/�^����>��%�*#[��>�\i#���g���������ج?8��?�c�?H����ع#?-��>�E���h¾�A�<4��>z�>�JP>�I�F@u>�t��@�x�>�;�?���?��?���0����V�=�}?vp�>C~�?�$R>�z?�d[=}3���!�:��=<�=;�f< ,?o�Y?���>�J�=�sr���4��.I�\�`�(�(���@�`~~>�	D?�M&?�}�>}��/;��������_2�h\Ѽ�0��!*<;&�P��x�>��Z>7�>�I#������?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji�|W	?������XUz��h�3H��+>��6?�q��P�>J��>���<��z��k��/j}�X�>?��?:�?w�>��?�5s��G��|(�o�_>�ہ?��?Ž��m�=�G?�{&�Fӆ�)H����Y?R�@L@��Z?䷘��hֿ����NN��R���t��=��=�2>��ٽO_�=-�7=/�8��<�����=g�>��d>q>M(O>�a;>Փ)>���K�!�r��`���W�C�������Z�?���Wv�Iz��3������q?���3ýy���Q�2&��>`��#�=��_?�V?22h?��?h;��>�� ��uF=����B�=��>000?��@?I?(0=߽���kl������ʭ��Ꮎ���>5>>�>>�>җ�>��̺�XF>��#>7_>;�=��"=���V=:[>ú�>�,�>��>�C<>��>Fϴ��1��j�h��
w�e̽2�?|���V�J��1���9��Ѧ���h�=Ib.?|>���?пd����2H?'���z)���+���>��0?�cW?!�>��U�T�1:>B����j�2`>�+ �|l���)��%Q>tl?�j]>s~>�0�m6�}?N��A��"S~>�'0?����&2K��	z���I��I߾�J>��>�=��e0�����*z�~s��t]=�U;?��>��۽����߸��P���#_>��_>B��=���=+TE>kvu�����1uH��8�<���=�|]>�$?�*>���=U�>L���t�T��¥>�J>>\A$>'/>?3�$?%T��M��bT����,��3x>_��>�>3�>��K���==��>��a>�u���u��u��Tg=�m3V>QZ��v7]���q���t=/���+��=��=M6�i�B��u+=ug}?C�������A�ξ��	�t�4?���>��l;�㌼��h*��+���p��?��@��?� �RR[��!?�P�?�q{�d��=�>��>��Ҿ7_H�.	?�I��w��x���o�g�?E�?����:7��l�i�t�>z�)?�ɾTh�>�x��Z�������u�U�#=M��>�8H?�V��)�O�r>��v
?�?�^�ݩ����ȿ3|v����>Y�?���?h�m��A���@����><��?�gY?�oi>�g۾?`Z����>λ@?�R?�>�9���'���?�޶?ԯ�?�=Ed�?xs�?�z?�t����)�ڵ���T�P=�[�>�W�>�Ԭ>�*����U��ͥ�p���og�`�M���>`�����>$��Uyu�p��=e���:��C}��Ђ>��>>wnR>�u�>**�>G?�>�#>�p=�-��7�0���K?���?.���2n��N�<z��=!�^��&?�I4?3k[�z�Ͼ�ը>�\?j?�[?d�>;��N>��F迿6~��y��<��K>*4�>�H�>�$���FK>��Ծ�4D�ap�>�ϗ>�����?ھ�,��<S��JB�>�e!?���>�Ү=�� ?��#?��j>-+�>bE��8���E�o��>���>DI?i�~?�?�Թ�c\3��	���硿��[�.N>N�x?CS?�ƕ>���e���5�E�%SI��������?�qg?�M�s?2�?��??��A?-&f>����	ؾ������>o31?$�1�>�I���C��B�\�0?m?�q
?�">y�����L�֭?�_��Ӓ?�r?>?�쾣�<��x��2��<)��=���=�-�<<%r�=@��Q��l�,=P�o>qhn>*o��S����潄��=ʛ�>vO>ұ{�y�k�:?˥�=N�n������2�2��7Q>�Of>v��ZP7?`�5�%f��]�����-h��0~?A=�?�<�?�����f��K?��?q�+?���><ʹ��\ھc�̾5�~��V�$y.��$>���>�,�*�#�i��rУ�s�i���==	�׵�>Uw�>� ?�V�>Q%>�Ӳ>�����i)����9�W`�ߣ��W.�,�$�xj��ᦾ�C��u	��(о�i����>VF��楎>�?MW#>ϖ�>>\�>H��;Ҷ>~f>�8_>|�>�cC>��>���=�+��N��!�`?�	�{+I�s��x����e*?�V?*�?�V�=����#�2a�>���?�M�?0��>���2E$�;?��-?�<j�o��>w��H��u�=Y�=.6>"{���	K>�#?UTB�r~}�6�u��y���?~�?D4>S��a���5����Oo=�N�?��(?��)��Q�6�o�3�W��S�}g�Q)h��c��A�$��p�C�`���$���(�?�*=��*?��?����)���$k�0?��^f>��>�"�>��>\�I>��	�\�1�� ^��K'��Ã��Q�>]V{?"��>��I?�;?=yP?vmL??��>*X�>J5���]�>��;��>
�>��9?^�-?50?Hz?�u+?�0c>Hp����ؾ<?��?�K?$?�?vم��uý���u�f�y�y�v���/�=�!�<Ь׽�1u�7�T=T>�M?��T�8������&k>��7?���>���>=�����ˬ�<V�>�
?�@�> ��xr�]X�ec�>��?���4=ܮ)>��=q�����ͺ�4�=z¼���=�\���W;�� <��=n��=.Xu��$;���:��;tX�<A ?��?���>�,�>����3y������r�=TW>�ON>�>�fھD���s���g�7�q>�?\�?զr="a�=LV�=ҟ����]P�Aÿ��]�<v]?��#?-lR?4=�?&L<?��#?<��=�������΅�Lꪾ!�?q!,?ۊ�> ����ʾ�񨿌�3�o�?�Z?<a����d<)���¾��Խ�>.[/��.~����D�u���-���y����?տ�?&A�i�6�Ky辉����[����C?!�>gY�>��>7�)���g�$&��,;>��>�R?��>��?لX?��u?��F>�U��i��p뜿�]b�|�-<+6?�c?�M�?M��?���>u(m>�3���󾾅]���7�!~��:��#a<��D>3�h>�F�>hN�>���=̄��f̽�׮��5=1�X>�y�>֒>��>UO'>�p�=�W?�r�>�o�?h+���i��av����O�n?���? �>=��=Q:�0w������	?/r�?���?���>�5����k=�c=B����f��Wk�>h�@>�A>���L8��>>��>G�?��/�A J�u�Z����c$?��1?�f�=,ƿ�{q��tr�~����<�ߏ�>�_��\��,V����=T���?�����Z�8w��QO��촾���m	|����>je�=��=]S�=<�<��ۼܩ<��M=�ԍ<r-=jm��w<C�9����@6��
���'�f<ױO=�.��ve��un?�HO?��?��x?A?��>EP�8�>��3>3a2?3�?]U�=�ӏ���j�����}��A�����3�߁��D�Ծ�k��m�����N>h�Z>$t>�{�=�2>,7�<�b���I�� r�<���=��=O9>n��>�#�>��w?�{~�2����\��[��#4?���>���<�8׾3*%?���=�p��gط���� �p?�>�?��?<�"?=dz�.v�>J�������6�;&;|�/y)>a
�=�+a�Y��>Q�=A:������-���?��@??����*$տ�h>Xu7>y,>��R���1�^E\��b� EZ���!?W1;��1̾J�>,E�=�߾|ƾ�.=5p6>�	c=�-�]C\����=	:z���;=�l=�҉>��C>9�=�
��7�=�zI="3�=��O>�M����7��v,���3=h��=�b>�7&>a��>��>DY?�6q?��>�w��|��ZZ;�u�=���Y�>��!=\�L>N�>&Y6?��O?S�P?m˅>v>�Ͽ>BƤ>��2�ڃ�l���:���<G;�Y�?��?�ve>�b���ܽ<���2�J|���?ם?��>?�>`G���߿��@���$�}��=¯�=2��=*���>��;>*�=���!2��!�=�Ƀ>p>�>��K>f.>Œ>zd=�M�>�߭=�����>zo�=�>��m=1?���G�=x'>��f����<���iϯ=x>���6+�*
>gh>R6�=��>jv>�/�>���=G��>�4>�:����M����=⸾��C�=c���y��a+��C6�Ņ9>;�H>Y^��������?n�d>��A>)��?�_r?�>����ɾ���tJ��G�H��=d��=��F�)P;�_��	O�^5ξ>��>���>�)�>��l>E,��?��_w=��� U5�C�>�]�����;��Bq�hC�������i��*��B�D?�B����=�~?
�I?�ӏ?\k�>�L��o�ؾ�.0>�2���|=���q��0����?�'?�r�>M쾓�D�J0˾���5@�>�3f�]�B�g����� �$�e=�.ȾE*�>^Ǿɘʾ��9�0���^(����D��k���>-m:?$��?�8���x�۸N��]��v ���?,@q?���=�y�>f�>�y�y���L�������Aqw?yL�?�X�?�e�=�c=����6�>���>��?�w�?�Dr?�A��>�>(T�<��J>ޑ3��n�=���=*b=o��=,?U�	?�P ?��d��g��P�5q�lr����<�js=8 �>��>�x>b,>b��=���=jXc>玏>%��>V�h>Gj�>��>����	��v&?�J<���=��?䧮=�([<��#�vи��ɩ����E�L�O�uK�:&�/&�����;���:�	�>m�׿왤?�fK>�h�b�?�27�\t���">��>6!> �>�F�>jş>���>]a�>�c�=�>�wH>rFӾ�>����d!��,C�W�R���Ѿ�|z>����
&�	���x���BI�n��<g�Bj�9.��@<=�dн<H�?�����k�4�)�����]�?�Z�>�6?�ٌ�E
��I�>���>�Ǎ>zJ��+���2ȍ�hᾐ�?	��?pec>ﯞ>��W?0�?��0��i4�6�Z��u��rA�&e��x`��Ս��y���1
��澽P�_? y?HA?+�<��y>Ջ�?@�%��я��I�>�/��5;�k�==��>_O����`�uqӾ��þ���2F>Y�o?��?2?V�OK���t^>4�)?#c�>ʃ?)9?;Q?�\�=��8?:1�>zr%?y�#?͸"?��>>��> 2�:�<E>}"[>sl��{8���=�f�B��5@�j!�;f	�<��8�� �=*pA=�=���=�%�<d̥=u<f����|=w�=��>c�4>���>�d\?F��>��>��7?m� �9��믾��,?�?+=�}�������ס�G.ﾹ[>~k?��?�|Y?P{e>��B�f�A�e>���>��'>�5Y>�7�>�g뽴�E�IL�=:�>��>���=hN������	�����#�<�;>�<�>�>����<iG���fϾΒ>p��� ��<��o���F�G�+ub����>ӴE?z�?���<3��������[?3M]?U?RŌ?�	�;_F޾</��G>�Z�c���>$K�=b���\������6�I���̽X��<	R���ޠ�Xb>���Et޾#�n��J�S��sJM=���YV=����վ6����=�$
>s����� ����֪�_1J?�j=x���bU�q����>���>
�>��:�G�v��@�V���&6�=���>� ;>_����~G�/8��L�>�BE?P_?Lq�?v͂�ns�*�B�a�������X˼?�?4�>�R?��B>+,�=�]������e���F�_�>��>7����G�i��}��̻$�uΊ>�>?��>��?h�R?9�
?߁`?E+*?�L?��>t���%��yI&?�s?���<{�7<&50<��$���%�n?��>ea��ސ>��>��?�m7?y�\?�?D�|>��/��'�|�>��{>}�O������=j|g?H�>c�[?���?�xA>�K��U|��S���=��>i9%?i�>3B?��>b��>L���m�=���>�c?�0�?�o?�=;�?�:2>O��>H��=���>O��>�?OXO?;�s?��J?��>���<v7���8��Ds�i�O��ǂ;xuH<�y=��3t��J����<��;/h��#J��a��G�D�
���Q��;'/�>�Pg>i����g>�~�����>�û�=�v
���ܾn;�:�>��%?j�L>�6��ͷ=Z�>b?c�(��-=?)G?r�?��O>�	��:侒�(QL>(|?��`=}����g���\��ɩ�L��?��r?	$羂��O�b?��]?@h��=��þy�b����g�O?=�
?5�G���>��~?f�q?U��>�e�*:n�*��Db���j�$Ѷ=[r�>LX�S�d��?�>o�7?�N�>0�b>.%�=iu۾�w��q��g?��?�?���?+*>��n�Y4�>�������D??��>�����?�vB���̾�ˁ�+��Z2ؾX䟾$����sT���7��Ӆ���̽õ�=�{)?�À?^	i?;*m?����|�o�h�#�|���L�D�߾64��S�hQ?�xJ�>�r��*�-S���ģ����=}�	��D�2�?V�?�[�����>&���	��,�@+�>|�V�	"�=�PI>��=X��=B���و��a�i�y�$??N
=H�>�`?�nI��>��U*�4�B����Q+�>)?v?�M=?�l+>��f�V���3��Ғ+��|ɾ�<v>7�c?h�K?,�n?�� ��1�j����!���.������B>��
>II�>��X�����n&�f.>�Ls����󁐾��	�kπ=ƥ2?��>Ed�>�?�?��?(�	�?뮾F�x�J_1��n�<)�>w�h?��>py�>�ѽ� �f�>���?�t?eM�>`�;����������
)�#N�>Uf�>^�?�8>eui�@z��K��������ci.�F#??�ĝ��9&��0�>�W?D�=�a��+">����n��&���'��(Q=���>|r�=_�>4�򾾣��|����u�U)?Z#?H~����*�E�|>�E"?�?�>�y�>�f�?
Z�>2�þ��⺀[?�^?��J?!�A?�(�>W='w���Ƚ�&��-=��>bY>@�o=���=F�� �Y�I�,H='R�=N�Լ|@���	<d��^6C<�Z�<�Z3>��ֿ��A�V�ݾx����߾,��_�����Ž��e�������ϒ�G]x�x).�%��[`���f������qO��N�?h��?fЃ��&>��=��`��&
�,`�>�t�E���ۺ�}L�9>��3񾬗��+����L���e�:�Q�S�'?º���ǿﰡ�
;ܾ! ?�A ?>�y?��N�"�ǒ8�M� >�G�<�(��l�뾫�����ο3�����^?���>��/��`��>��>��X>THq>����螾P/�<��?K�-?-��>��r�+�ɿ`���i��<���?!�@��A?��*��Pʾj��=0y�>H�>��>'�9�uP��A���<�>,�?� �?�w�=��Q�/V���P?O��=�P��"; !>�Q��G�g<����~0>U	�>m��G*;��8-����=��S>Mu{�������6���ǒ4>��W��L�=-҄?j\��f�`�/��Q����>��T?�r�>�@�=D�,?�AH�rϿ��\��a?l/�?���?\�(?�쿾��>B�ܾ�qM?�56?UΘ>e~&�p�t�t��=�Y߼����a�㾌V����=e��>��>�w,��s���O�/4��]��=@��������d&�8M��ѡ=F��;�p3�Eս�S���=l������.>�t�ݽ.�=5��=�H:>�ɀ>�#h>?�Q>��[?�m?e�>E�,>������ξ�ZԻ���ǈD�V����0C��V���y��9����o���X�yI���=�h�=�7R�Y���"� �t�b���F���.?g�$>!�ʾ��M�qR-<�mʾ����1���ƥ��.̾z�1��n�~˟?��A?����/�V���/��a��P�W?t'�����ի�=����-H=�&�>���=p��3�{S�St0?yn?�`��Ax��.X*>tE���&=��+?v?�VZ<�Q�>z-%?�+���нZ>��3>�s�> �>c�>]*��2�ڽ�?�vT?�T��0�����>ec��I={��`=��>o�4������Z>#e�<�x����Z�z�����<�(W?՘�>g�)�-�0c����|W==
�x?ߐ?f*�>kzk?��B?�B�<Sb��/�S�4 ��?w=��W?)i?��>Iy���о����5?g�e?V�N>jYh�=�龏�.��U�� ?��n?y^?le���u}�
��b���s6?��v?�8^�a�����iV�Z��>�m�>���>g�9��f�>�>?��"��I�������^4�ʷ�?��@>��?�37<B) �@�=�U?�h�>=-P�~zƾ�ɳ�Ⴕ��.o=���>q=��_,v�����,��@8?
l�?�F�>�X��G����=�T���U�?��?�o��U$o<���l��@���Ȣ<�ά=;d��a#�>��8�2ǾĐ
�ā��4����`�>RL@���sS�>^�7��3⿟VϿw
��%о�q���?5?�>+ȽI����j��fu���G��I������5�>���>Pa���<���Z���*��=�Q?~�����=V���
��O���	*f=��>�/�>ht�>p�ͽ0����?��dÿ����1N+��\�?���?Z��?��+?:V���rҾ�%�ߓ�=�;_?^R�?BRb?8\���/����j?�]���T`���4�HE��U>�"3?$B�>7�-���|=Z>���>�f>�#/�8�ĿAٶ�m���?��?K��?-p����>~��?xs+?�h� 8��	]����*�kY+�f<A?�2>E���ظ!�0=�eӒ���
?E}0?�}��-��5]?�eR��@x���0������>��z=��s������C����|��(����C����?���?�^�?�	C�d$*�+w4?���>��čݾK�ｪ.\>7ɽ>)~�> �G=q�)>�{#��g=�p�>���?��??�?�ؔ�����}��=�7h?d$�>��?7��=od�>hv�=A氾[F/�JV#>�3�=x�>�%�?J�M?i=�>���= $9�J$/�ISF��GR��"�Y�C�!�>�a?P�L?	Tb>tX����2�4!�Vbͽ�U1�((�Md@�D�,���߽F$5>��=>�>�E�AӾ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Da~����7�0��=��7?�0�$�z>���>��=�nv�ݻ��X�s����>�B�?�{�?$��>&�l?��o�Q�B���1=.M�>Ҝk?�s?�Eo���:�B>��?�������K��f?
�
@~u@`�^?(JRԿ5���ʸ޾o�߾�UN>ho�=J�1>�G`��,�=?�k>>&>�
=���=�{w>3UY>�1?>>>�S>V��=���t�`������S#F������@~����׾j)�T�⾬宾��о�B7�ޭM��u0�ǌ^�*�J7�����=/�U?R?Rp?Đ ?�x�"�>����j�=^�#�˄=t*�>�f2?}�L?=�*?K�=������d�*_��A���Ƈ�3��>zmI>l��>M�>�$�>�9��I>�5?>G��>�� >�N'=��h�=�N>�M�>W��>�t�>~K>E�>\B��f㱿�	f���P���E�ۀ�?��y���J�tD���!����i͞==�6?�� >�f��eoͿT��*tA?�]��9���D�.�w=1?z�X?��6>�-|�Bπ�W�>s���`l����=1C����M�2�/�lZ>�?uMg>�u>��3���8���P�zί�6�}>|�6?ez��G3:�H�u�'�H��mݾ��L>oZ�>�(����얿h�~��+i���z=DP:?�D?����좰���u�5�����R>�"\>�=��='L>�e�pƽF�F�X�.=?��=�]>�O?�X/>�p�=۹�>kҙ�N�l��>�>A>�Y*>;u??�%?���ݚ�#���|+1���t>a#�>�3�>��>��K��ɲ=
T�><c>���b����v��@��[X>A�w��W_���y��wy=ﭘ����=�ˍ=�����A�\�!=�Ty?������n���z��Z=!?�N0?�d>+Ž�B�0������m��?m-	@�{�?F��CM� \?�?�*��-�C=���>���>`h�^픾RN�>�0t���Ǿ���Iڈ����?0�?N�̼ ��J~�ަ<q�<?���Qh�>}x��Z�������u�K�#=O��>�8H?�V����O�c>��v
?�?�^�ߩ����ȿ6|v����>W�?���?e�m��A���@����>9��?�gY?|oi>�g۾C`Z����>λ@?�R?�>�9���'���?�޶?د�?XO>[H�?���?v�? ��Z
�v���i���m�D=�U>~_>��=vZ߾u�m�g����ݚ�CW�hJ��1>(ƈ����>�\�=�[���'=�j�����K6m�6>J��>/U=2m�>D4�>���>��i>�C���Z��}x���!�}�K?��?k��J3n��.�<!��=E�^��'?UK4?�[�$�Ͼ�Ѩ>�\?���?c[?�g�>���K>��Z翿*}��;��<�K>o3�>�H�>�&��1AK>��Ծ�8D�jp�>�җ>��.AھG+���V���C�>�f!?���>ή=0� ?ߚ#?�j>�0�>?bE��:���E�R��>���>bF?o�~?��?lʹ��V3�����塿֑[�ON>��x?�V?�˕>����ނ��7�D�u$I�캒�e��?|og?x形 ?�.�?.�??��A?g<f>���׾>������>:�(?���S3K��>U�첲���?+�:?��K?��
?�b�������5��K	����>�L�?7o?�n1��2m�$a�.�=��4=d/K=���<�0����=��ü�G˾��S=k0>���>�ٹ�v��-�r�h�=��>�C�>Nf�L��**?�%>��%��f=�6\��L	��`x>�2 >Y\��%�S?7�p��/U��|���r������p?5o�?�?|߽�d�+>?-[�? y?0¾>H����p ﾫ�@��C�Kq���=�J�>EA���ti����������u���,�?#�>���>��>��>�>����u+�������c�d��x�P��q	(�������r
Ͻ1U�;|&ž��w�3�>^��l��>�?�d�=��2>���>�B>�R�>.WL>H�>*�e>e9o>�O>�ʏ=ҋ?��U$�|�Q?@>վzE
��΢��cƾ���>78J?jC�>��d��艿H����H:? �?�.�?X�b>;k��';�]�;? b?f���?�=�<�P�<�>�Ԣ�����_ɽ�U�X!�=o�R�QzI��<_�:NI��&�>�?�\�=�w���h>���3�=8�u?؍8?�C&���b�@o{�_�V�J�E�G�������!�Nu���������gځ�Iw$�T��=^?>?�O�?'��i,���]ξ�Bw�
�?�0�E>�J�>{��>���>�	�=���pL,��MQ�����Oe��r�>��z?G��>o}I?��;?=�P?�rL?�>B�>`��k�>'��;|��>��>��9?B�-?�.0?'|?}�+?��b>|#��y���3cؾv?V�?O?�?4�?����<ý󺗼Q4c�X�y��� �=6W�<
׽}#t�$�R=~�S>Y?����8�����p k>�7?���>���>L��p/�����<V�>�
?�H�>�  �=~r�c�QW�>c��?)���=��)>S��=k����ӺS�=����\�=�9��lu;��f<�~�=��=��t��~|�.i�:�χ;�f�<X�?z�&?v̅>�Hf>��b��������fm�=�I>2�X>�an>����Z���������i�1�y>Lq�?�?�s�<05�=Zo>R�Q�}��� ��[�)f���>o<?glD?V��?��<?�C#?��}=��!��ݜ�հ��؂��3�?�%,?^5�>u����ʾ"꨿c�3���?�\?wNa�0��aN)�y¾޷ҽ�q>b//�'9~�_���i�C��~�����ߞ�����?U��?.�=��6�,���ʘ��i��DmC?�>�W�>���>�)���g����;>��>g�Q?�A�>���>�{�?��q?oss��IF��_���������s�y>�5\?�f�?aj�?|?��f>Ƨj=��*��Q��k���؍�j;־:��=�0K>�]->" ?(l�>�>c ���Kҽ��P�7>�c>��>Β�>���>��>��=�J?$+?2�˾��#�0{�tÏ>+"�=�J=?�6�?��$?(b+>�G7�Ygj�O��H�>M��?���?]�>�蒾��T=R�]=��7���̽ ��>d`?��|>�R��#�_��Ə>ņ�>Q�
?�#���.��zh�8���6?�k?�EE;�ǿW�r����� [��ƚ�>͝(���F�G�O����p�5>���xk�<zC���1o�{���P̈́�U0��ܵj������(�>���=�ߺ=OF�=�H+=(=��	=�y�=�ߴ<}3ϼ�ŽSm=?x���9��&��s�;R~�=$/�=�^E=�̾�}?��H?	\+?��C?��y>��>�7��M�>i���?��V>ګP��e���;���������hؾGG׾Uuc������>��H��V>�3>�"�=:�<E�=�s=���=��9��=%!�=���=���=W��=��>>b>�6w?V�������4Q��Z罢�:?�8�>y{�=��ƾm@?r�>>�2������vb��-?���?�T�?<�?7ti��d�>U���㎽�q�=Y����=2>���=c�2�P��>��J>���K��(����4�?��@��??�ዿТϿ4a/>�7>h8>ؿR�U�1�.�\���b��}Z���!?�H;��Q̾='�>�ͺ=�/߾��ƾ9i.=Շ6>�nb=4_��O\��ϙ=��z�	 <=��k=&Ӊ>��C>�<�=)@��r�=J=k�=��O>& ��5�7��,�
�3=6��=��b>�%>�7�>L�?�l-?�jz?���>����|6Ͼǒ����=��;��>G"�d�->��>Rv0?PTE?�e?o%6>7C�=x�>n�>�(�Ue�ś���,B����=���?s-�?j�>�]�=a]����7�,����<C?J`'?}��>�05>�S�*����$�;C�hW�>�&>_��=l�B=j]�>"xC>d�>�d�w=!�i>��=���Z�]>��<�7�>2�>1�S��ܭ=�B=�<Ǻ�>�4�����$�]���=���<��<k̼(��<m�<?�y=+t<�J�=�P�>��>�z�>F�=v�����.>d���m�L��+�=T>���B� d��?~��#/��6���B>�aX>�)��o)���?�fZ>6�?>�d�?��t?��>�~��Rվ� ����d��S�� �=xI>�$=�w;��N`��N�MoҾ�O�>Yg�>���>t?o>�`+��f?��u=xH�L�5���>�����}��a���o�פ����� �h���:3dE?*�����=`}?��I?7�?��>o���-ؾ�{,>�\����	=���8t�' ��v�?��'?�2�>���D��p���@�<xK�>�ٖ�̖Q��䞿�4C��s|�~���h��>sU¾����1�㌇��둿J{?�P�w�
.�>E{^?_��?�$9���w��(F�|������?��l?�F�>4��>�V�>㽙�������f>_s?4��?8�?��> ��=7��Y:�>=,	?q��?���?�s?t?��u�>��;q� >Ř��C�=��>���=�3�=yu?��
?�
?�g��X�	������q^�r��<:ԡ=�>�n�>?�r>���={�g=rr�=�*\>�ڞ>��>[�d>��>�M�>jʈ��ھ�>=?i�<)�.>�?l9�=c�f;ў/��f���}½�a��lf�2R��k�½��u<��T�N��=T��%u�>Z�˿V�?L^>�=�'�?'����J,;>���>��t=#u?�ؗ>{��>�>Mu�>}b�=�;�>|(�=�%Ӿ�J>���kK!��3C���R��Ѿ(_z>q���&��������H�bJ��Vd�;j�0/���=�c(�<B�?�7��K�k��)��C��V�?��>�(6?�Ԍ�¬��]>��>���>4������č��oΆ�?0��?�lc>�*�>ػW?&�?��0���3�cZZ�Eju��OA��e���`��׍�����C
�����_?��x?-A?P�<I�y>U��?ƭ%�{����E�>�.��;��>=�!�>
����_���Ӿ��þ�b���F>��o?z�?��?6BW�m儽�`">�9?�1?N9u?W�1?�:?�p��!$?�(3><5?�	?h�4?��-?l
?Q1>�O�=�#����#=�{���T���DϽ>�ǽ������2={!x=��:N<�r=B�<+4���Լ���:Fխ��/�<Z�F=@Φ=~��=���>�]?�@�>�Ƃ>�)8?F��x�5�����BB.?��>=��{�K���զ�V���� �=��j?`�?��Z?��\>$D�Ff>�ý!>���>�P>D�U>�̯>����P���u=p�>�� >���=�	z�-���+��-j��W�=Φ>4��>�4>���~�$>����{��d><WQ�$N��:.Z��TI�0
2��u����>o�J?�?߳�= ��;���?f�M�)?�G<?&DL?��~?��=uܾ3�9�:EI����I�>���<� 
�@���T����[9��9;�Nq>�%���ݠ��[b>A���r޾��n�J���羋2M=���OPV=��� ־�:����=_#
>h���� �-���ժ��/J?ڢj=�q��@_U�r����>潘>cޮ>��:�6�v�܆@�#���v8�=}��>��:>�o������~G�A8��Y�>	E?�\_?w�? Y���
s���B�����\��G�¼��?�ȫ>{�?�B>���=F�������d�(MG���>MT�>���G�QA���F���$���>H?��>U ?��R?�?W�`?��)?q?kb�> T��J���B&?r��?�܄=-`Խ�sT�9��F�� �>2p)?��B�mɗ>H�?��?�&?-�Q?�?ԓ>Q� ��0@�L��>�L�>��W�c��[�_>��J?`ϳ>PY?�҃?��=>�|5�Ԣ�����)\�=��>�2?�'#?@�?_��>��>8���y�=���>�c?�0�?$�o?J��=@�?�:2>J��>���=���>N��>�?XXO?;�s?��J?��>��<^7���8��Ds�T�O��Â;tH<��y=z���2t�|J����<�;Ii���J��&��z�D�3���%��;��>�:p>h���$>�ǾJ􄾙^I>&b��p~���ы��KH��R�=��~>��?O��>�r�=�/�>��>
�%M&?5?)�?�B�9Cc�ǻ־�<��}�>4�@?���=�vi����S�x���s=xZn?/\?)�Q�������b?"�]?@i�=�Y�þ��b��p�x�O?R�
?k�G���>��~?9�q?��>z�e�3>n�"��9b��j��Ŷ=�p�>�X���d��3�>w�7?�O�>�b>�v�=it۾��w��~��L?K�? �?l��?�9*>��n�2�q��퟇�	=Y?j�>�M���?��j��;þ7ʍ�����Wnľ~�󮱾�U��/����t!�5�u�����kU�=�=%?��~?o^_?ͪg?�o���Oz���c��?n���O�y����tA���=���G�M-f����V8����h���<=ȉ�XUE��4�? �3?m^����>/�,�K��{;�>	J��R�����P>�F =+��=�x�=ʨ����K!񾭹'?�'^<I�/>�Q?G�O��t<���O��EK��9���>�)?f?+�M?Pa>�@V����>���-s��c��k/v>p{c?��K?��n?_b�+*1�������!��0��f��S�B>;7>v��>��W�����2&��R>���r����2u���	���=��2?{�>O��>�G�?3�?js	��^��hOx��x1��c�<�2�>i?:4�>
��>�н]� ����>:�p?L��>��>꤄�g��|��ֱ�r��>ש>���>��d>�15��Q^�
6���ǌ�&'9�j��=Gd?�e��2�S�hK�>qT?KI<�E�<�B�>������,R��-�L>KE?y��=��5>��¾���o}�����U�)?Z<?_ʛ��@3���f>�,*?�"�>h�>���?�>h���3�Nl?xb?4P?�@? 	�>��<x7Ѽ�ͽ�S)��?=��>�-<>uyY<N>�= ; �1�i���A0=��=�xz�=��kC<`��<�<�#�<��">�BٿWC�<�ʾ_��FھU���������:���=�"u��di��S���̚%�p��^�ݐb�l���2\�v'�?�D�?f����tu����S_��ʫ��)�>9`w�Ѻ �!A��ń��;�����o2��w8(��N�*�]���`�Q�'?�����ǿ簡��:ܾ)! ?�A ?5�y?��@�"���8�N� >�C�<+����뾮����ο�����^?���>���/��L��>���>B�X>Iq>y���螾0�<��?6�-?��>��r�/�ɿ_������<���?*�@l�>?��9���ľ��O>��P=�SV>i����l�ȝ����?LǱ?��?H*a>l,D�D����S?8,>u	��+�<�d>(aE���t��l�='<#>F��>�>T=�獾��Y�Ӿ	=�A�=Y��^��8��p�c=�@>��!>H_�>:+?B�K�v�hvD��M���D�=d9T?���>eE=g%?��Z���ɿ�K��XW?(k�?�q�?R�,?�޾�è>>�޾�w.?P9?>7��>Ã�@s=����2����\.W�"`�=Ot�>=[>��Q�U����ɾ�='>c���)ƿ��#�����=婟�7�^��Y�N�� �Z���9�l����V�^=,��=��P>� �>[�T>�[>SW?4�k?%6�>yi>`��`�����ξG�ׂ��}�GQ��9��`���y��߾>c	�kh�C��H�Ⱦ!=�n�=w6R�䗐�t� ���b���F�p�.?�u$>Z�ʾG�M���-<�pʾ���;愼H䥽/.̾��1�p!n��͟?��A?�����V�����a�����n�W?�P����ꬾ���=9���|�=�#�>n��=3���3�2~S�iv0?�Y?,}���P����)>�� �Ê=��+?�?�^<P*�>^6%?�+���ʌ[>�4>Nޣ>��>-F	>����ڽ��?^�T?ڔ�`���,��>[P��{�T=a=�n>,5�:��)k[>m��<y���bU�� ���g�<��V?s�>��'�����V��}G�I=��w?�3�>O�>��k?r�F?B��<AB�EOL��k�D�=��]?�,i?p�	>�膽a־�����,?�8i?Ǹ>r�5��^ݾ41����.�?��n?�?�<)��#|�kc��{j�G�0?	|u?-�Y�������l�a�W��>��>qT�>�;��ߵ>+�<?�+�rz������y�3����?.�@���?�� <��㼳J=�O�>9�>_�N�O_��ݒ�}_��}��=���>d/���*x����s�$E?��?7� ?6W�����a��=�˕�oZ�?��?x}��Lg<���l��i��{�<cϫ=��-R"�h��D�7���ƾμ
������F�����>�X@�F��1�>~58�f2�8RϿ#���Sо�Zq���?��>&�Ƚ}���P�j�yMu��G�D�H�2���
\�>M�
>>Ɨ�A���r�F;��p��Yn�>MC��!x>~B��������?�=��>5�>�t>�]��o��R�?|���gPͿL%��]O
��Z?�B�?��?��?G�»�jt�-Qo�  b;a�D?v�k?SCT?��B�z/O�5�P�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*�{�+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.���_?��a�@q�(�-�K�ȽE��>�M0�1"\�u���2��\e�H���py�?�?�]�?A�?X���#�v&%?y��>����r�ƾ���<�l�>���>��M>oS`�?Vu>��	;�G	>���?hx�?X?����`���+>�}?Z6�>�ɇ?�J>���>:Q>�2����漆�0>@��=�Q��� ?�*G?���>���=�R�",�PF�m1T�����B�b�>�Pb?#P?0Ro>�j��d`���$����1�5��] ���1��X���۽+->Ds<>� >�n]�Tʾ��?�o�2�ؿ�i��2q'�"54? ��>�?C��q�t����;_?�y�>	7�,���%���@�`��?kG�?��?�׾�b̼�
>��>K�>��Խ����������7>�B?���D����o���>���? �@�ծ?@i�N�?��ؾ󶐿�\w���
�U���=O0?N!
�/��>D��>�*G=��w�䨢�g��T�c>��?���?��>��v?D�v�v7T����v�>'��?��$?U����DJ�=��>��{�������߈r?Y�@[c@�W?�!��v<Կ�W�����������=�9<Wk�=r�G���=#�=��=?&#=��=�K>5�>a�_>T�b>0>j�>k1~�������d����}9����H< �뫒����J2E����x���9٭���2~�y���u�����͈�ػ�=_�U?dR?��o?E� ?��y��t>W����z�<�#��M�=�Ն>�32?ΎL?=�*?�ޓ=Ǒ����d��R��6���ㇾ���>s{I>�#�>v�>M��>X�8��I>{B?>p��>�P>Q�(=�ĺ�j=��N>�-�>���>K�>�C<>��>Cϴ��1��o�h��
w��̽3�?5���L�J��1���9��ܦ���h�=Qb.?|>���?пX����2H?���k)���+���>k�0?�cW?^�>��b�T��:>3��˦j��_>�+ �Ll���)�{%Q>al?t�f>^�u>�3��8�FXP�E+���c|>W�5?�����h9��!v��H��޾NmL>��>��"��'疿L~�B0j���~=�";?�?�鳽���� �u��᝾H�P>�;[>I�=���=�L>�f��(Ƚ�DH���,=���=��\>f?�->T�=�>-/����P�	I�>�>C>��+>"@?_7%?�o�^�������	p-��$x>N��>�o�>�K>��J�d��=�x�>Ob>���HY�����˰?��bU>�����_�us��Hv=�x��b�=~A�=��\=���+=)�~?�z��&∿t�@E��^lD?�+?l�=�LG<H�"�E���aE��� �?&�@m�?<�	���V���?�A�?�����=�l�>6ʫ>�!ξȓL�,�?W�Ž����ˑ	��(#�P�?��?oS0��ǋ��l�X2>]%?��Ӿ-w�>#Z��P�������u�4�"=��>�AH?|r����Q�C�=�N�
?B
?��!�����ȿ�v��<�>���?i�? �m�/A���/@�(��>���?��Y?�/j>�۾�{Z��_�>��@??R?_��>FH�Ȕ'��?I϶?s��?BWF>���?��?d+'?|�=��Ͼ������b��zO>�(�<�52>�M�=����V�q�2��9Le��R����c�؊F>SѼ
��>A^*=�U���
�'�ۼ�cm�#�u�{	�>�h�>�G6>�ƺ>60�>��>��>�⾽=$������H���K?���?/���2n��M�<x��=�^��&?�I4?vk[���Ͼ�ը>غ\?e?�[?0d�>>��L>��;迿0~��֪�<��K>44�>�H�>%���FK>��Ծ�4D�xp�>З>�����?ھ-��0S��NB�>�e!?���>YҮ=J� ?O�!?d�f>���>tT?��Ƒ��BD�z�>��>:6?��~?�B?����cs-��q��?��_�\�Y.a>��x?^?>ꗏ�dם��¼�e��>5�D��?V�f?bz����?ﰈ?��??�)@?J�W>���+پ������z>�&?���G�pW[�<��t(?0h+?_�?
�>��r�����3��]¾\�?{T}?9;E?R����4�h�=��J�@�������=ƿὢ��M�G>�>6Շ>���>M<$>��Ľ%���!z뾇��=Z?�M>ζ��;���,?_�=1d]��Z�=8�j��8����>,�>w��Cu?7��x�w�N姿�|��a�\�xe�?���?���?�8��<a�jD?Ӏ?e�?4R�>X���,L���Sޞ�x�ƾ���Rt>5K�>9F�����剨�iT�� -|�vdŽ�����<?��>g�?5%�>���=�|�> 3��oT:�r��B��l e�x�&��,/��&���Ij��6X��x,X�ri¾�a����>���;geu>p�?�m>�`>�c�>�-�����>D�>8��>Jz�>�/>6�>���=����+�FI?H��\,������s���?�x�?4�$?�3�=~�������D?Q؊?6ޡ?�u�>���42�J?j�?V�?�O��>S]���þY=��Ä�=.d��ړ��ԙ>�7e>V�⾪�w�9	�-%��]?3
?��=�����=�������=��?��-?�h�S^��Pt���K�]�L��Fr�~�[��̗�(H&���s�4H���3��%_�����Kw=�OF?Y�?�K��v⾢�Ҿu"t���7�	��>�d�>`7�>.��>��>��	�3X/�[]��R9��Ȁ�C�>�j?��>HtG?d�:?!jR?�)M?�։>i�>pN���+�>U?�9=��>��>��9?��.?U�0?)�?��)?}n>]޽v���)�Ӿ-�?D?P*?�J?�z?�t�f�ͽ��ؼ�?I�NPv�Ɨ��q�=��=��K����Y=ob>Q	?��b�7�z��2_j>�=?c��>���>�僾7X��I鬻�3�>'�?
��>x��L�n�oq�ƕ�>pL�?���!	�<Ab(>���=�yI��m�����=��՞=ħлR`���;�C�=�y�=�������<x�X:��
���=�}�><�?)��>�:�>OR���� �:���=5,Y>O�S>�m>�Tپs}���&��:�g��y>ay�?u�?k{f=���=���=k���Q��������i�<ݐ?-.#?36T?���?��=??e#?3t>D��P��7]��^��+�?s!,?���>�����ʾ���3�ʝ?1[?�<a�-���;)�r�¾B�Խk�>![/��.~�n��.D�yׅ�����}��&��?ٿ�?�A�k�6��x�Ͽ��r\���C?K!�>�X�>t�>�)���g�b%�b/;>3��>DR?��>#�>�NV?���?�Wp>�4?�W�������(�@���a=�PH?���?��?%;�?�D�>!�K$�1��.���d�j-����Ͼ7��0�>��^>j��>��?@�=����p�=��=�~�=8��>��>]I�<�S�>@��>�6�;�YE?��>��H���E>Ѿ�ZN��w>Zj�?T�?]�L?/�=��(���R���7"?�e�?`�?�I?��2��^�=̞">z	��B�����>�gc>�Q<>�(�<�E��� �>�2B?j+�>�+�& ��=�ķ"��;?�D?�|k�� Ϳ��n���ýr�s�x��>��:�-�J@����.�=��<��;�j��,	��	~��*����S��᣾�g�3�>\��=U\�=BD�=���=��1uC�e�>�y�ȪŽ�ټ�r�;#W�����+�d��:L<.�J<��<&�A<�ž��?�[Q??W0?�GB?;�>[��=�P�8қ>g.W��z?�HQ>󣖽�̾�[�L����lE�r�оY�c��͠�H�>�Dw�XG>��*>N�=���;��=���=���=�
<�{=uN�=Aӽ=Kǃ=���=�_>�>�Uo?��b����,pW�(Pv���,? �>��=��dQ9?Le>��(���!��w?���?D��?���>�S�)��>�;s�ۼ&��;�8!�z[�=��	>�C��B�>u~>�U3�6��G'g<�V�?o�	@�O?������޿C1>έ7>#>�R�߉1�"�\���b��|Z�ޛ!?SI;�UJ̾M7�>��=�,߾�ƾ�.=C�6>�eb=0i�vV\� �=9�z���;=�l=�׉>��C>\u�=b0����=f�I=���=d�O>�:����7�&.,���3=w��=p�b>�&>��>AN?�.?VOe?�	�>�s��wξ�����7�>. �=���>I�=;>D>`%�>>�8?�@?BWG?<ɹ>�Ù=�^�> b�>�n-���n��m羲����-=]$�?�@�?F�>�Hj<d�9�'��_<�zսM?�$.?�(	?Y��>�E�¥ɿ�)۾�E���S>C��T�u<3s���3:�U�=�ت=T9�;�7�= _1>�>`%�=�W>�uû	v�=��>˿�=-�g<���<Y)�= ��<&t���=�k&<��>�W��;�c�<{U��BWU<�=q�_<Qg�kh!<[(=��>�??�^>:�>ﭹ=�ܝ���=���{�0��k�=���0�B�o�c�{�����?��,�^�>=�>�C�_F��0�?T٧>��>7��?>j?aq(���R���Ӿ�����������=x(�=*ו���;�W:o��{l��Eɾh��>[�>r	�>��l>E�+�! ?�0w=�⾴a5����>�r��^����-.q��:��WG	i��KǺ�D?�B��|��=� ~?�I?_�?r��>(7��\yؾ�0>oT���x=	�yNq�o&��?I'?t�>}�ԡD� #��<��<�r>���?@������6��YE=aȾ��>́�F���
z9�񝆿3㓿8�c��Xx�&��>.�@?��?��p�s�����g��4�h+=(?�Hc?Ӛ7>L)?9	?�ǽ'n��O�ɮ���WK?���?�%�?9)�=y�=1)����>�M	?u˖?.��?Ls?�8?�@��>а`;�-!>M䖽ȣ�=Ǹ>Sם="n�=#+?f�
?w�
?5����	�E �x7�3[^����<[��=M5�>.��>C�q>�@�=`[i=��=/Q\>�}�>у�>|:d>�0�>��>!j��j �h�E?տ�=IHR>B�?��N>�$��e��#�<���{�dQ�K�x�\q����a=Rㇼ�cp�k�I�<x�>��пۙ?3�>@���t?0�D���>�"�>� f<��	?*��>埨>��>W}�>���=iz�>�Ǆ=�Ӿ�G>����~�<5A�ЕS���Ӿ^Dy>���3�&�q�i^��B�K��A�����(.j������Q<��J�<M�?�
��l�d�)��\��?m��>b6?�F��kq�I�>���>�
�>[��nk���1��dw���?���?C;c>��>(�W?Ś?&�1��3�}uZ��u�,)A��e�Ѽ`��፿�����
������_?c�x?�wA?�O�<�7z>��?��%��ҏ�b(�>�/��&;�P><=�*�>z*����`�5�Ӿ�þ~7��GF>��o?�$�?MX?)UV��p�,�&>b�:?\�1?/ct?%�1?�t;?d����$?�S3>G?l?�-5?��.?c�
?�1>��=�I���7(=�Ց��Ί���ѽ��ʽ���-�4=aV{=,��8{)<kr=r��<NY�d�ڼ94;�V�����<�M:=�ʢ=��=��>\;]?��>�ڇ>��7?<�O�8�����
@.?��5=�'���2��{������8>̅j?[��?��Z?;8f>#B�.tA�$�>��>�(*>��[>�>�w��~F�P<�=�r>+p>o�=i�E�_����
�(;����<l�!>��>=�g>�6��E:�=Qȉ���̾�)]>����-
�Ԃ㽾�e�CI�Vg����>�!B?��#?�ٕ=2�ھ=tF;v8o���E?Ρg?ՃX?g��?�i!=0���D�^Z�����n�q>���<����;���S��X�2��"���7>�ͬ����8 d>�m����54q�`J�cྒ?�=k��2��<���J�ؾ������=j�	>\R¾��"�N������L?�]�=㩾��H�j����>�U�>( �>�Qͼa����CD�0~�����=br�>�6>�8ʼl��s�G����)�>2�J?��]?��?<5~���u��mH�ʿ �E[���0�E�?�h�>?W0>
��=wk���V�V�c��F�z��>�_�>Z$��=B����x����\"���>�N	?�>in?��T?5�?�]?�/?�Z?�ғ>�;ɽtžk�$?�
�?	Y�=����]�V�� 5�͆B����>�)?�.�/ܟ>Tq?�?��'?C�S???�y.>�3�HA���>=��>�2Y��Z��Ze>BF?�ò>��[?Oڂ?:�6>�U3�v���V�{�=`M>��.?ʼ#?�) ?ž>�D?�b/�{��=��>��E?No�?4J<?��=�{>?�R�>{� ?�d��>.�>R�?N�P?�^z?��K?0`?᣽h�2�l��y�q��%�<r��<�=�=-���<���������v���d��,8���<�&Ľ �ýĄ�=�_�>��s>x
��)�0>4�ľ�O����@>n���P��Fڊ�̎:��޷=���>��?���>�X#���=;��>sI�>Q���6(?��?�?@�!;�b�M�ھ�K��>=	B?���=��l�������u���g=��m?��^?g�W�p&����b?��]?�f�=��þ׺b�֋�S�O?��
?j�G�V�>r�~?��q?���>m�e��9n�����Cb��j��ζ=�q�>�W���d�0@�>n�7?N�>�b>�+�=[t۾��w�vo���?Z�?@�?���?�,*>R�n�[4��h���H��u^?�o�>�j���#?�4��ϾjI�����������{Ϋ��o��3m���$��僾�ֽ�s�=x�?7s?Eq?�_?�� �md��.^�����^V�u2�^!�$�E�P E��C���n�Z{��>��0����H=�YR��`��-�?|��>���?d�˾U�,�Ѿͼ�>��?�o&2�\ ]>0I�i�=�>->��_��~����׾��?*�?u�>��e?���xR��H�Y}C��nþY�&=M<�>'F�>|g*?u)���6n���!�aG��_�� �.�>��u?�	F?��u?a-���E��w����!��I�Y6��T=m>�h>�a�>�pM�����)��z�3�� v��p'��*�����h��=�*?SS�>���>9��?��?6\뾐����vp��b���J<���>�{y?���>�õ>[����2����>3�l?N��>�%�>ҧ��Z!�S�{�)�˽C��>\ҭ>���>��o>,��\��l�����\9�Z�=��h?����Zt`����>b
R?S��:��=<�U�>K�u��!���-�'��>}e?�˪=��;>(mž!��{��<���G)?�(?Ų���)�(�~>U"?-��>d�>��?��>\���_��{(?�0^?�?J?�_A?���>�j5=~T��"�ǽz&�>y=;3�>�1\>�){=\H�=��gS]��� ��>=f��=j�ۼɽ�0F�;>����3<��=pK7>��ݿ�;J��оS��,�Ѿ���daw��=�1����p�`Ⱦ�����u��m�(�����Qd���u��Sr��]ɽ�P�?��?l���췾5�������uL7�S�#?�j��m��{���|i�|=ҾQm���u��x�I�ha��lq�g�i��3?�?o��YԿ|���¾�Я>)L?�(�?zp#���;��,V�b�>�P"��3�=����J��*ʿkE�̹;?�<�>����2d<b��>�o>�4W>��V>O���>���H��>�;?HH2?*��>.ɸ��:¿%����n��m��?��?}A?�(�����V=1��>0�	?��?>�S1��I������T�>g<�? ��?;|M=`�W�W�	�,�e?x�<��F���ݻ�=\;�=PF=�����J>xU�>(���SA��?ܽ;�4>Bڅ>0}"�?���^���<k�]>��ս�:��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=$���ƿ�;�]��mP�=3��<S콽�����ӽͻ-��N��g^v��י�f0=�>�o>D��>��X>;+�>��]?VEs?���>]�=������������=����Zp������K4�{Ż�}��R���4��E,��i������B����=(=\��ʒ��V1���`��Y���P?Wr�=�8�� W�s�����G��y�Q��M��R���?�@kW�/�?^_M?�/���+?��3��2���s�=ƧR?{�X=���_����=5�����9>��>=ƙ<�&���R�>�i��l0?MO?"�������*+>����x�=��+?��?`�a<V�>F%?�+�9��n\>�4>���>���>?M	>t8��s�ܽkR?)@T?5� �	X��W�>=�����z�cXb={n>��4�s���[>|y�<]���K�P����*�<�(W?���>��)���Qa��s���Y==��x?��?'.�>_{k?��B?kӤ<�g��6�S���:ew= �W?*i?��>,����	оf���H�5?�e?��N>�bh�#��+�.�IU�g$?��n?�^?$����v}�q��B���n6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>��������>�vN�&�?)[i?T	�[�>Q=�x��-3��O�=/�P>W���N>����?8�/�������>J�S����%5>Z�@	j��9T%?в�NlΏ���1}z�,�H~��6?#�m>Մ��	"Ž;؈��N��u�A��$\��ȼ�@�>��>���e����{��r;�t���)�>R ��>��S��0��դ���6<p�>���>���>���� 罾�Ǚ?�P��M@ο����)����X?^h�?wk�?�v?&�7<Lw�v~{�ʈ�1G?��s?Z?�%��Y]��\8�=i?�����c���&��*B����=[F?i[�>318�W�^�Xk�=��'?���<D>��οd%��\��X��?�R�?԰ �( �>M�?��3?�W
�&���F��2V�c_׼�m?FTR>2�����ڨ\���ž�{�>%?o�^�[MҾ]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�$�>b�?���=Ls�>Xy�=����\2��E#>j�=�?���?��M?1H�>� �=��8�`/��XF�~HR�$+��C���>	�a?�|L?�`b>:;��02�f� ��ͽ�L1��꼨 @�1�,�
N߽�p5>>>�<>��D��'Ӿ��?Lp�9�ؿ j��"p'��54?1��>�?����t����;_?Nz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�>=�>�I�>B�Խ����]�����7>2�B?X��D��u�o�x�>���?
�@�ծ?ii��	?���P��Xa~����7�_��=��7?�0�(�z>���>��=�nv�޻��V�s����>�B�?�{�?��>"�l?��o�L�B�P�1=2M�>͜k?�s?�Oo���m�B>��? ������L��f?�
@~u@b�^?*�hֿ����_N��P�����=���=Ն2>�ٽ,_�=��7=��8�C=�����=t�>��d>"q><(O>a;>��)>���Q�!�r��\���S�C�������Z�C��Xv�Xz��3�������?���3ýy���Q�2&�)?`���=X�D?�D`?o��?��?�(��������s���ܯ<���>7_�>��>?��U?M�O?T�k>;���ꁿP���J˾G���T�>�,�=h�A>*J?�j?��^�w�>u@^>�և>�̉=fIO>�3輥Յ=��k>�C�>�s�>)��>Ԃ*>�-|>Ԣÿ�W������j��;�>S1�?��=�4���)�������h��>��>G�i��.����ɿ�拿#&Y?��|����E���>��>��4?��=�MǾ+f">�=�l>Z;���='�2ț�V�����>�'�>�b>�z>�m7���5��V�/��e΅>�;9?������Y�TE{�hF���2a>��>�#弈m��Z��g}�ybY�}=�@7?cx?�%��G{���m�����Q�Y>^7_>�<�f�=
�J>09:�J�ؽG�T�b�^=qn�=�e>�`?�|,>)�=���>}�����N�&o�>&C>e#->��??<+%?�������3d��&,�ox>i#�>6��>$*>ąJ��m�=��>�Ua>�?�怽�I�k@��V>Ӟ}��H`�K�w���y=a՘����=�$�=~V �_<�nR(=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾUz�>>��g����'�u�,z!=X��>\H?3c���1R���>�J�
?��?�����	�ȿ݇v���>���?��?D�m��5��*@����>؏�?�OY?~ai>��۾C�Y���>��@?x�Q?���>�&�6�'�.�?��?u��?��^>ﰛ?˶d?��>��콏;�;T��$ȏ��-
��0�`��>.f�=����:9�p=��������d�N��I%>q;��>�{$�TBx�}Em>o���������=Y�>�	>���=���>J#�>H�>T��>	$>�����a�� {ʾY�K?���?���2n�nV�<)��=�^�X&?1I4?3f[���Ͼs֨>��\?W?�[?d�>���X>��l迿e~�����<��K>W4�>hH�>�!��7HK>D�ԾZ5D��p�> З>N��@?ھ�+��u��fB�>�e!?��>�Ю=�� ?*�#?�j>C)�>WaE��9����E���>^��>�H?0�~?�?�ӹ�JZ3�����桿��[��9N>A�x?�U?�˕>Q���Y����AE��WI�����#��?�sg?�U�A?�1�?ӈ??g�A?I(f>(��#ؾv�����>��!?4��A��M&����~?�P?��>�5����ս&Eּ��������?�(\?�A&?����+a�T�¾�8�<��"���U����;�D��>&�>���D��=�>�װ=�Om�zF6���f<�i�=��>��=�.7��t��0=,?��G�~ۃ���=��r�?xD���>�IL>����^?kl=��{�����x��	U� �? ��?Zk�?b��@�h��$=?�?S	?m"�>�J���}޾6�྿Pw�~x��w�Z�>���>#�l���K���ڙ���F��_�Ž��\��o�>��>���>�k?�vi>��>g��(�*��6Ծk2 �?.x��*%�7�6��7��[�JP����O�*�=.�X��wXw>�>� ^�>�K4?Q:�=��I>�N�>p�=X��>+y�=�y%>3��>4t�>zfd>�7X>kں�1ǽ�KR?G�����'� ������2B?rd?Z2�>�i�J���t����?9��?Hs�?=<v>7h�-+�+n?>�>����p
?�Q:=3[��L�<�U�����2����̫�>�?׽g :�XM�\of�:j
?e/?���4�̾�:׽�Ϟ���=?�?�)?c*��P���p�E Y���S�
���/`�� ��m.#�Цo�@/��-Z��{烿8P(�|�0=3-)?�w�?U^�D�뾡k��x�l�G ?��f>7��>S��>7��>nI>R�
�Z$/��}]�V�'��]��[��>jmz?&��>��5?w�*?]L?��W?���>�o�>��v;�>��k=���>�5�>| 7?u?t�5?ò?�/B?��>`��Z�	�8?ྊ�?�
?l�?�u?'�>�޾/�r���:�;vǽ��G�t�;>d2;>��d��μ����E�<��:>�Y?r����8�a����k>��7?À�>��>����)���3�<��>T�
?�L�>����,yr�[]��\�>#��?t�fy=�)>W��=����uӺTh�=�z����=����r�;��<�r�=N�=�cr�0���t�:TN�;,��< u�>6�?���>�C�>�@��/� �c��f�=�Y>=S>}>�Eپ�}���$��u�g��]y>�w�?�z�?лf=��=��=}���U�����G������<�??J#?)XT?`��?z�=?_j#?ϵ>+�jM���^�������?I�/?^3�>��� Ҿ����l�4��e ?��?&a��ye�u�)��c�\&�8��=~@�������w!���=����a�����?�О?�����,�<�򾛷��(n��o�D?o4�>i��>K��>��9�V~t�s���86>� �>�#`?ɐ�>��h?�n?��h?��t>ӊM�%0��/X��A|��2�>�>? ؆?7q�?j�Y?6��>�M1>���*
�?�(�H����T��`�g<|=T>���>��><=�>��=ld���㊽��ؽDʚ=T/�>��?eU�>��?e�,>�����F?M�>d�c��3Z��Ux�g�9��}t?��?��*?^Ur=�,�nC�d���=�>���?��?m�0?ґV����=��Ҽ��¾�Iy�az�>��>�n�>EL�=ֺ=`�>�^�>��>�$���ԥ7�U��}�
?BF?m��=�ƿI�q���p�Xɗ�9�d<����Re��ؔ��[����=����Q��1Ω�I�[�-���H���S������C�{���>�n�=\��=^��=��<�eɼ�ؽ<��J=���<��=�p��!m<��8��Jϻؠ�������\<�I=1{����˾��}?:I?�+?o�C?f�y>�=>u�3���>�~��A?4V>r�P�����z;�x��������ؾ�t׾��c�\˟�iH>O\I�L�>�83>;�=8�<��=�%s=���=�?Q��#=�'�= S�=Z�=���=��>S>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��7>�(>��R�}�1���\�Ұb�
EZ�Ϧ!?/K;��Q̾��>�9�=6߾ւƾ�y.=�_6>u�a=�V�TQ\���=�@{�ȇ;=�bk=�>��C>W��=�0��O��=�I=�2�=��O>�����F8��e,�b�3=��=w�b>�&>"��>|�?y5?�:]?���>�R�l8���T���g�>VL.>�>�G>e[�>���>�K?�7F?�)a?���>�����k�>D�>	c8���g�=)��U䖾�6a=g��?�m�?���>$�4�t֓���C���+����(�>�3?��9?�>���'��p���:0�L�j��P�=������ll>��w=���ZY��r�=���>j#�>�-�>r:�>f(�>���>�&�>�$>���=
m�=�
�<a�1<�Ȕ���=U���<%���3�=	>�*L��k�<�߼��<,#��UϺ���=0��>� >F�>U�=fƵ���+>������N����=^觾?#E�:\d�N'����1��9>�?.>n�H>��[��ڔ�.�>�P>�e6>�Y�?>}?��
>@b�Zʾ�뜿�,[��+m����=,.*>Ra�8$4�%�W�5K��dԾ��>Rgc>W�>OM>�n���[�[�=$��֫R�2��>@����f������ǖ��ܸ��쟿�p�W���{e?�󥿿p�=�T�? #?� �?QN�>/��+����>���X�K=Wb���`��vQ<�5?�O?���>�0��w[��H̾����޷>wAI� �O�8�0�0����_ͷ����>�����о�$3��g��������B�Mr���>�O?a�?�=b�gW���UO�*���&��Mq?�|g?�>sK?�@?�$��z�ar���{�=^�n?���?=�?�>.r�=�\����>~	?̲�?j�?��r?T@�,��>�ݻ;X�!>�ٚ�;�=�/>uZ�=b��=^�?�F
?R(
?�/����	�79����C\�|�=��=9Y�>2_�>��p>6K�=�^=w��=�~[>���>F
�>j`>X�>_��>׹�z4<��Y+?,�T�|	?�h8?�d>����46�k��>~ý�~���Ҿ��F��%Ž#J�=��F&Ҽ��7k�?̿縖?9,������?*�����=�F>��>{��=��>�>���=r�?'d?1�Y>��>6��u>Ѿ�
>����U!�$D���R�;���>�f��RC.���
�t�콺�M�A���=���j�q7����=�0�<��?�V �Tk��*�\l���?�ب>�L5?����q�{���>
��>�3�>L�������V���p�G�?��?�;c>��>G�W?�?ƒ1�'3�vZ�+�u�l(A�'e�Q�`��፿�����
����*�_?�x?/yA?S�<*:z>M��?��%�dӏ��)�>�/�$';�@<=s+�>*��-�`���Ӿ��þ�7��HF>��o?;%�?vY??TV�}%I�� '>�(9?J�0?͏q?��3?�09?ZG��#?�k:>�v?�_
?�7?].?��?�=@>;�>��|��� =�ϕ�-H����ܽFxڽ�f�� =��=L��;6D�<��=cPf<����.S��A;4{�Ļ�<��<=��=TM�=^�>�q]?���>͚�>cT7?���7�'x��a"/?��A=�W��󱊾̢�5��z>)�j?��?g[?+�b>�>A�9�B�pO>�$�>�(>,`>v]�>x��dF����=?>�>��=&1\�rP�����f����{�<�">��>V0|>
���'>�|���0z�`�d>A�Q��̺���S���G���1���v��Y�>=�K?��?�=S_��,��uIf�:0)?�]<?�NM?��?��=��۾��9���J�y>���>X�<�������#����:��?�:��s>2��!Q���x>o��	��p��tL�ܾۧ�=ى�7ܼz��[.�r����w�=u7>�ݾ�R�d)���J���BS?�^�=⬾\���/)��Qc>�ˠ>d�>ځν�� �v@�2���^;�=l��>�>����,�>�� �OK�>_\?׿Q?�މ?�H��My����r��h쾇띾��k�>E?,��>+�>��<V�<�㙾0���r�\4�p��>���>�-�:qf�<���\Sž��.��>��	?��M���?:lS?3^�>�X?
pJ?v�4?Z�>��n�����2&?f��?}��=��ҽiMU�29��9F�]��>�)?��A����>V?�?;�&?�wQ?�
??>�g �|@�8+�>�L�>��W�p���f`>�HJ?̢�>�EY?�˃?�=>��4�����X.���t�=R>)3?�P#?��?�o�>���>@律��=؛>�]�?�d�?�b?Q�3�v�?>�>�o
?e�-�Ʋ?��?{Q?�}w?��x?�9?d�?���<2Ѻ���ğ��毌�<1<pw�=$�=�⁾��:����`��a��:�)˻���ů�& 8��~���"i�P�>k�s>?��e�0>U�ľa@��M�@>���De������0�:�e��=ߟ�>��?�w�>��#��T�=��>�N�>��*'(?s�?�?��3;�}b���ھ��K�8�>��A?�>�=b�l��~��|�u��vh=2�m?��^?e�W�F���b?6^?�s� <��Bľ��d�]��jvO?�u
?��G�8�>^
?��q?$��>��f�^n�����Yb�Q{j��&�=䭜>����:e����>�R7?i�>9�c>2�=q�ܾ�-w�t����q?��?��??�?&G*>�n��F��������Ue?.��>�����,?�$ѻ�eѾŘ���#��tݾ�����ư��˞�s���X��gy��G�AA�=b�?�Ks?>�n?�d?��
��5c���`��˂��{F�����;����=�خ>���U�_=r�R��������:�=7|�v�Y��>�?k�?�C#���?Ѡ�����vԾ�O>Y����t��M=������=�_=)JX���bV���"?E�>���>��A?4b��=�Xr6��]@���޾x�">���>�6�>N��>�;��7T�;��'Ӿ�Z�W���x�{>o�d?��H?�m?#��-23�T8����!��,�1���^V>��.>jn�>��Y����4���:�.5u�q��z����
�R�=Wk-?ˠ�>�ß>}�?/  ?����ߩ�dp�(�.����<c��>�ni?b`�>���>�R���� ���>��l?&�>N/�>�⌾v�!��|��'νM�>��>��>��p>6+��p\����3}���9���=��h?�\��%�_�|�>üQ?,��:e�1<陡><_o�h~!���]'��a	>�?A��=%y<>˖ž����{����9O)?�=?�풾��*��`~>&"?���>z3�>@0�?m�>�jþ;5\�ɭ?��^? 3J?�SA?�?�>b�=_���$-Ƚ0�&��~,=㈇>T�Z>lm=���=���;�\�*��l E=p��=e�μfX��<	����H<��<�4>G��ВK�|�쾡���5��j]��Ӏ���;�XO�#X�������þ�a�Y�0�ZZ�<Բ��f�#���>wH��m�?���?;���;4m�i𤿀-��̓��Ƀ�>�3�Le�-�=�����ɾ�g�#
�HQ��Sa��R��"<��,H:?��j��ʿ`١������>�<D?���?�\�"�A�1W���*>��~j">j �)ʔ�l�ο����=UR?K��>�ؾ��W��y�>���=�q>��o>.���\3���\>�?�f9?���>^�������>��(;$�hG�?V3@}A?��(�T��pV=W��>��	?&�?>T1�jI�����U�>�<�?���?�yM=�W���	��e?-n<��F���ݻT�=J;�=mC=a��T�J>�U�>����SA��>ܽ��4>.څ>]|"�x����^����<2�]>��ս�;��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=�O�,dȿR�"�p�զ�=��=%�>��&Ƚű�RR����>�w��M����R=�4�=��d>�˄>rmj>F�>��b?�Os?�Y�>]�J>/]��槾�LԾ�qK=�Ra�2�h�tO��5�?�VѠ�Uj��X4¾u#%���1�_:*��f��zR����=�hZ�B`��J�)�?
f���8��/>?�B�>�)�('S����Ȯ���幾Ԩ�=9U���Ӿ;@�]��"�?'�M?/P=b��1'��KϽ�'ҽ��B?�����j�׾O��=��T+=!�>r=�Jƾ:�>�6pm��.?�?�Ȿ;��81>�ƽ�2�=I4,?.n?4��<��>>!?	�;��
�R�c>�r0>�Q�>��>�>�ص��f����?�S?���ل�$��>��Ⱦ�ލ��=$�=�j;�.T�<%T>���;Tӕ�Ӯf��&��S<=��V?��>we)��z��
�����C=[�x?��?S�>�Ok?�B?@�<7���S��
�#�=��X?k�h?6�>�x��[ϾXW��6?F�e?W�O>�|i����>�.�n��#(?_�n?
%?#⣼��}�B1���4�E6?��v?s^�ts�����D�V�i=�>�[�>���>��9��k�>�>?�#��G������uY4�#Þ?��@���?�;<0 �>��=�;?n\�>�O��>ƾ�z������ۓq=�"�>���|ev����R,�a�8?٠�?���>������|�>�j��?���?��ﾃ�S=����녿I���{o>yG�=�T��wH�=��E���L��/��.��$@�iM6>��n>KL@+;!���G? ln��V�a˿�v���L���k=�d6?��>]��=�ľN*��;bc�)�M�<�j��M�H�>��>z�����t�{��r;�p�����>3��#��>P�S�'��ԥ����7<D��>��>���>�`�������ƙ?xe��<ο����e��޴X?�i�?�n�?�q?�K8<w��}{�����4G?|s?�Z?]�%��']��w7��(k?N��ǅ`�Y5���F�9�K>��3?`��>�-�tE�=��	>��>>�3,���Ŀ'���!� ���?���?j�^!�>�@�?�+?��������>����,���qD?$7>�0���3�T8>�}�����	?�h0?<`��k�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�&�>��?�w�=�c�>~��=������/�zX#>]!�=�?���?��M?]C�>�8�=;�8��/��WF�uKR��&��C�k�>��a?)yL?�ab>����1�{!�jͽ�^1�����J@��q,�0�߽�65>��=>�.>��D��Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>D�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*/bֿo:X������/�=�s�=��2>f�ٽ�-�=�7=�:��0�����=h�>
�d>-�p>BO>�\;>[�)>����!�;m������!�C����f���Z�O��.Uv�&j��7�������᷽X�½�У��P��-&��`�!�=W�O?��R?��k?<,?l�=�]�<�e��׃�q�u�5>�O�>k�/?�w7?�4?\/
>�l��V��<���7��ܑ��5�>�UY>vە>{��>�>]w�:�.T>�;3>�0>��<��=���=ü;=.�>��>�2�>g'�>g4�=�w>�����e�� )P���ܾu��=���?��˾��w�ʐ��y_Ⱦ����.�>Ų�>�fX�n���"���0簿�4l?�&�����ɐe�d�R>�?D�j?P"1>��\��>��u/нsL�=����c �>Z'����ü�-��q�>��.?�Qu>��r>gV7�yT:�HHO��������>��8?x��i�R���x�}LF���߾,�a>�+�>�y���i!�V/��F:{�ȩb��#m=��6? �?�(ƽ�Z���$k�`���a1Q>��^>]�(=u��=�M@>�2u���ϽM-H�Z��<`�=�>t>�?��.>b+�=m+�>gK��MA,�-ǲ>��R>��<>�\<?�i#?����m���3������m>�o�>��>��>pa����=���>4�r>,��;)�������^�E*>�����]�w���!��=����P�=�p=���;O��0\=�~?���*䈿��.e���lD?[+?� �=a�F<��"�G ���H��=�?q�@
m�?��	��V�:�?�@�?��:��=}�>׫>�ξ��L��?��Ž1Ǣ���	�)#�hS�?��?��/�Wʋ�8l�b6>�^%?�Ӿ�h�> x��Z�������u�"�#="��>9H?NV��H�O�	>��v
?a?�]�ϩ����ȿg|v����>/�?q��?,�m�SA���@�ʁ�>��?[gY?�ni>h۾�^Z�ڋ�>�@?�R?��>�9���'�J�?�޶?گ�?�Z>���?��x?��	?����
:�����r���ww�V >�o�>�4>�^����Z�G��c��nuf�T���M�>QN=
��>�e6�_�����=�����ƾV=0��>yZ�=.L>��>C��>HW�>R�>���#d��{��\�����K?ײ�?��&n��-�<5S�=^�^�~?�B4?\ \�ɩϾL�>��\?���?[[?�l�>����>���翿������<G�K>L-�>�;�>�ሽ�kK>��Ծ/2D��t�>�ė>۾���:ھr���B��Z7�>�g!?7��>���=��?��&?Z>gG�>�yE�υ���N��-�>�4�>�G? z?��?����Sn:�T�M��9�Y�U�,>��z?��?���>�s��-+��C/O�%Q����.k�?�Nb?�\�zJ?~�?.s*?�fI?��>�n��ƓϾ0"���]!>v!$?G6�,�E���(�f��?��
?�>�<e�����3`�f�p����?�U?�o ?�T	� l^�O���Zj�<�E���R�6<�r¼� %>ݢ> ��Py�=��>�H�=�CZ���A�eB�;3�=s�>�Ѫ=��,��<)��2,?��?�ᘃ��O�=�r��<D���>C�L>�A���^?��<��{�o���o���eT���?0��?��?�O��$�h���<?E�??�u�>���u޾=��.(x�]x�Տ�aH>c,�>�aj�����Ֆ�����JŽ/��@ն>�6�>C��>< ?�D�>z�>��t���!�8�վ�w��p`�~E𾯤��8��5��� ���=7��en���S->p���
b�>ό?j٠>\ě>Qq�>^uu�7��>���=��I>Y�>��>���>��n>�!��G����fR?�����
(��#龸�����A?W�d?���>)�d�Q����%��H?L=�?�}�?<u>�rh��d+��6?���>��/?
?O,9=K���4�<5������Ƈ�;�a>�"ֽ`�9�lM�a�f��%
?��?y+��S̾.Bӽ�Ɵ��Ls=l�?��)?�*���Q�]�o�mX�P
S�� �df�;נ�1�#�+}q�;���(����w(�;=*?�9�?���������k�!g?��Cg>E��>*ޕ>㚿>�L>e	���0���]�Ҧ'��d����>��z?�\�>�`:?�C?��T?z�@?�.�>h8N>�����>��=y��>���>[�?2C?��E?�0?Ί"?�5P>�z����İ��4$?�j?�?�	$?��?ُ��W .����=ݿݽ7��� q=�m=�p=�h���0������=���>nk?ն��q:��J��p�d>!T5?թ�>���>}Z���3���Յ<���>�?�-�>Yh �3Fr�Z$�n9�>:�?�c� ='1(>5��=�~��c;�3�= �ϼ\U�=�m*�c+��u�<�W�=C��=k�$+"��j;�u�;���<�t�>��?�>cF�>6��� ������=�xY>�$S>QA>>+پ���Q!����g��zy>�~�?���?�g=���=���=�e���#������������<��?�#?�@T?|�?l�=?�s#?��> &��R���b��fᢾ~�?�S??A�u>3\'����Z����1��g1?��?7_N��~���G�c3�滼=?y>��Q�*�������~0>���c��k�?^C�?<Ti���"�k~.�=ؘ��L���t?�n�>1�>�Z4?��9��8\�z^��oA�>��>�.?���>jb?�J^?6�N?@Ũ>�zD�UG���y��^��Y�=k�R?W��?��v?�TC?��>ڒ�>��
���P_���ؽy�i��d��{�ǣb>u�>���>�v_>�>�=��y���ҟ��M�=��>!?	�>a�?��>uHt�Y�;?hQ?X�����P�ξ����t#��S?�&�?��(?K�W>���a��4����>�O�?L��?]fH?�� ��Y�=k�U�jR��o����:�>'��>���>X>�@�<\��=�c>G��>,!9��%�9�*��ֽH�?��M?��>�ſYqq��Zr��0��ʀ<쐾Gb�m�����[�@��=����:�pl���EZ�����"u���Y��x�]y���>f%}=���=��=��<�������<U�O=�)�<��=�jm��;v<��3�P�c�������#;^w<�D=K9ʾ� }?UJ?Y,?��D?��}>2>�'i����>��p�K~?��Q>�~4��%��#�4��2������M�׾-�ؾ��g������>�ND��>X12>x!�=_��<�@�=�kb=e=�;PD=K��=���=�=*�=��>�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�J8>�>��R�Y�1�)�\���b��HY�s�!?;���̾���>/��=�E߾x�ž��,=�5>��^=�z��,\��=�b{�<;=Pl=l��>�BD>� �=Tt��׶=��J=�&�=�8P>{��J\8�H�,�R3=�z�=c�b>�'>.l�>�&?�/?/%j?��F>"�S�h�ؾx.�����>U�>� ?`�V=�kP>yB�>,|A?7�E?�j?ﻴ>e�&��>^��>oXD��(p���ȁݾ��<Iʛ?��?�д>��Z>���wL���/���f��1?�\?H�#?��>hT���TY&��.�Bn����8kH+=�`r�
vU������s�)��D!�=p�>���>��>�Oy>��9>6�N>��>�>���<�c�=3Y��V��<S������=������<�bż+q���H$��+�Lڥ�K�;��;l]<���;���=�%�>Ix>�o�>�З=p����<.>پ���7M���=ё����@� �`��x|�J�/��;��L=>��V>p)x����^?$�Q>Q>>��?o`v?�&!>�����Ѿ"n����[��c�ų�=�
>��6��h9�=4\�9CM�~`Ѿ�d�>�?>d>�>/h�=�7 �^�&���P=�:��E��h	?ޑ�����=�4�=�WQ�Vo��[�����h���3=�]<?T���L<=��g?�S8?�X�?�?��/��~Ծ*�>����HS>�jE�Rj���Ҥ��r?��?��?���9�3��H̾W���޷>�@I�-�O���R�0����3ͷ�3��>������оh$3��g�������B��Lr�Y��>%�O?��?c:b��W��HUO����;(���q?�|g?2�>�J?�@?;&��z�r���v�=�n?˳�?P=�?w>��=u������>�C?��?���?��r?́>�zk�>��;<�>������=��>���=��=5?�D
?��
?�g��]3
�X����𾶹\����<�6�=3��>mĈ>�s>���=�uh=���=1_>П>�{�>D�e>	d�>��>�y�
�I��?,ш��į>+R?p%�>*K�=qGT��c>���;�~�l�����l=��E���=8uH<�,L=.�;=K��>�hɿiP�?t�5>��j�?�(�����q>�"n>��&���>���=3��=���>�$�>,�>S�>��=r�Ҿ!�>A�հ!�#C��xR��о4~{>*����(����Q��LK�$q���B��%j��+���==��߳<4�?������k���)�Y5���?�ĩ>ż5?�N��-ه�`p>)s�>�~�>�F������Ί��F��P�?��?�;c>��>I�W?�?ؒ1�23�vZ�,�u�l(A�,e�T�`��፿�����
�|��.�_?�x?1yA?�R�<,:z>Q��?��%�\ӏ��)�>�/�&';�@<=x+�>*��*�`���Ӿ��þ�7��HF>��o?<%�?wY?=TV���a��U">]�:?x�0?�aw?5~4?ܑ8?p��W}!?0:>�?�l?|�7?f-?t7	?hWC>��=Hͻ.�!=ҫ��@щ��iҽc|����#�C%=.�=k�v:p�;=q�<O��<v��{r��r<!���iv�<_�a=�q�=^2�=�1�>�lU?D�>��>M$?̤۽z��QnG�:D?�=�(��"q���׾@p��-2>ޢc?�-�?�<�?��m>�FX��z�->��>�Y�>��>&�>n5��� '=E�;q�T>a�6>G弹߈�X�&�f�Ⱦ�[�=��;>���>�0|>����'>{��Y.z�ˢd>��Q��̺��S��G���1�Ӆv�=Y�>��K?��?���=>^龄4���If��/)?^<?KNM?��?�=��۾��9���J��;��>8!�<t�������#����:�͇�:��s>0���i��:sd>h�~�ྋo�/�I�����x=@k��0=����־7������=b1
>�Y¾׿"��������"<J?E�|=ӥ��
T�&���>$�>Q6�>��-��x���?�]���p��=��>�5<>| ��! ﾐ�F�1���l�>�f=?�l_?I~�?����|V�n!=�$����)�����?*�u>���>]�i>;X/>1Й�����Z��Fq����>�d�>�e��]7����O
����B�>0�)?�=M�>}�0?���>��R?^_%?�~#?���>���$�����*?t}?{�:>�N��`�~��2�9�:�Cu	?��a?Ŝ@��|b>�j->(��>��+?'�l?��?��>@�*����q��>��>TQ�D���W�.>0	?���>Cr�?�S�?c�x>X��n괾�ݽs	[=�kQ>w�9?�u2?>M?��>�T�>�}�1�?��}�>ȕ?���?J=l?.>mY?B->YW�>�h���T?n�?'d4?g��?��{?�X? ��>Ԛ=����$e��"Y��PP�u� <���<�n�<a��<w�������%�@�`��&Z=F�=�m�<��1=}����@���k�>��s>?���}0>h�ľ�D���A>������������l:�%|�=0`�>��?9Z�>Wi#��P�=�ټ>B�>����!(?��?�?��%;�b��"۾��K��3�>SB?���=1�l�Bz��)�u�&�h=n?gw^?L�W����E�b?.�^?\1��;�.�þ9�e�f��#BO?�s
?�SC��'�>��?��q?�>��d�;n��!��A&b�W&f�Hĵ=e��>����Zd����>FU7?��>�Ab>C4�=�ܾ��w�����@t?T�?��?��?7)>��n��1�ȝ޾Ĳ��VQh?�ۭ>'ղ��D&?UO�{�Ѿ�Ny�ԙt�p�ԾG:���]���-���~���7"�Bn�8��Î�=��?��y?�}?&m?��Kd�\d�a}��g�/���۾�6�C�G�L���[�wst������6��^�!=��g�
G���?Xn?p<����>`K��H(���ƾB!H>�̙�*]�.2�=[��M=��Y=�P�5`�H?��+s?���>)"�>��??�`a�"2>��5���8�+�о��S>�П>N��>�g�>�8��$-H�i�wM�8�z��Y뽩��>�z?j?]?s/�?��&��i.����._#�`��sW����>���=�!>Zg�䷅<T@���S��	�����vꆾ�)����<�`?"T>U�?�ܫ?�)�>z�徲�)K�>l�p ����>!b?�ʧ>�߾>4f�� �����>W�m?R��>Z�>Ϧ���"���}�yԽ���>_6�>k?1�w>\�.�H�[�����\���":��_�=lhi?u���J�\�t�>
Q?�;B�<�I�>MFt��"��򾜾#��=>��?�z�=��@>�ž�6�q�{��ċ��Y)?QB?�e���A(��v|>'.?��>q�>�D�?l#�>������?�@^?�K?�A?���>2Up=<��:н�0�ʌ-=�ԓ>��i>O�=@
�=s1��7t�n��wcO=���=�h��,֫��25�Nk��.Ȼ$� =�\G>g�׿�M�n�_���`ɾ�z��b�/�=�J���Xe�^�ؾ�����M���.��o�ar�/i���搾x�+�@%�?Bt�?�H���Aݾ^���v\u��ož�`?d���ࣉ�a� �k�'�>�������[���LJ��u�+�e�_;t�/U$?�+���|ſ������IW?l�?Z w?�)��%�j�9�Fw&>[�f�cO#�e�辏�$�Ϳћ���W?5��>{�ﾊ:���I�>|̅>K>4�v>��}�Ao���,<�K?��0?�a�>Z儾� Ϳ�o����=�(�?0Q@X�??5/�i�־�ѹ$��>S?�->L�/�1>��l����>Eٟ?w��?\�c=S�Hؼ�re?S�j=#�<��N;�p�=�z>�� =��7�[�5>!8�>��&���������;>qр>
"L�$@>�'Pj���<��3>�n��T½5Մ?,{\��f���/��T��U>��T? +�>V:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?8ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=x6����z���&V����=[��>c�>Â,������O��I��X��=�8���ǿY�.��T�r�=Ħ��z�Z�����!���Wf���J��a)�����G�|=���=7Q�>�Jr>eC>�p�>�pY?ijo?+�>L�R=+ɽ���+��jL�=b���B���	�Ǿ�v���蓾�A/�������%�������X<�@�=[�Y��S��i�'��Z�HB"�)�X?n�N=���<q���H=Q�~�\����+��r���1�b^����?�d?����a�ZB����@kI=Pjo?�O�b��q2��5�=B܄�a��=iQk>#�:���$���0���M�
�0?��?����Î��>4/�/�=؏7?�$?U�;=1�>�I?dw0���j�<��>�^I>%�>���>��>����q�@w?�-b?�=5�A�`�e7�>h#�#
��
>1H>�F����<��E>��p눾a���.ν x=�%W?T��>A�)��	��h�����.>=��x?-�?P%�>$ik?��B?���<0e��v�S����x=*�W?i?��>�ā���Ͼ�k��5�5?��e?n�N>�h�����.��H�l#?��n?�i?����io}�������Wn6?��x?��)�bm��2i��I��=� ?1��>�V�/Q>��-?у���P����ƿ�`�mC}?���?X��?�6=�2��X�=�+?���>ë���TϾ��4�>Z���a�=�?9g����g��*�ـ��|&%?H�?'��>q����mH0>'�n��ֺ?F)t?�"���>=�n9���y�)Zx�C�S>�x�=e�<zҽp-���P���վ�#'��㶽}<>5P2>g�@�H��O4?���\@�Y6��s��M��F�w=�r@?�P�>����!���Y-~��Et���d�(�f�r���N�>��>������*�{��n;�W6����>�����>��S�~(�������5<�>���>	��>BF��=�xÙ?�_��x>ο������k�X?f�?�n�?r?o�8<D�v�ۑ{��M�}-G?C�s?[Z?�T%�9]��7�&�k?������`�uu4��[?���>G�4?Ct�>�!7���\<�>?��>���=��;�7Aƿ⍱��jھ�ܧ?)X�?���f�>d�?�)?���@K��D�����%�X�;�F?$�>I:����"�H@<�Q'��YK?F�+?�����]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>gH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�$�> �?Y|�=�c�>�`�=��X�-�5i#>�$�=��>���?Y�M?fK�>�Y�=��8�/�m[F��GR�""���C��>��a?�L?�Ob>����2��!�_qͽ�h1����o^@���,�ْ߽�,5>��=>>g�D�$Ӿ�%?�$��%׿�?��F�-��?�8�>�r�>�}+��>Ѿ��=w{{?,i">�,��L��O}���(��:�?�s�?�
?K+��$�=���=���>��>�fw�_Z�I�c�b�>l5?T�`����W���>,{�?|��?��?m6T��K	?���f��j�~��M���8�B��=Hp7?O��+w>��>vŰ=�|v��Ǫ�VQt��A�>!!�?�l�?p��>Mhl?f�n��B�5=�y�>�Pk?G
?�f��]��zZE>�p?x+�X��:�)�e?b�
@0C@�a^?ݢ��a߿�j���긾��ܾ�E>���=�>tq��p�=�ҫ=!/�������G>��>��m>q>{�}>H�{>�t>����#�/K���ˈ�`�,�F�
�2 ,�B����[�b�#��9ߑ������6t��4��s�[�}��0Kݼ��»(�>��N?��X?�
p?�Q�>��7=���=����=R�ѽ�u|=��=�}?ĎN?��3?�ϩ�T���7���i������˻�����>�j#>���>���>���>��1=N�>�n>a��=ß>خ=���"�"=� �>��>���>��>E�>��=>�=��B��8�r��E�� ��W��?���Bc����2{���6Ⱦ�̓=ȍ!?J=)����ʿ!L��r�I?�OK�*�����	�q=�?,Z?�>�X���g0�t�>�G���A�=C>�j��������*���3>��
?�.>��>�_G��O�"�i��`�bַ>�T`?�iɾ�AӾ�����I�'l��*�>�?�>�UT��C]�	�� s�i�(���<G�9?��(?�����p ��(�
�B��>B��>��*>?��=�Ć=M%�Mߡ��[��.>�e>.��=��?:0.>��=N|�>����S���>�nB>�'>��>?+�#?������Ʌ���1�Qw>U]�>���> >[OL���=T��>i�f>���r�rg�v�E���Q>xqP�;%a�j�q�{��=An�����=� �=���s0C� �=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�e�>���Vu��uTz�o�t��"�&�?e[?���O٩��c��.?�8r>C�%�����sӿ.O�u�>��?B�?uyJ��e���XQ�8#?���?QC�?2N>�/������'�>7�P?��e?�>z�^��i��;;?��?A�?0)�>.�?��?o#%?'U��?�H�Rȿ)Z��2�c<�`�>UN?���>�z;��P�
뎿;��N�\x��P�?�L=���>]���K���)�>D�p�4��R>�o>9�>�F�>��>͓?,!?N�?�h��Q�����W�`�|�K?ﲏ?v���.n�0�<#��=6�^��&?8L4?5B[���Ͼ�ƨ>��\?���?�[?uc�>A��J>��H鿿�z���u�<~�K>�+�>�D�> &��
MK>��Ծ	D��p�>�̗>��9ھV-��q��%H�>/g!?���>�=��?+Z(?��>�>��G�b����O�p��>?��> �?zR�??o���(x4�P��^!��-^���B>�P}?^?Z�> ���癿&hv<>��g,ν�{�?c�_?���̚?��?��D?�H?�Q�>��aӾ:Dǽ�>+�!?��	�A��F&����E�?MN?(��>r��p�ս��ּ@���q����?�'\???&?t���,a��þ�Q�<�t#���W��.�;�D�*�>ڃ>n��Xմ=�>���=�Rm�G6�j�f<3��=`��>+
�=�-7��u��*�2?�ʐ=jhB���:��v��;`��Ϥ>B�&>�\
�JD9?�k���E��1��z����hؾiu?tн?ъ�?� ����\��c$?9�?l�>�`�>|Hm���پ,��-9r� ���ם�~*}=�0�>0�=���$��uP���i�*����`�.S�>��>�?�T?��h>���>r����*������U�%��hB2�k`.����Ґ��6���Ҽ�tǾE��/g�>��#�N�>T?��X>'��>-��>��׼���>OgZ>m�>:�>�ey>��\>�h�=�|��`�˽�8R?	���[�'�\���u��OEB?�ad?���>�k�D��������?8��?h�?��u>�hh��+��j?03�>k7�� M
?��7=�2���<�������������o�>�׽7 :���L��%f�!�
?xY?�C��޶̾�#׽MX��د�=4Z�?^z)?b�+�PqQ�r�o�s�W��JP�p'��>c�8���&��r��ꏿ�b���f���2'���:=��)?5��?����q龌S��C�k���=�_kd>b��>OB�>�g�>'O> t
��(1��[_��(��}�i��>��z?%Y�>�(?k0?vfc?�bX?@��>���>�C����?��>_y�>dF�>q??��:?��*?�?�%$?!�=Cp��d�6yľt�?��+?��I?��?��> ���6��%/�qSp�J�1��n&>��/>��$�h���r��D��K挼N?���p�8�ѿ��&3k>d�7?0v�>t��>,���3�����<��>2�
?e8�>H����`r�S�lL�>~��?"G��=H�)>i2�=艅���׺V��=��,�=_F��j�;��$<Gg�=�Д=�d�L�E89��:'9�;�H�<���>�?�r�>���>Wㆾ�$���o��=��U>�R>m>k@ؾ����#c��-Zh��x>�w�?Ot�?�Rf=���=�[�=�9��Fu��T�<����<�?��"?��T?4�?�]=?�`#?�>
�����xH��⢾ys?��?Xo�>j��Jl̾���v8��v?x�?�U���}�e;�W����T�T�=���I������E��1ν��'���A�?�	�?��+���$�@���j�����K�A?%�>�n�>'�>7�:�"ke��`�~�>A`�>N�>?���>��X?I|?@+]?Q�;>I>�5��K��$�л��[>��T?9<�?�#�?�sn?��>ʺ�=g]`��<�Ѿ"�$��`齿w���7=e�v>�G�>�>��>��=�������jm��-�=��>�O�>^��>6��>�8>�LR�DqH?M�>,���>!�Ů������ZC��Z�?L��?��?��,=�A1��F9�|�����>H�?���?�6%?	&���G�=���3�ھ�:�h�>���>2]�>�=;����T>��>�k?��̽Bs��V;��� ��_?��o?���>ƿ��q�u�q����~�c<����je�$*��"[�'�=ݾ������1���~[�
���?��ﻵ��e���{�5��>�:�=q�=2��=�&�<q�ɼP�<?!M=��<ߡ=F p�g<sz:��̻d̈��_��]<2�J=�ۻ�R˾�9}?��H?�a+?h�C?Y�z>�0>�6����>�����?�V>ΏM��Q��Sp;��"���ڔ�PyؾS׾C�c����t�>iI�Y> �2>���=�a�<^�=\	s=�,�=W5h���=���=f�=3ì=/�=>.�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>X8>N>:�R�h�1�I�\���b��	Z��}!?l];�Ry̾7(�>�3�=$v߾o�ƾ �*=D>6>$9d=���H0\��=�z�ӝ>=��m=7��>��C>�˹=�د���=�rK=2:�=�yO>����\9�Ϧ+��6=�M�=C|b>��%>�C�>��?U�0?��d?��>i/l��Ͼ����ג>*�=�;�>�W=�m>>���>B�8?k�C? �I?�B�>Ͳ&=��>�N�>�s+���m�k�從G����<q�?#h�?�5�>�s5<�J��r���;�ȴ�"�?��0?��?�}�>��B����c�2��_h���/��͗�=蟾��ڼԙ5>�m��;���>&ٷ>�)�>A�?��q>&�>LQ�>�=�>��N>����`>�:!� ����1�=$�D>��!U�������=���g潙�u�=ۺ�=���>2�)>���>�8^>4cE>/�X<ۮ��4VT>7�̾}g�/��=�|����.��kZ�F�y���F��w��aj>aR�>���������n�>H��=�>���?��?�n�=�d~�7(���ߎ��N"��&����>�|�>�7�<�-��V�2�K�H,���,�>rf�>��>�q0>��$�F2���=�q����>�}4�>�����w���
�L�i��������[�z=Q.@?ؚ��S��=S�g?�G?�'�?�{?7?��Zlھ�D>�+���OR=�m�<L����<�'?Ŗ'?�n�>Z����[<��˾Eٽ��۶>�H�o?P�����X/0��9��෾�ݯ>m'���Ͼ�3�����CꏿrC�W�r�)��>�9O?nڮ?��a�|q��jMO��'�P����?ݙg?Y�>��?T�?Os���_�I����=*n?'��?J�?�i>���=�p���y�>��>l�?�-�?'cc?�e�����>���,�=�v�lM.>ge>�wE= >`B?�?��?������m������a��Rم=�K�<rK�>u�>�S4>1��=@�I=b��=��H>N��>O�>�b9>��r>lS�>��h�#n�&^?�ؕ�}�>L�G?ܴ>nT�;�?g�����U�ؽ��ؼS-U<��Z�#�5x=[��=��K>J�>nP�>q�ÿ�d�?l3�;�+�;�>�����<�M�>hF�>DM��o�>֛_>f?A>��>'%B>M�L>�)�>�.>B�Ⱦ��>%��Hd��iM��pT�����@�>	ə���m�"�����U*���7оh��G]v�����{7�2De�o��?��
�qki�z,!��E���5�>���>�8?���Žv�l>"�?Xb�>�Y�[o��A~��"���y�?��?<c>��>@�W?5�?�1��3��uZ���u��'A�e�3�`��፿������
�����_?��x?�xA?xB�<f:z><��?��%��ӏ�x)�> /�';��D<=�+�>$*��(�`�ȯӾ��þ�7�aIF>��o?)%�?ZY?TV�\&s=$k�=�`?��5?�K�?��g?�.?8N���4?�N/>�r�>1d�=��2?�&?� ?-p>���=��.�&�=s���E���tf���%g��9���<F�< ì=�����*=W�p=�F=�E����
�7���=�@=��>��}>	r�>�Y]?i��>�C�>|�6?*��O7��=����/??=�7��������ﾞ >��j?�ݫ?ʚZ?��c>�nB�x�D���>fi�>�?)>2�^>?y�>���NJ�&��=��>l�>*4�=�aJ��ɂ�k�	�q���R�<3i">���>e=|>�ލ�D�'>rh���z���d>V�Q�%���^�S�B�G�^�1��tv��\�>��K?k�?M��=r3�:��h9f��)?0^<?:eM?��?۹�=��۾�:�&�J�����>vc�<���T������S�:�U�:�s>=���3����c>��I��ldo���I���ʢd=���<=���}Uվ-���y��=��	>����v\!����;T��J?��}=E=����Q�,P��R�>ꆙ>T=�>��;�Ziw��@��C����=�a�>��6>J̼ش�
�H��=�s�>T�K?F�b?�-�?ݷ����l���N�w��'���]�;~�&?1ݷ>H��>(*,>ݸ4=j��)���nk�%z<��H�>���>��!���J��yj����G�*��]�>_?�/�=rl?8�G?��??Xc?�6?W��>M��>�q���þE&?6��?��=h�ǽ��J�QO7��jF�g�>�f,?i@=��>�\?[�?`�&?nR?�?��>�� �#�A� Ŕ>b��>�|W��G���A_> eG?a��>�[?ܼ�?x�:>��3�r���>H��.��=��!>9Y3?��%?�;?�>1��> �����=V��>�9c?��?�o?��=� ?K3>��>��=|r�>�>�>�c?�XO?;�s?K?o�>D��<A���񮶽��m���?��ܘ;|/Q<6�s=�d�M	q����օ�<ǻ�;���������$�J�����<�_�>��s>����0>�ľ�7��D�@>����J��e�����:���=���>��?���>�M#�옒=G��>:J�>*��\9(?\�?#?w�;V�b��۾B�K���>CB?���=��l�䅔��u���g=8�m?ׇ^?��W�u��%�b?��_?�����9�����lh��Q�z%M?�?tH��+�>4?}?Up?��>�b�Al�H��]�d��so��^�=��>�,��xc��W�>�|5?���>�jf>l�=�\ܾL0y�+r��,�?:�?RP�?�R�?�^&>�cm��>࿅��H��*�_?O��>��P�'?��ջʙξ�ㇾ0ē�������@x�������ӡ����u��$W�����=��?eYt?*�p?�mf?�� ��Of���_�!����P��e��E���rC��VI�f&E�V�m��2����	��9Z=��O���T�ֈ�?�?(M���?���B�پk<���ƺ=m����⽓�}>�{��D�=s�=�;{�O���헾�R?��>�*�>��]?@^P��FE�o�7�$N��n���Om>'>�>�+�>���>�-���d��=3��ʼ�By�� 赽�̎>�m?��D?�
j?�9�4�3�5싿���N�N=½��WG>��>���>?���i���b�:��S��S.��
��`�n�<=A(?�Ix>钙>ފ�?i��>���;���k숾�B-�qK�=�>�>�yj?���>3{>�׽�19����>Y�l?��>��>�U���I!�E�{�˽���>��>��>cuo>P-��,\�f��4~���9�No�=c�h?鏄�; a�ƺ�>�R?�[�:
R<�}�>f�u���!��ء'���>�?�Z�=�;>Hgž��e�{�n-���B)?��?�x����)�>�>�G!?�`�>oc�>���?ᴜ>H\��%Z����?�y]?&=K?mB?���>ʊ,=;�����ƽ��&���4=�4�>9�[>��u=���=�k�śb��S���H=n��=�ॼNj���p<j޼��;<�K==�:>��ɿ��7�)��#�Z�߾��YS��<�<{��� 'm�?oþY��+���]��r;HcX���V���A��l�p�?	��?��Ⱦ U��3������X����>Ӆ���+�x�ﾬ�+�#c������ʾ��H�V�����{� b��g0?�Fu�в˿*۞�Z�ľ�q�>LV<?7�?�8��D��7]�㹺>,K=s���܊��	����˿�u�<�l?J��>*&龔s�^�>�׀>��Y>��>Xؾ��վ?O���� ?- ?���>y�@��ĿMj�����[�?@�A?6[*���J
N=�(�>�?�:@>{�-����\��~��><��?4.�?g�K=�_V��I���c?n1�<W�E�
h��g;�=�V�=5=���w�G>�!�>G6#��h:��(ֽ��4>�i�>��4�a=�C0X�w�<��[>��ϽXߗ�5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�򉤻{���&V�}��=[��>c�>,������O��I��U��=���F���o� �.��=R[@=e�c�ğ��q����X�e5���6��������>��>�^>�֙>j��>�FR>�*Y?��m?d��>�O�=/���6���L��8�T=�����R�{���� *�ᅥ�Ֆ�Wܾw>��P,���z�پG�4����=}�W���U3,�``^���3��G7?���=n�
S���	;Nݾ���k�%����پ98.��g�6�?��G?�����F�&��q�\�G�{-O?Yl��t �z����'*>��W\;8/�>�̙;�����D�S2P��n0?��?�d��~萾�s,>� ��G=�D,?��?�m<.u�>�$?+*�T��?V^>�5>�>�>�U�>d�>s®�1#ݽ]?ܑT?�2 ����>�>����H�|�� d=�+>*�4������\> e�<,썾�+~�����T�<P,W?Y��>�"*���}L��)| � A=r�x?�b?{��>Dk?�2C?ͬ�<VK����S��]�Y?t=��W?�7i?	>�偽o2оmi���5?A�e?cxO>�i��꾧�.�1D���?��n?�]?�o���t}���P��ʕ6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������i�->쒣�X��?5.�?F�̾�	>C�����A���\Y�=y��=����(��%!1�X$���N��˂�-K�=Ihz>|�@�~�'?������:�ȿ�)���9��]��<��6?Oҥ>�×��n��>֔�"�k�#� �5�u|��M�>��>Ͳ��V����{��q;��"����>���	�>��S��&������5<[�>���>��>�*��d罾*ř?�c���?οA�������X?-h�?�n�?q?;u9<��v��{�-s�Z.G?��s?AZ?�o%��=]���7���t?��o��u�4�#�p>�Y���u?w�>Hme�/{t�����|�2?"�=v-E��п�ſJ1�ɗ?@��?v�ž/�>]��?7A?(�+�CO��g���A���d=<`v?^��>������K�P�+���A?�&6?�.�!n�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?m*�>f�?N��=e�>���=����÷0�^#>�a�=X?��?�M?N�>���=��8��/��XF��PR��)�t�C��
�>��a?w}L?�Hb>%
����1�t!�m�ͽe1��鼊b@��6,�k߽�<5>u�=>(>��D��Ӿw�?}k���ؿ�h��8l'�)4?̓>��?g�� �t����?_?�o�>�6�/-��+*��o����?�F�?�?q�׾��˼W>��>�D�>{�Խa��������7>q�B?I2�zA���o�<��>���?%�@[Ϯ?Y�h��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*����z���|[����}��P�;�fA>U\>0Ͻ-}=s�=p˼�rl<���>���>8�e>��>ޓ�>Z�_>���=��|�ژ�.&���d���EX�х
�NOѾT^_��6辇�,������꾻]�=MT�#�J��"���9�9s�:>�+X?� O?*�z?�?S}뼿J=gh���R;Ɠ���7>��>��B?�"F?"�<?��>��}�d
�������㔇� ��>��L>@�>LH�>/��>�h7����=�{>��q>ٯ9=7��<r�9� �=X�r>�v�>� ?���><�;>z>!̴��,���i��x�sȽL�?gD���K�&@������<���_�=�.?ܠ>���
п߿��^>H?0ғ����)�a1>��/?�W?�>������S���>r0�6�i�G��=Ji��mn�V*��OM>!�?X>ǖ>�B�~e5��!t���T�>�>?��۾���������)�_�꾥��=��>@~ ���5�6���?r��!�q��=��<?�^?�L��3߾������h�>�|>�V�=�k>3�P>|���?W�Z����	�<�Z�=GfA>�X?��+>6Ȏ=�ۣ>�Q��v8P�i}�>��B>D8,>�@?�/%?u��l֗�녃���-�+*w>�`�>�>�O>!WJ�կ=sj�>��a>%�����3����?�	WW>��}�6~_��hu���x=��#��=/�=	� �.�<��B&=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿa �>Bָ��̙��u���Re�r!ҽ��>p?�:���*����%�@?j��>T��z����{̿�p���>�C�?mw�?�s_��m����D���?m��?3?~?g�p>��x���U��=�D?<2S?o�>#���s����>���?���?4�>���?o�?@?�*&���#��p��.I���/g>
�=m�
?~p~>B���x@.�㞉�]�_��\T��K=��8>��=I��>���.v��}J�>�d�-�꾡��=Jy�>L�=ؽ9>���>.��>��?��>�S9<r��j̾��ɾOZJ?�D�?����V�E�f��=_��<󃰾���>�<?���B���?�><2Z?'��?��\?���>`�錄��ƿ%h��
:���>>),�>���>�yb</��>=aԾ�,��ݿ�>���>|�/��ѱ�5y�����=���>�'?
�>}�C�<� ?�#?ZNk>�> mE�"*���F����>���>h??��~?s?�.���N3�B���ǡ�$�[�!M>��x?�G?���>�������V�2��I�7r��]��?�jg?�N潍�?�#�?�M??��A?�g>��)�׾I3�����>��!?���A��M&�V�+~?#P?	��>�4���ս�Fּ���O�� ?�(\?yA&?ޜ�f,a�j�¾�8�<��"�N�U���;�D���>a�>0�����=�>װ=�Om��E6���f<�l�=��>��=A.7��x��0=,?��G�|ۃ���=��r�?xD���>�IL>����^?hl=��{�����x��	U� �? ��?Zk�?`��@�h��$=?�?S	?o"�>�J���}޾6���Pw�~x��w�U�>���>�l���K���ڙ���F��X�ŽBl�	=�>��>{� ?��?�?i>���>�o��Y|>���ž����h��*�;�E���.�X��qԻ�����=�P���餾�d>�*���^�>�-2?��>�D�>{b�>ѳ]��iY>iQ>�>^�>��Q><�D>A�>߇�y��Q?�ž%�Ӎ辪A���D?T�c?6��>�k��ƅ��.�K'?�ړ?���?��v>J,g���*��D?�v�>A}�6m	?�2P=�h:��<����\v�����fs缾Z�>��ӽH|8��aM�4Zk��-?�i?ڌ����ɾ�ٽ44����r= �?��(?E*�R��ko��MW�i�R������h�d�����$�&�p��я�W��� ��.�(�:�'=�m*?��?���"�J2����j�/?��f>�^�>��>��>��K>�	��1��3^�'Z'��Ԃ�J�>�6{?V[�>2hI?��;?3�L?YFS?5��>*�>���a�>�� =\V�>�\�>��2?��%?�:?� ?v�1?�>���[���)ݾ�S?�?��?Z?�\?M���/{	�Y8�;'gм+^k�񜂽���=�F<�q���ڽ�=w�v>q\?v��C�8�t���H�j>>u7?���>��>�%���G����<x�>%�
?�;�>�	 ���r��j�-]�>���?���:q=X�)>�=�܅��:Ժ�d�=jüϰ�=󁼼�:���<�p�=)��=�5~��_����:��;���< u�>6�?���>�C�>�@��/� �c�� f�=�Y>>S>�>�Eپ�}���$��u�g��]y>�w�?�z�?ƻf=��=��=}���U�����G������<�?=J#?(XT?`��?{�=?^j#?е>+�jM���^�������?
~+?q�>$%���ʾ|�����4���?[�?'_a�����H*��!����ݽhT>�$/��~����[�C��s��%�O���8��?�n�? 5��]6���� ���^����B?� �>ާ>�{�>�2*�V�h�λ��=>A��>AQ?��>TQd??�l?^�U?�u�>;������y�>�`�=g�6?�Oi?JN�?Ȣp?�(�>��>��M��v�7�ټ���p�:J��y�=o6i>�t�>S�>�G�>�|=Xk�i�R��p��<>F�>���>�y�>��>�A=>�K���D?���>�˞���	���b��Nz�C�ҽ'�?�Ӛ?�L)?�f>�����C���۾���>���?��?K�$?4E��^1�=.%=���Ñ�y�>���>{��>�?>�b)���>���>�/�>Sɜ�ap"���%�T�z�b�?~OH?lI>nƿլq��p��ӗ�dNe<b��d�Sʔ�G�Z�4��=���M��
Ʃ�C�[�奠��x��Uᵾ+�����{�K��>L��=���=��=�t�<�yɼ �<!K=3��<��=4"p���m<o�8�*Eϻ�������\<��I=A���˾��}?�;I?�+?��C?�y>�:>�3�M��>�����@?WV>��P�����N�;�<���� ��o�ؾ=x׾�c�ʟ��H>�`I�/�>�83>�G�=�K�<��=�s={=�R��=+$�=�O�=xg�=��=�>SU>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�6>��	>T�Q�N^/�h�m�?ts��W���!?@t:�Ѫ;�E�>B��=?�⾮�˾�_=�=(>�z-=��!�Lv[�4�=�����b=��y=zf�>�@>Da�=K)��wX�=�eT=8m�=�6d>�B���Z�K�p��R=�8�=`_u>
�.>��>��?�1?Vh?�t�>��
�q(ʾn����W�>� >��> ����=���>ۥL?�EX?5+O?��s>RP����>G�>�J:���|�־���Ee��w�?	>�?�ɚ>o,�=�>�S�)��l4�c�
3?]�j?J�'?a.�>�0����¿�l/�@�W�͛�<Ϗ>��>UP$��=��}>^`��5�S#��H�3?�u�>��>(�?���>��&>t �>��>�k>=s��<DA�=,�<�:��}4<���2�Qno<�X�=mq۽i�c�\��䉽�宻:��=-+w=d�>���>�Y>GL�>��>���X�>-a��d�W�V˃>(f��6F��v�R����1���Y��=��d>_�y=�Ǐ����>�	>/?>D��?w��?�=��ƽoj���t��`~�d���7��=��Y>2?��>�#�éV���D������4�>o��>���>��>�VG�,�X�<�>��&�)���+?�����F�=\�Id��X�e3��
�\�Rd=�XP?3���VK�=��?/"?�b�?�b?W�þ�ھ�>�:O�>$>�2J�o�����3?]A6?���>���n/��E̾&��fٷ>�=I���O�_Õ���0���_ͷ���>z���i�оD%3��g�������B��Vr� �> �O?B�?g=b�,U��ARO����,(���n?W|g?K �>�I?F??���u�.u��dO�=o�n? ��?�=�?u>�ý=����ZK�>�"	?J��?���?zys?_?�Fd�>n�;ٱ >�Ș�]��=F�>Y��=(�=�g?��
?��
?tN��k�	�����^���<z��=�k�>~�>{�r>X��=S�g='c�=�\>��>���>>�d>��>�A�>��r��;#��9*?[�C=���> �j?���>G�=�|q�a%8�����5Y��_G>�Ѷ��X.�}㼂ݽ>�>Yp�=�%�>U�п!�?p�%>��� =>?D���|�=��>ݹ�<��þ�?�W?\2�>fZ�>nW�>�KI>�c�>����ܷ���7>��H����O�^�d�����j�>� ����U��R��H <>�������a	��Cp����E�2�!v�#�?k�!��eW���$��C��V ?٘�>�'@?!�;�琽d�=��!?�G�>�D�A՘�_A��`Ǡ�v��?���?�;c>��>J�W?"�?��1�!3� vZ�+�u�d(A�%e�M�`��፿����
�I��/�_?�x?)yA?�Q�<,:z>O��?��%�aӏ��)�>�/�$';�l@<=�+�>*��$�`�{�Ӿ��þ�7��HF>��o??%�?|Y?;TV�ѣm��#'>6�:?}�1?BPt?��1?��;?U��\�$?8r3>�F?o?N5?I�.?n�
?�	2>��=������'=3�� ���q�ѽ�uʽ'��<�3=+i{=1�ڸ*�<�=��<�t�	�ټw�;����Y�<:=y��=��=B~�>9�`?�H�>�a>��D?oiʽ:E*���t���A?!�=Hh��h۬��؂����O��>e�v?l��?��Z?!��=�&�o�b��:>m��>U[>C^�>A<�>�m�����=UQ!>���=b�>����K�Z�!��þ@�>� �>���>�0|>p���'>�|��`1z�@�d>��Q��̺���S���G���1��v��Y�>%�K?��?֜�=�_龪-��TIf�0)?�]<?�NM?��?��=��۾��9���J�%>���>�\�<�������#����:�-u�:�s>�1��m���J�>�v���!�(��W�j� 1��[ֵ>T��)Ӏ���V��{U���=>S�S=v.	�|�N�n����}��`CI?M��=,ꗾrxǽ�\��I��=B�>�5�>9�v���9���R��eѾ�ٵ=x��>W
>�<�5���f*��s��n�>N;E?P_?zr�?8���Z�r�K�B�����Z��R��� ??Z��>�J?��A>�}�=���W��a�d��G����>�j�>����H�)$��CX���=$�~��>�?_ >�?��R?�1?�-`?*�)?�<?��>.�������)&?��?{a=we��{�H���5��qA�r��>~v?�I�#�>i~?��?�y ?4�S?}�?��9>]��Q�K��c�>���>��V�ZC��\�?>�=?̌�>d`?L�?S{H> �3�ȩ��Ľ/�=��>0�.?�+?�%?�L�>o��>˙����r��f?�P�?T�?[Hw?ND5�M�?�6d=��?z���F6?�z6?�?%�k?�"Z?�6/?���>�R=�ؽ�y��9=
�}DE����>=>���<̽؏;=�� >~-�.t4�r�S��U4�qNx=�=���<�_�>��s>�
���0>��ľ�O���@>�����P���ي��:�*߷=���>��?d��> X#����=p��>vG�>��T6(?�??l";L�b�!�ھ&�K���>b	B?���=��l�����Q�u�3�g=9�m?i�^?y�W��%����b?��?Q���/���kþ�1�K�;?�?�D��	q�>�Ӛ?H�J?m<�>
�ؽ��?�����l���ߪ�q��=0��>�Y%�c�M����>��?EE.>�n>��$>�f����C�����!?���?Q��?��?B:�>�������j�ɾ����@�w?��>�N��F�+?�ɽ��ھ<��L�?�L��<KZ�|_ľ@��A����������v��sk�=��?��?3mX?��u?�D�Pqo�؏W� ���B��I��o���G�;�J�:�X�ջz�߱���~���4s�=�^�RT�OM�?8�?I�Z� ?����dŬ��ct>�%������\?=����;=�:0=C�V�w�ս�բ�f�&?�C�>�>eXJ?_+r�g 2�i�1��7��žh��=��E>���>��>�#n�ag#�k����J�e�R�.��Jv>�vc?��K?��n?�`��$1����ʘ!���0�jQ����B>->`��>��W��~�"-&�&L>�9�r�)���x����	�vX=��2?2�>���>�M�?��?{	��B��/$x���1��y�<x!�>�i?�8�>�>^Ͻ� �f��>��l?j��>�>p����Z!���{�1�ʽ�%�>�߭>7��>z�o>��,��#\��j��d����9�rt�="�h?�-�`���>bR?�%�:��G<_|�>�v��!�����'���>^|?}��=��;>]ž�$���{��7��QJ)?3?�䒾]N*��x~>d"?ߡ�>�!�>��?^i�>8�¾����<�?u�^?�@J?�AA?%��>V�=�����~Ƚ��&�� .=L��>c�Z>��n=��=����<\�J��UHE=��=�lɼi3���u	<�d���	C<��<��3>?/ӿ
	@����.S	�����J���v�6g<*k[�����#�Ǿ1\��z��B�����AO���ɟ�J+�������?��?��ǣо���A���I2����>�Ͻ��Q����Ὣ=e��Ef����c���/؄�Fd�P�;��I!?��9�͠����]����>��3? �?�4վ��G�P�Z�0}>�̮���m=� �s�����̿����n;?�}�>����d="Ӻ>�{s>�m�>�n�>��ξ�(��$��=3?t�D?�f�>"�����Ŀ����c=���?�c@�|A?��(���쾮OV=���>�	?=�?>EW1�7M�W���,Z�>;�?���?��M=��W�"j	��ze?l�;�G�Ä޻u��=!L�=JZ=���ٞJ>Ic�>����fA�.�۽��4>̅>�N"����v^�ђ�< �]>�fս�Q��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=s6��{���&V�}��=[��>c�>,������O��I��V��=f� ���ĿB�.��^��g3=Yo<��ȼV�߽q�ǽ�V��-:���ϡ�F��T��=^ >kU> z>a�>S�`>�DW?��s?���>�!>��ݽ�����<پ���<���d�|�����v����ǾrH ��H��)5��.��0�����7���>FL�ʃ���gN�k�x�˧��U?*�A>9S�
�P��>5v��T�����%��M1,���#�5�$�ED�?O;?�^���]�]$��y-��$�<�J?�������㑾�i<>����I�F>S��>��>���T1�(K�k2?��?IBľ%J<��I>���,(�=�<?���>d�3>cv�>}%?2&ս�+۽�K�>G 9>�%�>v5�>�i>N*���3�Sa?�I?[�~�	�*��c�>ȏ�V�}�s�=��>�Ys�UR>P��>�_�����`��d/�x(�=!V?K��>�%��l
������o����=Y�?BJ?O�>2�j?"{;?$��;�2���3�Ū��'>	._?��e?��=Hq��u���;���?�4?�8_?��>񟈾̏��� ����M"?Izu?�K!?�r��q�y�\�3��	A?��v? s^�vs�����P�V�_=�>�[�>���>��9��k�>�>?�#��G������rY4�$Þ?��@���?��;<��Q��=�;?k\�>�O��>ƾ�z�������q=�"�>	���{ev����R,�c�8?ڠ�?���>��������;>�Þ�]��?#5�?R�����<��.�Yiw�[:־�|&>�8�C�����d�ǭ1��M�[˸������?�_=U�>�@���C�?=Aؾx��H�ƿ�x������t>?�G9>	u�ԧ��`��٧s���I��3T��/��H�>��>!�J����{�Ds;�j��b�>x
�� �>��S�D��잟�dn5<��> ��>���>{7��&㽾&ę?�\��G>οת������X?(g�?n�?�n?�E9<��v���{�����.G?0�s?Z?��%�DC]���7���j?����_�K�4��ZE�oS>.&3?-��>��-��y=�>�7�>�>�X/�`�ĿW���q&��SӦ?-q�?�X꾼e�>���?�+?�5�82������5+���G���A?�N1>Id��%4!�T�=�e����
?�0?�<����]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�U�>#�?;��="H�>���=���jE��`#>P]�=z�?�D�?"�M?��>�_�=�B8��.��2F�_�R�1n�ݤC����>��a?�mL?�\b>6巽�1��� �9�ν֧0��鼳�@��,��޽�5>�>>�>u�D�VIӾ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*l���:���\�:(¾���=(�>!��=�0K��jT>�5�<�5ջrn���=}"�>5��>���>�o>�F>�DH>h�������=��:ӟ��Y"��4	�F.��VI��� ��Ι��������ξ����]��G#�
?0�D����;��8>�>O?*3/?'�w?��>�,���9;�R�� �!��w�R>t!�>?E?P�???/?�1�=7F�T3S�$���O����t�>ݛ>���>hh�>�F�>�E�u>pS�>P�>+�=�<<��׽��=�G.>��>��?�P�>N�0>%N>ʹ���a���ks�����,�.��?��i��n�񳝿���_�����>��?)4�#��qĿ���ιG??Ht����J�
���=�3?�`?2��=-���[�k�Q8�<�-�UZ&����="�'���^��G���l>w_?��c>��>$�4���=�\�T�����9��>J�B?����Iz�}�b�E�F�ݾ�i`>8��>�JT���%�§���+~��:L��)�=f29?/` ?.���bҝ�PE�
*��`>��W>�Rj;'O�=��T>u*_������G���`=v�>pVZ>�n?�2>�Bi=�٧>�$��b<H��Ϯ>�I>�J1>S�D?�l)?�DT�I]E���x�jj��p>�R�>ߵ�>4>]�S��w�=B~�>�!o>Ϲ���3�>���Ԍw�j�F>���*�_��ɽ�|�=�6M��F�=Vtu=�S�&�C�
�"=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�g�>lu�?Z������u���#=+��>�9H?/T����O�J>�Yv
??	]򾧩����ȿ�|v����>f�?e��?Y�m��@���@����>���?hY?�ki>6g۾�]Z�H��>�@?zR?��>�9�i�'���?�޶?���?�I>w��?h�s?�l�>�Hx��Z/��6��Ԗ��4p=1\;Vd�>�W>�����hF�Pؓ�_h��r�j����-�a>�$=��>�O��4���8�=����)I��)�f����>)q>��I>2X�>�� ?�a�>���>2n=�o�� ှk����L?M�?ʋ ��9�&=a�7��W�>qg�>�佄���M�	?��P?��V?i�L?��>ĮԾ�Y��b�ڿ���@{E����>a�?��>� @>|ܽ>U쾤�վ�_�>��>TE8�z�������?��c>a�;?q�#?�:e�¶'?�X@?�:�>4��>�A]����� xi��h�>�o�>e?+�x?��/?�9�V�f�uĝ�z��a�Y��r�=�Lh?�h?� ?a������Y5�>������?EHN?�/ʾ9�$?k��?_?e?+e[?:f?�d����ž!�S���Q=��!?���C�A��H&�
���t?I@?M��>�1����ս�<ּ��w��2�?'\?6@&?���n6a�1þr�<Q�#�6LU���;8D�W�>��>뗈�<O�=>���=Zm�E-6�h< g�=���>51�=57��Ǝ��=,?CG��܃�i�="�r�5wD���>�aL>���p�^?�]=�9�{�#���w����T����?e��?l�?����<�h�� =?A�?�	?#�>LF���o޾ϒ��Uw� }x�1v�1�>���>��k�a�7���i���zF��K�Žaa!�wh�>~�?qպ>�+�>t�">� �>�/���Gd�㲾,'���^��)��6�бD�E�����'
�=��ϾJ+����>P�ɽ\��>�8?U\.>���>�u�>�+�<&�>'=p��=_^�>&�q>��F>��>�d=��
��KR?����&�'�@��|����2B?�qd?2�>i�p���d��,�?h��?Cs�?�;v>4h�!-+�8n?�=�>���&q
?qY:=�:��:�<@U�����5��F�U��>BE׽F :��M�xnf��i
?L/?����̾�9׽Ȳ���ɩ=G��?�5?`W?���M��2|�?\��\F�O�"=�[�s��<5;�����BS��~���A}���t&��=��#?�ג?� �q��SI����n�p�<�寅>H��>�&[>���>��>^d
�)&���_��/�������>��m?�"�>i�.?�[%? qa?k�@?���>��>O�A0�>:>�4�>z��=c�~??F4?|�9?�6?�|&?U�g>[e=�c�0���&?��&?�]&?M�0?���>uM�Viн8j9�x0�-=����5>{ca>*�$=�8h=����*��@��<pX?֖���8�����j�j>�7?J��>���>���,���<Y�>z�
?�F�>O  ��}r��b��U�>q��?����=��)>���=
����Һ�`�=Q���(�=�;��u;�02<+��=G��=.\t��ҁ����:+[�;c^�<�{�>��?���>�B�>�A���� ������=�-Y>�HS>�5>|<پ�z��_!���g��jy>�{�?Q|�?��f=��=�h�=\u���;������뽾���<K�?)>#?VKT?⍒?P�=?�j#?
�>H+�LJ��a��a����?X%?���>õܾ����@��QKG�~�0?D?�7D��Ԯ��T�.z���݇�A=HS_�Ce���G��֠��r�=q���N����?�v�?t]�;15B�6,"������Ja�?�>�m�>�P�>5�o� |����:>`�>�;k?TA�>��K?X�p?�p`?��[>��.�쑩�o������1H>�J?�}?)��?4�n?)��>/}+>6���d�־bX�!����������.F>��z>�g�>��>aY�=Bi�n�K��-��Z>_
A>|	�>X�>��>fK�>��{;8H?3s�>%)ž,v �I���̏����A��?��?��<?��>X��n2C�N���>~��?o�?(G?�Sx�nC�==��rE���}/��$�>i��>���>�_>!�#>�>�]�>W#�>(QU��]�;�%�������>��A?���>��ſhq���q��M��*5<链�0d�Mȏ�IYZ����=������I��s>[�Š�Z����;�������z����>�z�=E5�=���=?��<�Լ4��<v*P=��<��=,uo� �p<'8���A!������Z�N<zAH=�j��s˾�}?�2I?��+?��C??�y>�>�4��s�>x8��H?�$V>�P�B��#S;�ۙ����9�ؾ�׾5�c�˟��a>LI�r�>,3>ҝ�=;�<���=�s=�=��M���=_��=ln�=9s�=�7�=��>�?>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�7>[�>��R���1� �^�'�d���Z���!?��:��;Rv�>�l�=d߾0�žj�-=�4>q�V=�E�n\�o/�=��y��:=#�k=���>�B>��=�r��k*�=�F=n��==�N>����?1��*��q8=���=Nb>�#>X�>f�?߼?�KO?_#�>gcw�3�ľ�U��w.�=���>n�?lc�=�x>sw�>7dE?�^B?^�e?�V�>�3r��>3֨>�+�E�^���tǾ��<�ܓ?��?\��>��r� D��b��b?�'�r�NE?R?��'?���>u��`�޿��8�;y0��(K���=Qct<|~V��>�==F���ʾ���>�ܴ>��>�T�>���>F�>��>F�>B�>�������=ϔ;�r�;>�=<F�=�<Q���9��B6�����2����=U>�=6S��F�=г=o�=;I�>��>�>�3�=T����0>����˫M����=C$����A���c��t~�h/���6���?>q�T>KM��Jc?Z>.R=><��?�v?t�!>8L
��վ]���0_�Q�W��,�=AK>�;��m:��_��NM�g�Ѿ�׺>,Dx>x?$@�=w3��]��=�����y����>����^&>|0��u��w*���מ���m��C<���F?�-y�}�<���?��?�Ì?�g?ٰ\�D������]=��o>C�9���S���8ٹ%?
h?Z��>���kn)��G̾p���>:MI�y�O�P�����0�-��{ٷ�"��>����L�о[&3�
f�������B��Qr���>f�O?��?�Lb�U�� RO�N������k?<|g?�$�>�K?6@?Y���w�i��L��=��n?��?�;�?!�
>V�=���.��>}o?�Ŗ??k�?�{s?kHO�=��>�\<y�&>|��b�>7v>V�=��=�t?W�?	?���"?	��	�~� �X�Y=���=�i�>j�>=Ik>up�=�^=*(i=gU>|͖>j�>4�d>���>TJ�>F�����/��m?�*/���>T^2?�3>1��<-�j��ul>�U⽣MM�]*��1W۽}GA���Y�	0�<;��<���x�>�/ʿ숁?~��>?h����2?�\9�:N8��'?2��>H�⽣�?�I�>��=���>�ϩ>
��>}��>ǿ��~&Ҿ>���@S"�^�C���R��Iξ��>�(��0�0��z
����� I������x�j�Aw���C<���<���?+����i���)��"��v?2�>-�3?y���Mӂ��	>���>I��>�B��Jh��)������ċ?j�?�;c>��>P�W?�?ʒ1�%3��uZ�&�u�w(A� e�S�`��፿�����
����%�_?�x?&yA?>S�<":z>H��?��%�Rӏ��)�>�/�-';�L@<=�+�>
*��'�`�u�Ӿ��þ�7�IF>��o?@%�?zY?`TV�Sd��N�=F� ?��N?�3�?HNU?5�C?�ߚ�ۘ&?мD>��?�r�>�FA?k�0?+B?w�>�S>n��=L0'=�C��~��V	�"
�+`^��J:=�g�=��+<Ǝ>wp*��C4:���<�튽�=#����=�p=Ǯ�=���=|
�>�]?ĳ�>���>p3?֥!�~p7��К�~/?0�=Ho��鈾[4�� 6�l>ji? �?��]?��d>Y�>��*F��>GN�>�+>#s\>D�>4o㽥�G��}=�J>�,>eB�=�"��v���
����qSA<�A>���>�C|>�(��j�'>t���*z��}d>��Q�&ݺ�`�S��G���1���v�b�>�K?��?ν�=�b�騖�qDf��#)?�`<?�VM?��?6>�=��۾��9�P�J��	�s"�>�<�	�����v����:��a�:��s>H ������)_>�����vl���H�
~���e=���D�=��
�zҾč}� ��=M�>�@��i~��ʖ��h��p�I?�́=&y��[�V�������>a��>��>�8�Tq��_>�S�����=av�>I@>�C�����ۢF�=w��K>�L? 2a?��r?�ό���m�"�K�E��[�������>^��>%K? >*��=瞠�0���?f��M����>�?�	��N�P�3���B��Q|3�`P�>Qh?�ݫ=���>7�X?�I?N?�m ?n��>�F>̺�
о�B&?�?��=��Խ��T�� 9�QF����>E�)?t�B�θ�>w�?��?��&?ՅQ?�?��>�� �gC@�F��>Y�>��W�:b��&�_>]�J?���>�<Y?�ԃ?�=>��5�M梾�ة��R�=k>W�2?�6#?��?ͭ�>���>ã���"�=���>� c?)3�?��o?�k�=��?��2>a��>��=&��>%��>� ?FO?��s?_�J?՜�>lI�<[i���󶽒Cr�U���~;�G<�B{=?2��t����r��<i��;䗻��Mh��D��(����;<��>BRu>�Y��5�>]�׾�]��8t>�d�<�^��u!���BP��؍=�&�>�?UI�>BC�z�m=|=�>N��>Z#�G@(?�V?��?�cD=��X��
Ҿ3�l�*ˡ>�W7?�ӊ=ʩd�����Wt�IO�=˞j?��K?�=����O�b?��]?@h��=��þ{�b����g�O?=�
?4�G���>��~?g�q?U��>�e�+:n�*��Db���j�#Ѷ=]r�>KX�R�d��?�>n�7?�N�>-�b>+%�=iu۾�w��q��g?��?�?���?+*>��n�Z4��I��y���$�a?���>s桾a�(?��&<r�پ�����j�2r��᧾Y���s���s���(�X�~��ֽ:��=��?�Sm?�j?�\?�#� g�ؾ\�Dkp���M�E|�W�@�H��x>���D�v�i�d��R�HǊ�Yw=�	��%U�
�?9�3?#���(?���ü�������>T�ʾ�Oi�,o'>���|E�;f	>`�9�X��Jc'�T�+?*�?�J�>-d'?E f�o�`�;X��a�zS㾛��=��#>G�P>bq�>#,==.�.͏��L��DL6�!܃�r�u>w�c?q�K?q�n?2t�?M1�����!�<�2��r����B>q_>.�>�V��0�&�"_>��r����"O����	��!=��2?"1�>���>�O�?��?�w	�}Ʈ�j�w��1��y<�%�>��h?��>�>��н�� ����>��l?���>��>ؖ��gZ!���{��ʽV&�>�>��>��o>�,��#\��j��L����9��u�=)�h?
���a�`�[�>�R?��:�G<�|�>~�v���!������'��>X|?;��=��;>,�ž�$�x�{��7��H>+?��?������#���>y?���>�˟>���?W�>�už�p+���?Hc?�K?F�??���>�~H=�_��@Tɽ:H*�C�J=�M�>B�T>BjO=�'�=����O�,;�J�m=��=W���Ǣ�~�<�S����u<��=hm1>��ڿ��K�.=۾ǹ����F�
�_�4�������_X��F���f����}���@�9��?O��\��X����p�/,�?7��?�Α�e���陿�~�]W�����>ڿr��ow�Tͱ����Ց�!"�`�������EM��j���e���?�耾uu¿����Y��a$?��>H^�?��'��&�]g���l=�c�<W
=�xt�PX��Mʿ?�5���Q?�%�>�����J��P_�>�Q">�U+>�A�>��S�G& �t�%>̈́?��?�c�>5��D��+iʿ��=���?=@�}O?Ix��׾R�=�p�>m�?i�>	9��7
�E�оE�>�è? ��?�~��3d��S/=�gz?U�=G I��:�L�>4�S=(�<� ��c�>:T>�!��"ƽkz��gE�=�ӕ>r��<׈>�Ŵ���m=��i>ڰ$�L�5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�����{���&V�}��=[��>c�>,������O��I��U��={~����ƿ�85�d%�4���B��얼�io�B����f���>��8������*>��<��>�R�>�$C>ց�=�D?��l?���>��ҽ��
�LJ��sn��ِ�矼�!��(VC�zqh������o־?9�e5����O��᪽�^b��"��x�2��R��f(�q#?��/>�Ҿ�8���=*��4�����9��|�=1i4�?n;�W�� �?i�??�Ge��0d��žR��=�>�5??ob8�
������r�=��=&+ ��|�>t�=�?۾�1��jK�w�0?`S?枾��現�(,>� �V�
=�5+??J2^<��>F�$?9�)���߽�Z>4>��>!#�>�'
>S䮾*ܽ0�?~�T?�z��Y�����>ƽ��qx�r�e=B>�5��S��.^>�q�<����Pp�bގ�}��<�:X?�ȍ>��(�n��q������0=��w?*,?V(�>ak?>IE?a'�<s�����T���� �=�X?�f?W�>8nv���Ͼ0ɦ���6?-,f?P�H>H s�|�8-�h��R?{�n?�? 7򼂞{�����&��>6?'�v?�a^�Oh������V�F5�>1E�>���>�9�v5�>�>?�"�6=�������_4�T?��@ϊ�?�'8<�뵎=�*?�H�>O3O�ƾn��򳵾�r=�>򚧾�=v�y��5�,�o_8?���?���>ܞ�����)ԃ=�����?�Q�?C}��E�=���d�s�������=9�<3�/�r�=�p羾V(��뫾��N|Ǿ����Ȩ�>&@��>�dը>�dN�m��i@տ�g�\������M�>�2�>�J��n��_Z��rv��xC�T�.�������>4%>i��=,���ڪ��%S�yӗ=��>ć��׫�>z��������/��<Ԣ�>�'�>�O>�M��%N�����?�3���ο��������O?2��?���?��?1���E���H�I��1����5?�o?�N?�I�=B�۽����qX?Q��Nc�b�@�5�I�#f>`jC?+�?~Z8�6|̺��=>�
�>�>Z�5W�������JϾߜ�?���?�Xؾn��>��?-%4?0b0�Č������2�"��0n>�$?�ý�^���l˾�_������!?��?<ބ��V�^�_?(�a�K�p���-�n�ƽ�ۡ>�0� f\��M�����Xe����@y����?L^�?h�?Ե�� #�g6%?�>e����8Ǿ��<���>�(�>*N>NH_���u>����:�	i	>���?�~�?Uj?���������U>�}?G��>R6�?$,�=���>���=�����I�!>��=7�;�L?��M?T��>��=d�7��.�LfF��R�9Z�nC�S�>"�a?oL?�mb>�y���90��:!�sϽ�/��5ۼ��@�'�0�<�ܽ�5>h>>�>�D��zҾ��?Mp�8�ؿ j��#p'��54?3��>�?����t�����;_?Tz�>�6��+���%���B�^��?�G�?<�?��׾R̼�>*�>�I�>��Խ����J�����7>%�B?Z��D��p�o�j�>���?	�@�ծ?hi�	?���P���`~�<��m7���=�7?m0�q�z>=��>(�=�nv������s����>�B�?�{�?c��>��l?e�o�w�B�!�1=3N�>��k?Ds?��o�+󾗰B>��?3������"L�f?��
@wu@p�^?~����ꚿ(ӾJ,�ln����<c >�Sɽp>n/U=��>	��b�����>XC,>yRq>�ps>F?�>��p>dQy�7���ÿm���	C��_7��r���!�g�޾��޾����[�������a=ܳ�v5ݻ�3��
����܄�[�=v)p?"�\?�$^?��>Q�0�!\�;rY��мx�#�~*�=T�>��5?��G?P;3?�Yw=�����_�����?����}�(v�>˃>��>���>r��>�ށ��G�=��>���>~U�=����k=䊄=��6>MG�>a�>(a�>�x�=�5<>����
��������w�� �?�����q���b��䙾������q<�<?�-m>�}��,�ʿ2��"�>?j>�����O԰�_�B>�O2?��>?��>�~־���<WՀ>G*Y��s���/>0^�=����T&/�M��>�A?Dhf>Z�t>�3�x8�P�P�Nw��6	|>r36?ض�+�9��u�a�H��Qݾ��L>���>	6?��_�Y����!�1/i��^|=�[:?wt?�m������Ʒu�%!���:R>R�[>�="�=uqM>�b��ƽ��G��6,=�s�=��^>�u?��+>ah�=��>��wpP��C�>�OB>�K->�??�$?�[�k	������g�-�?�v>'D�>�j�>>�hJ�F��=c��>Wb>n�b����8���?�uX>6�|�ц_�A�t���u=qH��g�=���=ґ �'<��8%=�~?���(䈿��e���lD?S+?b �=
�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��N��=}�>
׫>�ξ�L��?��Ž5Ǣ�ɔ	�0)#�jS�?��?��/�Zʋ�<l�~6>�^%?��Ӿ4g�>h���Z��F���u��#=[��>�@H?�q���O�ۻ=��i
?�?�P�գ����ȿ�rv����>��?�?��m��5���@�U�>���?�rY?�Ti>�A۾�aZ�`�>�@?
R?��>cF�{'�F�?5ն??JR%>1��?$�t?��>�Ʀ�)�8�|%��|����o=�)�@>O�s>C����M?�.���@����e�b���=�=�Cb=��>諢��Qľ�#�=�D��FW�����Ɠ�>�}�>�Av>�>�>U �>�J�>�&�>	v�<�-ܽ��J�"���N�K?���?����2n��M�<e��=&�^�`&?YI4?�b[�m�Ͼ֨>�\?Z?�[?�c�>P��>>��@迿�}�����<��K>G4�>�H�>�$���FK>�ԾX5D��p�>aЗ>�����?ھs,��fE��BB�>le!?x��>;Ӯ=�� ?5�#?�j>P9�>+hE��7��S�E����>��>mP?��~?Z�?i���IX3�����ࡿ'�[��7N>(�x?�]?�ϕ>ǎ������ΔI�NJ��Ғ�ҡ�?�mg?:��� ?�(�?}�??B�A?�Gf>Zv�A ؾɰ���Ԁ>P�!?6,���A��k&����|?�1?=�>"i��RFֽ ʼ���̔��S�?�2\?��%?����`��t¾���<�A'���U�Q�;�8L�P�>(4>�爽�˳=�>�G�=�Bm��\5�de< ��=�>�K�=�W7�/ь��=,?ٲG�ۃ�/�=��r��wD�>�>�IL>B����^?k=�h�{�;���x���U��?(��?Tk�?���ڝh��$=?��?�?�#�>OI��|~޾����Mw��|x��w���>`��>�l����n����F����Ž�a�>��>��>��?�ކ>)?Cc��7P��k���#�Y�(�Q��`��6!��?�1��)cD���>V���Eھ7-�>Gy�=N\�>��?{��>�i=��>%�]>4$�>T�~>Ͳs>s0N>�<>Xt>7�>��'�+�%��ZM?!k����&�Fw��Ǿ]4?��j?�?�>�!��4ჿ�y���?�~�?��?�U>G l�V�%�#�?��?����?���=R=)
�<`ɶ��9��;���J�k+~>��32���N���a�^
?A#?��D�]^���^�������s=1J�?
�(?��)��CQ�Cko��W���R�����k��C��o�#�(p�̔�������ك�%�(�l�%=Ќ*?.[�?���G[��ϭ�_�k�|�?��.i>��>�k�>Ǝ�>��K>�		�c1�ia]��Y'�J3��ϕ�>�z?�[�>��E?�D<?J�V?GP?�0~>w�>�ְ��d	?U"�<ۓ>���>O�0?�:?R
4?��?#(?��~>g(Ž`���)�ؾ�?sM?��?m��>�?^�~�����Wx	<��Q<�b���l4�=-�:=������ �=��Q>
�?�.��;I�����{>�f0?T�>?~t㾠r}���}>xۨ>g��>R>�5þ닿��d��>�ȉ?�b��}��d4;>Ѝ�=�����"���s>9L��n��=n�ȃ��q�y�>�8=��W���g�,�>TJ�i��=2u�>3�?���>�C�>l@��� �b���e�=�Y>�S>z>�Eپ�}���$����g�"^y>�w�?�z�?9�f=��=��=�|��cU����������<ˣ?FJ#? XT?H��?i�=?Wj#?Ե>+�\M���^�������?��+?0~�>����ʾ��3���?�?o a�^�:4)���¾ �ҽ�->:H/�,@~��毿´C��W�Q���N��;��?Y��?�a=�
�6�A�]���=T��\OC?/{�>�.�>��>K�)���g�&���:>A~�>{�Q?��>n�}?-Ղ?�E?�h>�9J�q��������̽)�>q�.?6��?䮇?x�s?�4�>`�
>x�����R��=�"��i2.�	�l>f�T>#��>TH�>��N>��ؼ��=�8=Ln��2���>���>�w�>{y�>t�> T�=��g?�	�>���i;Ǿ��ؾ�+�����<��t?,tz?��>��">-MϾ t(�M��Tͭ>���?�;�?�A?x�����>��%�����u����=?��?�b�=�K����=�������>�4?6&�&!��_�D=v=�T:?5!K?�� ���ÿ�n�񗉾Є����ܼՓ�Fe�P�X���M��Ri=1󞾸����`��� |�q��iR{�:윾�򬾝ȓ����>QO�=���=DT�=BG=�˻c΂����=��s�����۔Q�Rg�:�ۼf��ǝH���)��Us���)=���˾��}?�AI?��+?��C?->y>�>�4���>�����?X�V>բN�����`O;�����1����ؾ��׾��c�2���]>%�I�Q�>�3>�=�G�<���=�2t=@f�=��Q��=L��=]��=C_�=�h�=��>rK>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��=��=j?b�:�J�J5L��]c�FN��j�#?�%�D	��`g>!��=��̾b�׾w*�;��>��&=�|�<z���>�T�<Ⱦ��=�=�>�R>ה=.���5��=#c�Zj>��>Qˋ=��;�i= �=�IͽN&&>q�>	?�>x�?-3?�~j?\��>��z�[�־�:¾�>�>�\�>�b1=\K*>,��>yv;?��@?�iI?n��>1V�=<��>��>N����g�i��LO���W=d��?�x�?f��>��=�P.���sr>�A�ؽ�?�7?��?�<�>�U����SY&���.�������>��+=/mr��PU������l������=�p�>)��>�>�Ty>��9>�N>k�>�>V5�<$n�=0ߌ��µ<��約=8�����<�{ż�u���e&���+������;���;��]<��;��
=bT�>.>�V�>���=�����א>�4f�+�S�q�:�ȾDA��g���q�w���3�����=���>��T�/4����>&-�>L~T>��?�wz?��>(��z��S����8���h��"!�B�O�G(���3���c�JUV��㶾�J�>�
�>��>��R>�P.���?���=�NȾ��2�  �>�Ș��\c��:��d��響z����e���=��C?�)��!-�=��?�J?46�?,g�>Y|������=.s|�U�h<hz�r���H�pv?u4"?AB�>Jl���@��˾龽mk�>-�D���P�_����0���0�X���8�>(3��� Ҿ�
2�.��v���Q�A�)�r���>�O?4�?5�_�CP���aO����9��td?�h?>��>!U?�?b������~��m�=&on?j�?���?k)>:��=���
1�>?�?���?Vg�?r�o?)O����>� �<dq>����m�=\�>WD�=*�=�
??�?�����W	���r��ɪf���<®�=.A�>���>'ok>���=H,=��=ȟW>hG�>���>�[>�>���>�^�>51�~�?j>��>��\?o��>�A����򽿳3>�a���O��~������~5ڽ<�ļR>����ӽ�� >
��>z�¿�#�?�}�>ԅ�_*?U�����O�>�3>d���>v�>}G�>g8�>��?�`�>t��=$c�=)FӾ>f��Je!��+C�P�R�־Ѿ2�z>�����&�����z��DI��m���e��j�r.���;=�:ν<�G�?����r�k�L�)�C���	�?h\�>�6?
܌������>I��>
Ǎ>�I������ȍ�g���?1��?�<c>�>n�W?��?�1��3��sZ�i�u��&A��e��`�`፿G�����
������_?��x?xA?א�<�Cz>Ϣ�?��%�dԏ�� �>�!/�Y%;��<=]*�>;+��G�`��Ӿ��þ�4�oNF>C�o?$�?SX?TYV�x����N>JB?3�7?�4m?d�<?�=?��C�_�?�|>���>uc	?�d3?Vi,?z�?Z>2>�N�=g�漶r�=��)������������(���M	=� 4=N(>=-�B=�ž;�E-�(���6���?��9,j�v�;��v=خ>��>��#?#2D?r0?R?��_?�f�<�:���߾J�{?�f�=���	�˽�c��%�]�W�F��\?|}�?&5b?Jc�>]�L���M�95�>���>:3	>�N>��>��b���w�>��=w�<��c�<h%>G��@پh���P�4>�(�>�n�>�|>�`����%>�/���{��h>kWN��
��=�V�H�Z�1���t�IO�>�#K?�d?��=���=u����f���(?Ѽ<?58M?�a�?�{�=O(۾��:�b�K��y�s�>�t�<��
��ܢ��d���8:�)u8�,r>����٠�κO>V��RPݾ1h�bhK�ڲɾ��=z%��u��
��/���v����=���=A��N;�h������<?�<�=�ҕ��6��\��R��=mC�>��>_͉�����c�L��Ä���)<� �>%�u>O&���g��(HP��G�%/q>�79?�b?�?�?�U���i��C"�˫پ����dSG�iB�>\�P>�W�>X�X=���=:���[s���`��:��	?�?��ɴn�bھ��Vo$���?�M#?L�='�?��~?�?!$C?TD?��?��|>�䲽>���%K&?�?�y�=�eֽN�U���8� �E�o��>�)?�
D���>�?��?�g&?�Q?��?�>�� �lC@��C�>�>��W�n���$^>>�J?6��>{@Y?�܃?{+=>f�5��e��ˆ���f�=�� >3?6�"?e[?萸>̖�>Ei����>���>y�V?���?em?��=��?v�2>���>�K�=h�>;��>Z?�Y?�{�?��7?*�>,�a���Z�	�������;53�< �M=P�>O�Ē��C����2;�-4ǽ�<�Ń9���<$�P=���>u7W>������1>��ܾ#i�P�s>�1�"}��h�ky��'�=Wv>�+?ϔ�>�P ���=Ƽ�>ɶ�>�%���4?�@�>�?p݅=�Xj����'q6���>2Y*?��.>�(j��/��}U��^I�=K�t?��J?O����ܾ<�b?X�]?~d�#=��þ��b������O?z�
?��G��>:�~?��q?>��>��e��6n����Eb��j�w�=!p�>%Y���d��9�>e�7?)Q�>��b>�3�=4u۾��w��h�� ?*�?X�?2��?�(*>��n��2�R$��/N��f�Z?2��>?���ϱ&?��ü�;�ð������SӾ����f���n����l���6�;����+ֽI�=�?�m?��q?�2\?����]k�Zyh���y��aR�x��l���>��s8��W?�.�`�����ې�[�W=�]��B�C�)�?�*?�J����>)��(n �Sƾ�HO>������4���=�è��7�<HP�<��t��]*����	�?��>�F�>�e9?��[���H��>��4����>��>_�>��>����m�]��O�⾽�x�r����f>;b?��O? om?�p����6�"����#����c���P�6>b�>�@�>Z�2�f��O��i>���q�=
�Q#����؟;=k�8?�)�>��>r�?���>r��4墾�9w���-�����̃>}�R?Ĕ�>�x�>���<��L��>��l?��>��>����sX!��{�D�ʽ0�>�ޭ>b��>D�o>}�,�e#\�j��ۂ��?9�p�=J�h?�����`�I�>2R?%��:lH<	~�>v�K�!�x��N�'�6�>7y?�u�=�;>3~žT"�h�{�C7����T?��>`�E�%��q����D?�H?��>[n�?N�>O�3�^�9> 0/?.˂?�CV?�J<?�J?Z�=6f�'�̽2*T�6�ѽІ>�c>/n=ܑ=�D�0�V�"��뱘=n����.h��c����T����pM�=�Ԇ=�|/=���W�d�g|��p��D������ā���Nܼ�1��3:V��7h�{f���9��� /�p��<�P3�`{�z>T�%K���?A��?���pP��g���a��y�x��>�혾 �Ľ��T��q��qȋ����� ����$��jZ��	i���e���?��@�(+Ŀ����U����>}��>��?��1�"+'�u^��~��>�t��G%�7^�E����ѿ����J? d�>���¼��+6?��?z��>�=����������>n�D?�W�>6��>� 2�S�ƿ�y���>���?˥@�8B?�)�3��-�[=�f�>KH
?D�E>�"/�3�{���i�>�u�?�P�?H\=W�V��Z��oe?��<*�F��|���V�=���=B =���K>Yw�>��VY@��Wֽ|72>(�>p!&�Y��V%`��(�<B�`>&̽�F���Մ?]{\��f���/��U��\>��T?�*�>�H�=��,?�9H��{Ͽ��\�,a?Q0�?!��?�(?�ڿ��Ӛ>��ܾ��M?B6?e�>�a&���t�(e�=�2�C4��b�㾽"V����=ե�>�x>b�,����?�O��������=��%�Կ�8-������c>�3���pI���r�R���x�#���	��"��τ��(ڼr�D>�jo>_��>���>�h>ȿ�?�Xq?�L=%��=59��/f�?�;�=,����>����ǋ��Q�����S�ž �������ξ��.�4�=�Z��h��3�$�z�r��	"�U�?��8>����B����=����ǃ�0y`�2nK;!'����Q�%o��+ˋ?��>?U�\�U�p��	��)��ཱིnn?g�_�o��� 2>����{=��>Z8��+�no0�5�8�%^0?2�?EԾ��:����*>���N!=��+?T�?#�A<��>�$?�m+����2�\>5>P�>z��>�k>>��Ipܽ�?�sT?���;����E�>�྾�T}���b=�i>ID6���0�\>w��<ꀍ�EV��΍�ض�<�'W?N��>��)�&��N������3==�x?��?�1�>t{k?��B?(�<Gc��B�S��$�mw=��W?I.i?�>����Yо�w��*�5?�e?5�N>�fh����,�.��R��?��n?�Z?R����o}����\���r6?��v?s^�xs�����L�V�g=�>�[�>���>��9��k�>�>?�#��G�� ���{Y4�$Þ?��@���?��;<��X��=�;?k\�>�O��>ƾ�z������8�q=�"�>���~ev����R,�f�8?ݠ�?���>������k��=8����?%�?�J��E�<e��L�u�N�����O=��=Ҥڽ#b'�?꾮�4���Ͼ}��������=�ō>��@q������>��W����/8˿u�t�񷾾�:�(?�*�>�+.���|�� D�n``��}U�B�)���j���?��R>�
�=\���ξ�������[T>Hu%?��@>~)�=h�	�ES{>q�<�Jý?k�#?X��=�Ů��۾Ϗ�?��)�*���c�w��o3��}?�٫?|D?z�5?n�>�1�4�=�z�>TCl?��\?;r9?���=oi�<OT}���c?( ��L�]���5��u.�b�>�?!˫>��/�d��=˹p>��>ݘ>"a�ǿ$����J¾�?eQ�?����?�~�?'?P�6��񆿖����R�$�P=�-?lC>��˾��6��k���k<�d%�>t�?g _�U�0�F�_?ʚa���p���-��ƽzݡ>k�0�
b\��!�����$Ze�>���8y�j��?^�?V�?���� #�=5%?h�>񡕾	9Ǿ$>�<�~�>+�>f1N>OX_� �u>����:�7e	>��?�~�?�h?�������b^>t�}?w�>/�?|c�=�{�>�;�=���I2�	�">�T�=>�>�+�?�M?tG�>�]�=+�8�I/�OQF��=R�����C����>��a?��L?�tb>o���91��� ��Iν�1�n��@�.�)��x�4>�=>��>�D���Ҿ��?21 �39׿h�������7?kCg>3T?�J�e�U�4-<~(V?�0�>���A���9������<�?&��?�?+�;���;T�>D�>b��>C,����ҽ�B}��M>��;?� ��������s��3�>/1�?ۣ@��?��^��	?���P��Va~����7�c��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?Qo���i�B>��?"������L��f?�
@u@a�^?*�hֿ����dN��K���h��=���=��2>	�ٽ=_�=��7=��8�+<�����=k�>��d>3q>n(O>�a;>��)>���H�!�r��X���K�C�������Z�@��Xv�Rz��3�������?���3ý1y���Q�2&�_?`���=<�M?!Oe?!aj?�]�>�'��@�>� ���k=��1�ݡ�=�3>�&?��J?y�'?}zD>ή��vd�OCg�@�¾$���i�>�5�>�>���>-/�>����O�=b5�>�Γ>pLA>�Ӊ�ɖW�@	��}0>��>UV�>�B�>�>W�P>�5��0߾��cg�s�۾5o���"�?7^��nn�ۘ���8	��rѾ{��=a�4?�U�=h!����̿	>��f�:?6Ys�`��/+���
V>$�3?9?��> ����d����=`>�����Hp=�b<��wD��"�>�<?K_b>p�s>&z4��8�7�P��+���}>��4?J��s�B��et�. F�;�߾Q?M>\��>�˻/�|[��P!��ګg�6A�=n�9?Y�>q!��ȃ���ht�{q��ϾS>��U>���<X��=�G>!�X�(~���N�u�=P��=ZB[>�?/:+>}��=��>�<��aYP�)P�>��A>��+><�??�%?��<���Tl��n[.��w>�Y�>���>>�TJ��m�=[�>tPa>*+�
ʃ����D@��fW>��}���`�ar�1Bx=[��;��=��=�h �[>��X!=d��?D��ՠ��Z��O����F?>?7H�=zg�<ܓ�t���֫�*��?	�@��?I����Q���?E��?tڒ����=�'�>�>��̾4sB�œ?T�ѽw��3����*����?��?��ʼ=�����m���#>a�(?��׾�l�>����\������u��.$=N��>m>H?"]���aO���=��w
?]?�S�/����ȿ�|v����>�?��?��m��8��%�?�?t�>u��?YXY?�Ri>V^۾+$Z����>�@?R?`�>�K�s'���?o۶?��?�:>�B�?�sk?]�>���,�;�}���Ζ�����= l>ܜ>>`���H"�����8���怿�B��ɏ>�2@=�?*�*����xMn=*H�Pַ�j�d�k.�>҉�>m�]>;�>E�"?���>�ٓ>��K=��=U�R�iη�Q�K?*ʏ?� ��m����<���=��`���?�e4?2$b�jϾ���>��\?�?��Z?镔>�0�@��򋿿�������< J>_��>l0�>X�����K>6�Ծ?H�ݝ�>��>�F���ھ�(��i����=�>� ?���>�~�=(� ?G�#?�j>h,�>�ZE��8����E����>���>MJ?��~?7�?й�HV3�����䡿4�[�B=N>	�x?|T?���>R��������E�]�I����7��?Rug?K%��?�3�?�??ͥA?!9f>̃��ؾ����\�>�%!?��B���%����X�?�#?"6�>C֒��ڽ��˼N���X��V�?�2[?�u&?����a��ľM��<����Dvl���;��N�_Y>�V>E:��ZP�=��>�H�=q�i��5���q<���=E�>���=�c:��ᓽF=,?ҾG�@ۃ���=��r��wD���>IL>�����^?�l=���{�k��ax���U�� �?���?.k�?M����h��$=?�?@	?A#�>�K���~޾���Pw��~x��v�	�>w��>��l�<���������F����Ž�wl�R2�>o�>��1?#8!?f|>��>�\���U�`\��@ھKb�PF���G�s�Y���0��ф�,��1�&={�̾�W��b�F>wLؽ~M�>�o�>��>�ŉ>��>cĐ=��=�->���=LP8>#;�>�;>���=��g���ڽe?��پ	k�Jľ���{(M?�G?�_�>t��<+~b�A�&�)?���?x��?e�>��P���(��>4g�>H���_8?����WD��Z��=H3վ?�������㜼L/J>��:��A��q]�p9���<?Q�?���ؗ��$f������	cv=��?�d)?@p$���O�ݺp��<Z�3�Q����-]��5���V!�BJl�/)���]���*��L�#���f=�(?�m�?���Pv��㬾@r��^@��d>o�>�c�>�B�>��a>l��M)�@/T�%�(���R/�>uw?�Nm>��A?�fP?يJ?�C1?�]w>˃�>����j��>���e'�>�y�>�m? !?i�2?��%?%� ?���=3K)�}��YD���[,?�c#?��>"�?��>?Hо�`���=fFC=	w/��/�����=c���s���N�ݤ�=E�F>�1?����H1X��B��y�>�A?��m>Gp ?X�־\$�V�'>QN�>��?K&>��.�����F?�2�?�%�����x0�>�>?�/�po�=c�=���~O����:�����½8l>I!�-�R�	�>h�=�c�=�rR>�t�>5�?���>�C�>�@��-� �a���e�=�Y>;S>{>�Eپ�}���$��x�g��]y>�w�?�z�?�f=��=��=}���U�����F���2��<�??J#?'XT?_��?{�=?^j#?ɵ>+�iM���^�������?l!,?芑>�����ʾ�񨿍�3�ĝ?H[?�<a�3��i;)��¾��Խ��>�[/�q/~�����D��ʅ����y��(��?�?�A�C�6��x�ѿ��\��~�C?�!�>\X�>!�>��)�q�g�|%��1;>��>R?Gơ>V�?�(y?+�
?x�ۼ@t��/������G�>��>��?�@W?�?iߔ?��w>A|�<��6=F���������JF�_}��L'I��g�<���=�D�>�޵>3�==�����@ ��1�<���>
�>��>]1�>��]�����H?���>gֽ�����A��J���m���au?�Ő?WA,?L;�<[���C�����\��>�E�?Yɫ?T�)?,�U���=����4z��}�l��_�>qk�>٣�>{C�=H=V�>��>���>!�ϖ��8���`�u�?�F?���=ɕ��w�|��e�����4^��ٖk�ۧ��;�=�g�����	�=x]۾(���ʾ6�h��Jɽ�Af��iٽ#Qo���?ލ�=���=�D>w���߽*�=�=ѻ�8=FvS<f�q��--=
���"�=ʚo�1(>E�c=쬼�'��;�ʾ��y?�pK?�x0?��A?��y>�>c
m��>}���$�?��H>�n��V��zb:���D����ھH�־�[g�y١��q>����>�0>��=Mʜ<-�=ZҀ=�ts=�V߻�,�<�;�=2�=a�=@��=��
>��>�6w?X�������4Q��Z罥�:?�8�>f{�=��ƾq@?|�>>�2������xb��-?���?�T�?>�?Bti��d�>L���㎽�q�=H����=2>k��=w�2�T��>��J>���K��H����4�?��@��??�ዿТϿ7a/>��=L7��٘`���
�D�o��#��UI9�W5?�%���A�>�Ǽ���纾�F�I�>9g�=�W!��X��h�=n=��<^�f<:@p><��=|=>�.�+�=�,�<�����>if�=qT<eܪ��_�=���=o<hB�v��>ж?6�0?��d?O'�>+�l��Aξ���z��>���=���>�=�A>(t�>��7?��D?cL?���>w�=���>>��>�,���m�9V�{|��Q|�<��?�ކ?�.�>lA< �?�f����=��u½�v??,1?�[?F�>���>q'�3�-��럽�I�9{�=��l�z=a�W��)
��n��Y8�=��>M�>�b�>��x>j=>��L>5�>�>�=�<���=�1��k�<,<i�߃=8]��Or�<}F���������9�P�ռ\<i}�;r].<t�;��=`��>��>8V�>��=��}�->[�ub���4>n#��j�\��]�dZ���F�1p��%%S>H�>��<p����
�>�bn>�n>P��?w�U?(>r���ݾ҄�������#%�=< }�<���:g3��mJ�k,?����v��>4R�>���>kd>��,���<�=@�����9��%?��L�CO&�X��MV��g��L���O���>ܸR?z���w��=)(�?RL`?�?�>�>a���Q���`=�m=�6��C:0�:������=�?3,�>/x�>߾V_�;H̾ ���߷>;I�N�O�j�l�0�����ͷ�>����/�о�$3��g��n���^�B�9Mr���>H�O?��?|7b��W���UO����*��q?�}g?��>wJ?�@?��y� r��F~�=
�n?C��?�<�?�>2=񮦽@	�>�?�ȏ?n�?l?��~�0~�>ۑ=��<>(Uu��Ȭ=W�3>h��=�.">��?�.�>p�>v²���9����e���qF�Z\=� �=�ל>�+�>n%m>��|='��=Ԇ>�l>�n�>l �>D|�>G��>�>�>�+��K�Y"?�>Ȱ�>��H?Hc�>Q��椽.�#>��<�|�mId�����<�H�x�����<��c=�j,=���>.r¿��?Oϊ>�		���?�(�\����>��>����ҷ>R�=>��T>_��>���>/�c=�'>�$>��Ҿ��>��L|"�PC���R���о��~>�<��-*��		�.��bI����އ���i�q���;=��`�<o�?���ٹk��)���C	?�Ҩ>�6?�ߎ��;���>}��>�Վ>�A��Q���'��FF⾏��?Q��?M&c>��>��W?��?�q1�!'3�KdZ���u�X)A�b�d���`��⍿����5�
�
��_?5�x?.dA?~��<�Yz>��? �%��돾|�>C/�5 ;�3�==�>�>� ��9�`�$�Ӿ�þW)�+�F>Z�o?��?�S?M`V�?���F�>�2J?.6<?`�d?�8?��4?�ZS�MS0?�.c>�q?�~?#2#?1�1?x�?B��>Fr�>�4�A�<䔨��X��Z1��4.��m��?�=�.�=l!�=�y�=Z��<rV�ɪ� �r=Ť�<����$3=/�=D�=��>�l�>�o]?@��>�v�>ע7?���38��$��g/?;=$����������p@>�k?h��?Q�Y?֭c>�$B��|C��>~G�>K�&>�G\>	 �>U<�5D�7�=�p>>�5�=2L��ށ�Ɏ	����,��<U0>"�?�7�>o��=J�=U���8~����&>d��˧S=�1��1�����>k�Ǹr>��T?ga>?<��=� ���;������v?lD?�_$?z~�?�RѼZ+�cj��S��̭��}?=�%�����4��Ⰶ�ǩ��&<�^>'W������)_>�����vl���H�
~���e=���D�=��
�zҾč}� ��=M�>�@��i~��ʖ��h��p�I?�́=&y��[�V�������>a��>��>�8�Tq��_>�S�����=av�>I@>�C�����ۢF�=w��K>�L? 2a?��r?�ό���m�"�K�E��[�������>^��>%K? >*��=瞠�0���?f��M����>�?�	��N�P�3���B��Q|3�`P�>Qh?�ݫ=���>7�X?�I?N?�m ?n��>�F>̺�
о�B&?�?��=��Խ��T�� 9�QF����>E�)?t�B�θ�>w�?��?��&?ՅQ?�?��>�� �gC@�F��>Y�>��W�:b��&�_>]�J?���>�<Y?�ԃ?�=>��5�M梾�ة��R�=k>W�2?�6#?��?ͭ�>���>ã���"�=���>� c?)3�?��o?�k�=��?��2>a��>��=&��>%��>� ?FO?��s?_�J?՜�>lI�<[i���󶽒Cr�U���~;�G<�B{=?2��t����r��<i��;䗻��Mh��D��(����;<��>BRu>�Y��5�>]�׾�]��8t>�d�<�^��u!���BP��؍=�&�>�?UI�>BC�z�m=|=�>N��>Z#�G@(?�V?��?�cD=��X��
Ҿ3�l�*ˡ>�W7?�ӊ=ʩd�����Wt�IO�=˞j?��K?�=����O�b?��]?@h��=��þ{�b����g�O?=�
?4�G���>��~?g�q?U��>�e�+:n�*��Db���j�#Ѷ=]r�>KX�R�d��?�>n�7?�N�>-�b>+%�=iu۾�w��q��g?��?�?���?+*>��n�Z4��I��y���$�a?���>s桾a�(?��&<r�پ�����j�2r��᧾Y���s���s���(�X�~��ֽ:��=��?�Sm?�j?�\?�#� g�ؾ\�Dkp���M�E|�W�@�H��x>���D�v�i�d��R�HǊ�Yw=�	��%U�
�?9�3?#���(?���ü�������>T�ʾ�Oi�,o'>���|E�;f	>`�9�X��Jc'�T�+?*�?�J�>-d'?E f�o�`�;X��a�zS㾛��=��#>G�P>bq�>#,==.�.͏��L��DL6�!܃�r�u>w�c?q�K?q�n?2t�?M1�����!�<�2��r����B>q_>.�>�V��0�&�"_>��r����"O����	��!=��2?"1�>���>�O�?��?�w	�}Ʈ�j�w��1��y<�%�>��h?��>�>��н�� ����>��l?���>��>ؖ��gZ!���{��ʽV&�>�>��>��o>�,��#\��j��L����9��u�=)�h?
���a�`�[�>�R?��:�G<�|�>~�v���!������'��>X|?;��=��;>,�ž�$�x�{��7��H>+?��?������#���>y?���>�˟>���?W�>�už�p+���?Hc?�K?F�??���>�~H=�_��@Tɽ:H*�C�J=�M�>B�T>BjO=�'�=����O�,;�J�m=��=W���Ǣ�~�<�S����u<��=hm1>��ڿ��K�.=۾ǹ����F�
�_�4�������_X��F���f����}���@�9��?O��\��X����p�/,�?7��?�Α�e���陿�~�]W�����>ڿr��ow�Tͱ����Ց�!"�`�������EM��j���e���?�耾uu¿����Y��a$?��>H^�?��'��&�]g���l=�c�<W
=�xt�PX��Mʿ?�5���Q?�%�>�����J��P_�>�Q">�U+>�A�>��S�G& �t�%>̈́?��?�c�>5��D��+iʿ��=���?=@�}O?Ix��׾R�=�p�>m�?i�>	9��7
�E�оE�>�è? ��?�~��3d��S/=�gz?U�=G I��:�L�>4�S=(�<� ��c�>:T>�!��"ƽkz��gE�=�ӕ>r��<׈>�Ŵ���m=��i>ڰ$�L�5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�����{���&V�}��=[��>c�>,������O��I��U��={~����ƿ�85�d%�4���B��얼�io�B����f���>��8������*>��<��>�R�>�$C>ց�=�D?��l?���>��ҽ��
�LJ��sn��ِ�矼�!��(VC�zqh������o־?9�e5����O��᪽�^b��"��x�2��R��f(�q#?��/>�Ҿ�8���=*��4�����9��|�=1i4�?n;�W�� �?i�??�Ge��0d��žR��=�>�5??ob8�
������r�=��=&+ ��|�>t�=�?۾�1��jK�w�0?`S?枾��現�(,>� �V�
=�5+??J2^<��>F�$?9�)���߽�Z>4>��>!#�>�'
>S䮾*ܽ0�?~�T?�z��Y�����>ƽ��qx�r�e=B>�5��S��.^>�q�<����Pp�bގ�}��<�:X?�ȍ>��(�n��q������0=��w?*,?V(�>ak?>IE?a'�<s�����T���� �=�X?�f?W�>8nv���Ͼ0ɦ���6?-,f?P�H>H s�|�8-�h��R?{�n?�? 7򼂞{�����&��>6?'�v?�a^�Oh������V�F5�>1E�>���>�9�v5�>�>?�"�6=�������_4�T?��@ϊ�?�'8<�뵎=�*?�H�>O3O�ƾn��򳵾�r=�>򚧾�=v�y��5�,�o_8?���?���>ܞ�����)ԃ=�����?�Q�?C}��E�=���d�s�������=9�<3�/�r�=�p羾V(��뫾��N|Ǿ����Ȩ�>&@��>�dը>�dN�m��i@տ�g�\������M�>�2�>�J��n��_Z��rv��xC�T�.�������>4%>i��=,���ڪ��%S�yӗ=��>ć��׫�>z��������/��<Ԣ�>�'�>�O>�M��%N�����?�3���ο��������O?2��?���?��?1���E���H�I��1����5?�o?�N?�I�=B�۽����qX?Q��Nc�b�@�5�I�#f>`jC?+�?~Z8�6|̺��=>�
�>�>Z�5W�������JϾߜ�?���?�Xؾn��>��?-%4?0b0�Č������2�"��0n>�$?�ý�^���l˾�_������!?��?<ބ��V�^�_?(�a�K�p���-�n�ƽ�ۡ>�0� f\��M�����Xe����@y����?L^�?h�?Ե�� #�g6%?�>e����8Ǿ��<���>�(�>*N>NH_���u>����:�	i	>���?�~�?Uj?���������U>�}?G��>R6�?$,�=���>���=�����I�!>��=7�;�L?��M?T��>��=d�7��.�LfF��R�9Z�nC�S�>"�a?oL?�mb>�y���90��:!�sϽ�/��5ۼ��@�'�0�<�ܽ�5>h>>�>�D��zҾ��?Mp�8�ؿ j��#p'��54?3��>�?����t�����;_?Tz�>�6��+���%���B�^��?�G�?<�?��׾R̼�>*�>�I�>��Խ����J�����7>%�B?Z��D��p�o�j�>���?	�@�ծ?hi�	?���P���`~�<��m7���=�7?m0�q�z>=��>(�=�nv������s����>�B�?�{�?c��>��l?e�o�w�B�!�1=3N�>��k?Ds?��o�+󾗰B>��?3������"L�f?��
@wu@p�^?~����ꚿ(ӾJ,�ln����<c >�Sɽp>n/U=��>	��b�����>XC,>yRq>�ps>F?�>��p>dQy�7���ÿm���	C��_7��r���!�g�޾��޾����[�������a=ܳ�v5ݻ�3��
����܄�[�=v)p?"�\?�$^?��>Q�0�!\�;rY��мx�#�~*�=T�>��5?��G?P;3?�Yw=�����_�����?����}�(v�>˃>��>���>r��>�ށ��G�=��>���>~U�=����k=䊄=��6>MG�>a�>(a�>�x�=�5<>����
��������w�� �?�����q���b��䙾������q<�<?�-m>�}��,�ʿ2��"�>?j>�����O԰�_�B>�O2?��>?��>�~־���<WՀ>G*Y��s���/>0^�=����T&/�M��>�A?Dhf>Z�t>�3�x8�P�P�Nw��6	|>r36?ض�+�9��u�a�H��Qݾ��L>���>	6?��_�Y����!�1/i��^|=�[:?wt?�m������Ʒu�%!���:R>R�[>�="�=uqM>�b��ƽ��G��6,=�s�=��^>�u?��+>ah�=��>��wpP��C�>�OB>�K->�??�$?�[�k	������g�-�?�v>'D�>�j�>>�hJ�F��=c��>Wb>n�b����8���?�uX>6�|�ц_�A�t���u=qH��g�=���=ґ �'<��8%=�~?���(䈿��e���lD?S+?b �=
�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��N��=}�>
׫>�ξ�L��?��Ž5Ǣ�ɔ	�0)#�jS�?��?��/�Zʋ�<l�~6>�^%?��Ӿ4g�>h���Z��F���u��#=[��>�@H?�q���O�ۻ=��i
?�?�P�գ����ȿ�rv����>��?�?��m��5���@�U�>���?�rY?�Ti>�A۾�aZ�`�>�@?
R?��>cF�{'�F�?5ն??JR%>1��?$�t?��>�Ʀ�)�8�|%��|����o=�)�@>O�s>C����M?�.���@����e�b���=�=�Cb=��>諢��Qľ�#�=�D��FW�����Ɠ�>�}�>�Av>�>�>U �>�J�>�&�>	v�<�-ܽ��J�"���N�K?���?����2n��M�<e��=&�^�`&?YI4?�b[�m�Ͼ֨>�\?Z?�[?�c�>P��>>��@迿�}�����<��K>G4�>�H�>�$���FK>�ԾX5D��p�>aЗ>�����?ھs,��fE��BB�>le!?x��>;Ӯ=�� ?5�#?�j>P9�>+hE��7��S�E����>��>mP?��~?Z�?i���IX3�����ࡿ'�[��7N>(�x?�]?�ϕ>ǎ������ΔI�NJ��Ғ�ҡ�?�mg?:��� ?�(�?}�??B�A?�Gf>Zv�A ؾɰ���Ԁ>P�!?6,���A��k&����|?�1?=�>"i��RFֽ ʼ���̔��S�?�2\?��%?����`��t¾���<�A'���U�Q�;�8L�P�>(4>�爽�˳=�>�G�=�Bm��\5�de< ��=�>�K�=�W7�/ь��=,?ٲG�ۃ�/�=��r��wD�>�>�IL>B����^?k=�h�{�;���x���U��?(��?Tk�?���ڝh��$=?��?�?�#�>OI��|~޾����Mw��|x��w���>`��>�l����n����F����Ž�a�>��>��>��?�ކ>)?Cc��7P��k���#�Y�(�Q��`��6!��?�1��)cD���>V���Eھ7-�>Gy�=N\�>��?{��>�i=��>%�]>4$�>T�~>Ͳs>s0N>�<>Xt>7�>��'�+�%��ZM?!k����&�Fw��Ǿ]4?��j?�?�>�!��4ჿ�y���?�~�?��?�U>G l�V�%�#�?��?����?���=R=)
�<`ɶ��9��;���J�k+~>��32���N���a�^
?A#?��D�]^���^�������s=1J�?
�(?��)��CQ�Cko��W���R�����k��C��o�#�(p�̔�������ك�%�(�l�%=Ќ*?.[�?���G[��ϭ�_�k�|�?��.i>��>�k�>Ǝ�>��K>�		�c1�ia]��Y'�J3��ϕ�>�z?�[�>��E?�D<?J�V?GP?�0~>w�>�ְ��d	?U"�<ۓ>���>O�0?�:?R
4?��?#(?��~>g(Ž`���)�ؾ�?sM?��?m��>�?^�~�����Wx	<��Q<�b���l4�=-�:=������ �=��Q>
�?�.��;I�����{>�f0?T�>?~t㾠r}���}>xۨ>g��>R>�5þ닿��d��>�ȉ?�b��}��d4;>Ѝ�=�����"���s>9L��n��=n�ȃ��q�y�>�8=��W���g�,�>TJ�i��=2u�>3�?���>�C�>l@��� �b���e�=�Y>�S>z>�Eپ�}���$����g�"^y>�w�?�z�?9�f=��=��=�|��cU����������<ˣ?FJ#? XT?H��?i�=?Wj#?Ե>+�\M���^�������?��+?0~�>����ʾ��3���?�?o a�^�:4)���¾ �ҽ�->:H/�,@~��毿´C��W�Q���N��;��?Y��?�a=�
�6�A�]���=T��\OC?/{�>�.�>��>K�)���g�&���:>A~�>{�Q?��>n�}?-Ղ?�E?�h>�9J�q��������̽)�>q�.?6��?䮇?x�s?�4�>`�
>x�����R��=�"��i2.�	�l>f�T>#��>TH�>��N>��ؼ��=�8=Ln��2���>���>�w�>{y�>t�> T�=��g?�	�>���i;Ǿ��ؾ�+�����<��t?,tz?��>��">-MϾ t(�M��Tͭ>���?�;�?�A?x�����>��%�����u����=?��?�b�=�K����=�������>�4?6&�&!��_�D=v=�T:?5!K?�� ���ÿ�n�񗉾Є����ܼՓ�Fe�P�X���M��Ri=1󞾸����`��� |�q��iR{�:윾�򬾝ȓ����>QO�=���=DT�=BG=�˻c΂����=��s�����۔Q�Rg�:�ۼf��ǝH���)��Us���)=���˾��}?�AI?��+?��C?->y>�>�4���>�����?X�V>բN�����`O;�����1����ؾ��׾��c�2���]>%�I�Q�>�3>�=�G�<���=�2t=@f�=��Q��=L��=]��=C_�=�h�=��>rK>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��=��=j?b�:�J�J5L��]c�FN��j�#?�%�D	��`g>!��=��̾b�׾w*�;��>��&=�|�<z���>�T�<Ⱦ��=�=�>�R>ה=.���5��=#c�Zj>��>Qˋ=��;�i= �=�IͽN&&>q�>	?�>x�?-3?�~j?\��>��z�[�־�:¾�>�>�\�>�b1=\K*>,��>yv;?��@?�iI?n��>1V�=<��>��>N����g�i��LO���W=d��?�x�?f��>��=�P.���sr>�A�ؽ�?�7?��?�<�>�U����SY&���.�������>��+=/mr��PU������l������=�p�>)��>�>�Ty>��9>�N>k�>�>V5�<$n�=0ߌ��µ<��約=8�����<�{ż�u���e&���+������;���;��]<��;��
=bT�>.>�V�>���=�����א>�4f�+�S�q�:�ȾDA��g���q�w���3�����=���>��T�/4����>&-�>L~T>��?�wz?��>(��z��S����8���h��"!�B�O�G(���3���c�JUV��㶾�J�>�
�>��>��R>�P.���?���=�NȾ��2�  �>�Ș��\c��:��d��響z����e���=��C?�)��!-�=��?�J?46�?,g�>Y|������=.s|�U�h<hz�r���H�pv?u4"?AB�>Jl���@��˾龽mk�>-�D���P�_����0���0�X���8�>(3��� Ҿ�
2�.��v���Q�A�)�r���>�O?4�?5�_�CP���aO����9��td?�h?>��>!U?�?b������~��m�=&on?j�?���?k)>:��=���
1�>?�?���?Vg�?r�o?)O����>� �<dq>����m�=\�>WD�=*�=�
??�?�����W	���r��ɪf���<®�=.A�>���>'ok>���=H,=��=ȟW>hG�>���>�[>�>���>�^�>51�~�?j>��>��\?o��>�A����򽿳3>�a���O��~������~5ڽ<�ļR>����ӽ�� >
��>z�¿�#�?�}�>ԅ�_*?U�����O�>�3>d���>v�>}G�>g8�>��?�`�>t��=$c�=)FӾ>f��Je!��+C�P�R�־Ѿ2�z>�����&�����z��DI��m���e��j�r.���;=�:ν<�G�?����r�k�L�)�C���	�?h\�>�6?
܌������>I��>
Ǎ>�I������ȍ�g���?1��?�<c>�>n�W?��?�1��3��sZ�i�u��&A��e��`�`፿G�����
������_?��x?xA?א�<�Cz>Ϣ�?��%�dԏ�� �>�!/�Y%;��<=]*�>;+��G�`��Ӿ��þ�4�oNF>C�o?$�?SX?TYV�x����N>JB?3�7?�4m?d�<?�=?��C�_�?�|>���>uc	?�d3?Vi,?z�?Z>2>�N�=g�漶r�=��)������������(���M	=� 4=N(>=-�B=�ž;�E-�(���6���?��9,j�v�;��v=خ>��>��#?#2D?r0?R?��_?�f�<�:���߾J�{?�f�=���	�˽�c��%�]�W�F��\?|}�?&5b?Jc�>]�L���M�95�>���>:3	>�N>��>��b���w�>��=w�<��c�<h%>G��@پh���P�4>�(�>�n�>�|>�`����%>�/���{��h>kWN��
��=�V�H�Z�1���t�IO�>�#K?�d?��=���=u����f���(?Ѽ<?58M?�a�?�{�=O(۾��:�b�K��y�s�>�t�<��
��ܢ��d���8:�)u8�,r>����٠�κO>V��RPݾ1h�bhK�ڲɾ��=z%��u��
��/���v����=���=A��N;�h������<?�<�=�ҕ��6��\��R��=mC�>��>_͉�����c�L��Ä���)<� �>%�u>O&���g��(HP��G�%/q>�79?�b?�?�?�U���i��C"�˫پ����dSG�iB�>\�P>�W�>X�X=���=:���[s���`��:��	?�?��ɴn�bھ��Vo$���?�M#?L�='�?��~?�?!$C?TD?��?��|>�䲽>���%K&?�?�y�=�eֽN�U���8� �E�o��>�)?�
D���>�?��?�g&?�Q?��?�>�� �lC@��C�>�>��W�n���$^>>�J?6��>{@Y?�܃?{+=>f�5��e��ˆ���f�=�� >3?6�"?e[?萸>̖�>Ei����>���>y�V?���?em?��=��?v�2>���>�K�=h�>;��>Z?�Y?�{�?��7?*�>,�a���Z�	�������;53�< �M=P�>O�Ē��C����2;�-4ǽ�<�Ń9���<$�P=���>u7W>������1>��ܾ#i�P�s>�1�"}��h�ky��'�=Wv>�+?ϔ�>�P ���=Ƽ�>ɶ�>�%���4?�@�>�?p݅=�Xj����'q6���>2Y*?��.>�(j��/��}U��^I�=K�t?��J?O����ܾ<�b?X�]?~d�#=��þ��b������O?z�
?��G��>:�~?��q?>��>��e��6n����Eb��j�w�=!p�>%Y���d��9�>e�7?)Q�>��b>�3�=4u۾��w��h�� ?*�?X�?2��?�(*>��n��2�R$��/N��f�Z?2��>?���ϱ&?��ü�;�ð������SӾ����f���n����l���6�;����+ֽI�=�?�m?��q?�2\?����]k�Zyh���y��aR�x��l���>��s8��W?�.�`�����ې�[�W=�]��B�C�)�?�*?�J����>)��(n �Sƾ�HO>������4���=�è��7�<HP�<��t��]*����	�?��>�F�>�e9?��[���H��>��4����>��>_�>��>����m�]��O�⾽�x�r����f>;b?��O? om?�p����6�"����#����c���P�6>b�>�@�>Z�2�f��O��i>���q�=
�Q#����؟;=k�8?�)�>��>r�?���>r��4墾�9w���-�����̃>}�R?Ĕ�>�x�>���<��L��>��l?��>��>����sX!��{�D�ʽ0�>�ޭ>b��>D�o>}�,�e#\�j��ۂ��?9�p�=J�h?�����`�I�>2R?%��:lH<	~�>v�K�!�x��N�'�6�>7y?�u�=�;>3~žT"�h�{�C7����T?��>`�E�%��q����D?�H?��>[n�?N�>O�3�^�9> 0/?.˂?�CV?�J<?�J?Z�=6f�'�̽2*T�6�ѽІ>�c>/n=ܑ=�D�0�V�"��뱘=n����.h��c����T����pM�=�Ԇ=�|/=���W�d�g|��p��D������ā���Nܼ�1��3:V��7h�{f���9��� /�p��<�P3�`{�z>T�%K���?A��?���pP��g���a��y�x��>�혾 �Ľ��T��q��qȋ����� ����$��jZ��	i���e���?��@�(+Ŀ����U����>}��>��?��1�"+'�u^��~��>�t��G%�7^�E����ѿ����J? d�>���¼��+6?��?z��>�=����������>n�D?�W�>6��>� 2�S�ƿ�y���>���?˥@�8B?�)�3��-�[=�f�>KH
?D�E>�"/�3�{���i�>�u�?�P�?H\=W�V��Z��oe?��<*�F��|���V�=���=B =���K>Yw�>��VY@��Wֽ|72>(�>p!&�Y��V%`��(�<B�`>&̽�F���Մ?]{\��f���/��U��\>��T?�*�>�H�=��,?�9H��{Ͽ��\�,a?Q0�?!��?�(?�ڿ��Ӛ>��ܾ��M?B6?e�>�a&���t�(e�=�2�C4��b�㾽"V����=ե�>�x>b�,����?�O��������=��%�Կ�8-������c>�3���pI���r�R���x�#���	��"��τ��(ڼr�D>�jo>_��>���>�h>ȿ�?�Xq?�L=%��=59��/f�?�;�=,����>����ǋ��Q�����S�ž �������ξ��.�4�=�Z��h��3�$�z�r��	"�U�?��8>����B����=����ǃ�0y`�2nK;!'����Q�%o��+ˋ?��>?U�\�U�p��	��)��ཱིnn?g�_�o��� 2>����{=��>Z8��+�no0�5�8�%^0?2�?EԾ��:����*>���N!=��+?T�?#�A<��>�$?�m+����2�\>5>P�>z��>�k>>��Ipܽ�?�sT?���;����E�>�྾�T}���b=�i>ID6���0�\>w��<ꀍ�EV��΍�ض�<�'W?N��>��)�&��N������3==�x?��?�1�>t{k?��B?(�<Gc��B�S��$�mw=��W?I.i?�>����Yо�w��*�5?�e?5�N>�fh����,�.��R��?��n?�Z?R����o}����\���r6?��v?s^�xs�����L�V�g=�>�[�>���>��9��k�>�>?�#��G�� ���{Y4�$Þ?��@���?��;<��X��=�;?k\�>�O��>ƾ�z������8�q=�"�>���~ev����R,�f�8?ݠ�?���>������k��=8����?%�?�J��E�<e��L�u�N�����O=��=Ҥڽ#b'�?꾮�4���Ͼ}��������=�ō>��@q������>��W����/8˿u�t�񷾾�:�(?�*�>�+.���|�� D�n``��}U�B�)���j���?��R>�
�=\���ξ�������[T>Hu%?��@>~)�=h�	�ES{>q�<�Jý?k�#?X��=�Ů��۾Ϗ�?��)�*���c�w��o3��}?�٫?|D?z�5?n�>�1�4�=�z�>TCl?��\?;r9?���=oi�<OT}���c?( ��L�]���5��u.�b�>�?!˫>��/�d��=˹p>��>ݘ>"a�ǿ$����J¾�?eQ�?����?�~�?'?P�6��񆿖����R�$�P=�-?lC>��˾��6��k���k<�d%�>t�?g _�U�0�F�_?ʚa���p���-��ƽzݡ>k�0�
b\��!�����$Ze�>���8y�j��?^�?V�?���� #�=5%?h�>񡕾	9Ǿ$>�<�~�>+�>f1N>OX_� �u>����:�7e	>��?�~�?�h?�������b^>t�}?w�>/�?|c�=�{�>�;�=���I2�	�">�T�=>�>�+�?�M?tG�>�]�=+�8�I/�OQF��=R�����C����>��a?��L?�tb>o���91��� ��Iν�1�n��@�.�)��x�4>�=>��>�D���Ҿ��?21 �39׿h�������7?kCg>3T?�J�e�U�4-<~(V?�0�>���A���9������<�?&��?�?+�;���;T�>D�>b��>C,����ҽ�B}��M>��;?� ��������s��3�>/1�?ۣ@��?��^��	?���P��Va~����7�c��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?Qo���i�B>��?"������L��f?�
@u@a�^?*�hֿ����dN��K���h��=���=��2>	�ٽ=_�=��7=��8�+<�����=k�>��d>3q>n(O>�a;>��)>���H�!�r��X���K�C�������Z�@��Xv�Rz��3�������?���3ý1y���Q�2&�_?`���=<�M?!Oe?!aj?�]�>�'��@�>� ���k=��1�ݡ�=�3>�&?��J?y�'?}zD>ή��vd�OCg�@�¾$���i�>�5�>�>���>-/�>����O�=b5�>�Γ>pLA>�Ӊ�ɖW�@	��}0>��>UV�>�B�>�>W�P>�5��0߾��cg�s�۾5o���"�?7^��nn�ۘ���8	��rѾ{��=a�4?�U�=h!����̿	>��f�:?6Ys�`��/+���
V>$�3?9?��> ����d����=`>�����Hp=�b<��wD��"�>�<?K_b>p�s>&z4��8�7�P��+���}>��4?J��s�B��et�. F�;�߾Q?M>\��>�˻/�|[��P!��ګg�6A�=n�9?Y�>q!��ȃ���ht�{q��ϾS>��U>���<X��=�G>!�X�(~���N�u�=P��=ZB[>�?/:+>}��=��>�<��aYP�)P�>��A>��+><�??�%?��<���Tl��n[.��w>�Y�>���>>�TJ��m�=[�>tPa>*+�
ʃ����D@��fW>��}���`�ar�1Bx=[��;��=��=�h �[>��X!=d��?D��ՠ��Z��O����F?>?7H�=zg�<ܓ�t���֫�*��?	�@��?I����Q���?E��?tڒ����=�'�>�>��̾4sB�œ?T�ѽw��3����*����?��?��ʼ=�����m���#>a�(?��׾�l�>����\������u��.$=N��>m>H?"]���aO���=��w
?]?�S�/����ȿ�|v����>�?��?��m��8��%�?�?t�>u��?YXY?�Ri>V^۾+$Z����>�@?R?`�>�K�s'���?o۶?��?�:>�B�?�sk?]�>���,�;�}���Ζ�����= l>ܜ>>`���H"�����8���怿�B��ɏ>�2@=�?*�*����xMn=*H�Pַ�j�d�k.�>҉�>m�]>;�>E�"?���>�ٓ>��K=��=U�R�iη�Q�K?*ʏ?� ��m����<���=��`���?�e4?2$b�jϾ���>��\?�?��Z?镔>�0�@��򋿿�������< J>_��>l0�>X�����K>6�Ծ?H�ݝ�>��>�F���ھ�(��i����=�>� ?���>�~�=(� ?G�#?�j>h,�>�ZE��8����E����>���>MJ?��~?7�?й�HV3�����䡿4�[�B=N>	�x?|T?���>R��������E�]�I����7��?Rug?K%��?�3�?�??ͥA?!9f>̃��ؾ����\�>�%!?��B���%����X�?�#?"6�>C֒��ڽ��˼N���X��V�?�2[?�u&?����a��ľM��<����Dvl���;��N�_Y>�V>E:��ZP�=��>�H�=q�i��5���q<���=E�>���=�c:��ᓽF=,?ҾG�@ۃ���=��r��wD���>IL>�����^?�l=���{�k��ax���U�� �?���?.k�?M����h��$=?�?@	?A#�>�K���~޾���Pw��~x��v�	�>w��>��l�<���������F����Ž�wl�R2�>o�>��1?#8!?f|>��>�\���U�`\��@ھKb�PF���G�s�Y���0��ф�,��1�&={�̾�W��b�F>wLؽ~M�>�o�>��>�ŉ>��>cĐ=��=�->���=LP8>#;�>�;>���=��g���ڽe?��پ	k�Jľ���{(M?�G?�_�>t��<+~b�A�&�)?���?x��?e�>��P���(��>4g�>H���_8?����WD��Z��=H3վ?�������㜼L/J>��:��A��q]�p9���<?Q�?���ؗ��$f������	cv=��?�d)?@p$���O�ݺp��<Z�3�Q����-]��5���V!�BJl�/)���]���*��L�#���f=�(?�m�?���Pv��㬾@r��^@��d>o�>�c�>�B�>��a>l��M)�@/T�%�(���R/�>uw?�Nm>��A?�fP?يJ?�C1?�]w>˃�>����j��>���e'�>�y�>�m? !?i�2?��%?%� ?���=3K)�}��YD���[,?�c#?��>"�?��>?Hо�`���=fFC=	w/��/�����=c���s���N�ݤ�=E�F>�1?����H1X��B��y�>�A?��m>Gp ?X�־\$�V�'>QN�>��?K&>��.�����F?�2�?�%�����x0�>�>?�/�po�=c�=���~O����:�����½8l>I!�-�R�	�>h�=�c�=�rR>�t�>5�?���>�C�>�@��-� �a���e�=�Y>;S>{>�Eپ�}���$��x�g��]y>�w�?�z�?�f=��=��=}���U�����F���2��<�??J#?'XT?_��?{�=?^j#?ɵ>+�iM���^�������?l!,?芑>�����ʾ�񨿍�3�ĝ?H[?�<a�3��i;)��¾��Խ��>�[/�q/~�����D��ʅ����y��(��?�?�A�C�6��x�ѿ��\��~�C?�!�>\X�>!�>��)�q�g�|%��1;>��>R?Gơ>V�?�(y?+�
?x�ۼ@t��/������G�>��>��?�@W?�?iߔ?��w>A|�<��6=F���������JF�_}��L'I��g�<���=�D�>�޵>3�==�����@ ��1�<���>
�>��>]1�>��]�����H?���>gֽ�����A��J���m���au?�Ő?WA,?L;�<[���C�����\��>�E�?Yɫ?T�)?,�U���=����4z��}�l��_�>qk�>٣�>{C�=H=V�>��>���>!�ϖ��8���`�u�?�F?���=ɕ��w�|��e�����4^��ٖk�ۧ��;�=�g�����	�=x]۾(���ʾ6�h��Jɽ�Af��iٽ#Qo���?ލ�=���=�D>w���߽*�=�=ѻ�8=FvS<f�q��--=
���"�=ʚo�1(>E�c=쬼�'��;�ʾ��y?�pK?�x0?��A?��y>�>c
m��>}���$�?��H>�n��V��zb:���D����ھH�־�[g�y١��q>����>�0>��=Mʜ<-�=ZҀ=�ts=�V߻�,�<�;�=2�=a�=@��=��
>��>�6w?X�������4Q��Z罥�:?�8�>f{�=��ƾq@?|�>>�2������xb��-?���?�T�?>�?Bti��d�>L���㎽�q�=H����=2>k��=w�2�T��>��J>���K��H����4�?��@��??�ዿТϿ7a/>��=L7��٘`���
�D�o��#��UI9�W5?�%���A�>�Ǽ���纾�F�I�>9g�=�W!��X��h�=n=��<^�f<:@p><��=|=>�.�+�=�,�<�����>if�=qT<eܪ��_�=���=o<hB�v��>ж?6�0?��d?O'�>+�l��Aξ���z��>���=���>�=�A>(t�>��7?��D?cL?���>w�=���>>��>�,���m�9V�{|��Q|�<��?�ކ?�.�>lA< �?�f����=��u½�v??,1?�[?F�>���>q'�3�-��럽�I�9{�=��l�z=a�W��)
��n��Y8�=��>M�>�b�>��x>j=>��L>5�>�>�=�<���=�1��k�<,<i�߃=8]��Or�<}F���������9�P�ռ\<i}�;r].<t�;��=`��>��>8V�>��=��}�->[�ub���4>n#��j�\��]�dZ���F�1p��%%S>H�>��<p����
�>�bn>�n>P��?w�U?(>r���ݾ҄�������#%�=< }�<���:g3��mJ�k,?����v��>4R�>���>kd>��,���<�=@�����9��%?��L�CO&�X��MV��g��L���O���>ܸR?z���w��=)(�?RL`?�?�>�>a���Q���`=�m=�6��C:0�:������=�?3,�>/x�>߾V_�;H̾ ���߷>;I�N�O�j�l�0�����ͷ�>����/�о�$3��g��n���^�B�9Mr���>H�O?��?|7b��W���UO����*��q?�}g?��>wJ?�@?��y� r��F~�=
�n?C��?�<�?�>2=񮦽@	�>�?�ȏ?n�?l?��~�0~�>ۑ=��<>(Uu��Ȭ=W�3>h��=�.">��?�.�>p�>v²���9����e���qF�Z\=� �=�ל>�+�>n%m>��|='��=Ԇ>�l>�n�>l �>D|�>G��>�>�>�+��K�Y"?�>Ȱ�>��H?Hc�>Q��椽.�#>��<�|�mId�����<�H�x�����<��c=�j,=���>.r¿��?Oϊ>�		���?�(�\����>��>����ҷ>R�=>��T>_��>���>/�c=�'>�$>��Ҿ��>��L|"�PC���R���о��~>�<��-*��		�.��bI����އ���i�q���;=��`�<o�?���ٹk��)���C	?�Ҩ>�6?�ߎ��;���>}��>�Վ>�A��Q���'��FF⾏��?Q��?M&c>��>��W?��?�q1�!'3�KdZ���u�X)A�b�d���`��⍿����5�
�
��_?5�x?.dA?~��<�Yz>��? �%��돾|�>C/�5 ;�3�==�>�>� ��9�`�$�Ӿ�þW)�+�F>Z�o?��?�S?M`V�?���F�>�2J?.6<?`�d?�8?��4?�ZS�MS0?�.c>�q?�~?#2#?1�1?x�?B��>Fr�>�4�A�<䔨��X��Z1��4.��m��?�=�.�=l!�=�y�=Z��<rV�ɪ� �r=Ť�<����$3=/�=D�=��>�l�>�o]?@��>�v�>ע7?���38��$��g/?;=$����������p@>�k?h��?Q�Y?֭c>�$B��|C��>~G�>K�&>�G\>	 �>U<�5D�7�=�p>>�5�=2L��ށ�Ɏ	����,��<U0>"�?�7�>o��=J�=U���8~����&>d��˧S=�1��1�����>k�Ǹr>��T?ga>?<��=� ���;������v?lD?�_$?z~�?�RѼZ+�cj��S��̭��}?=�%�����4��Ⰶ�ǩ��&<�^>'W������)_>�����vl���H�
~���e=���D�=��
�zҾč}� ��=M�>�@��i~��ʖ��h��p�I?�́=&y��[�V�������>a��>��>�8�Tq��_>�S�����=av�>I@>�C�����ۢF�=w��K>�L? 2a?��r?�ό���m�"�K�E��[�������>^��>%K? >*��=瞠�0���?f��M����>�?�	��N�P�3���B��Q|3�`P�>Qh?�ݫ=���>7�X?�I?N?�m ?n��>�F>̺�
о�B&?�?��=��Խ��T�� 9�QF����>E�)?t�B�θ�>w�?��?��&?ՅQ?�?��>�� �gC@�F��>Y�>��W�:b��&�_>]�J?���>�<Y?�ԃ?�=>��5�M梾�ة��R�=k>W�2?�6#?��?ͭ�>���>ã���"�=���>� c?)3�?��o?�k�=��?��2>a��>��=&��>%��>� ?FO?��s?_�J?՜�>lI�<[i���󶽒Cr�U���~;�G<�B{=?2��t����r��<i��;䗻��Mh��D��(����;<��>BRu>�Y��5�>]�׾�]��8t>�d�<�^��u!���BP��؍=�&�>�?UI�>BC�z�m=|=�>N��>Z#�G@(?�V?��?�cD=��X��
Ҿ3�l�*ˡ>�W7?�ӊ=ʩd�����Wt�IO�=˞j?��K?�=����O�b?��]?@h��=��þ{�b����g�O?=�
?4�G���>��~?g�q?U��>�e�+:n�*��Db���j�#Ѷ=]r�>KX�R�d��?�>n�7?�N�>-�b>+%�=iu۾�w��q��g?��?�?���?+*>��n�Z4��I��y���$�a?���>s桾a�(?��&<r�پ�����j�2r��᧾Y���s���s���(�X�~��ֽ:��=��?�Sm?�j?�\?�#� g�ؾ\�Dkp���M�E|�W�@�H��x>���D�v�i�d��R�HǊ�Yw=�	��%U�
�?9�3?#���(?���ü�������>T�ʾ�Oi�,o'>���|E�;f	>`�9�X��Jc'�T�+?*�?�J�>-d'?E f�o�`�;X��a�zS㾛��=��#>G�P>bq�>#,==.�.͏��L��DL6�!܃�r�u>w�c?q�K?q�n?2t�?M1�����!�<�2��r����B>q_>.�>�V��0�&�"_>��r����"O����	��!=��2?"1�>���>�O�?��?�w	�}Ʈ�j�w��1��y<�%�>��h?��>�>��н�� ����>��l?���>��>ؖ��gZ!���{��ʽV&�>�>��>��o>�,��#\��j��L����9��u�=)�h?
���a�`�[�>�R?��:�G<�|�>~�v���!������'��>X|?;��=��;>,�ž�$�x�{��7��H>+?��?������#���>y?���>�˟>���?W�>�už�p+���?Hc?�K?F�??���>�~H=�_��@Tɽ:H*�C�J=�M�>B�T>BjO=�'�=����O�,;�J�m=��=W���Ǣ�~�<�S����u<��=hm1>��ڿ��K�.=۾ǹ����F�
�_�4�������_X��F���f����}���@�9��?O��\��X����p�/,�?7��?�Α�e���陿�~�]W�����>ڿr��ow�Tͱ����Ց�!"�`�������EM��j���e���?�耾uu¿����Y��a$?��>H^�?��'��&�]g���l=�c�<W
=�xt�PX��Mʿ?�5���Q?�%�>�����J��P_�>�Q">�U+>�A�>��S�G& �t�%>̈́?��?�c�>5��D��+iʿ��=���?=@�}O?Ix��׾R�=�p�>m�?i�>	9��7
�E�оE�>�è? ��?�~��3d��S/=�gz?U�=G I��:�L�>4�S=(�<� ��c�>:T>�!��"ƽkz��gE�=�ӕ>r��<׈>�Ŵ���m=��i>ڰ$�L�5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�����{���&V�}��=[��>c�>,������O��I��U��={~����ƿ�85�d%�4���B��얼�io�B����f���>��8������*>��<��>�R�>�$C>ց�=�D?��l?���>��ҽ��
�LJ��sn��ِ�矼�!��(VC�zqh������o־?9�e5����O��᪽�^b��"��x�2��R��f(�q#?��/>�Ҿ�8���=*��4�����9��|�=1i4�?n;�W�� �?i�??�Ge��0d��žR��=�>�5??ob8�
������r�=��=&+ ��|�>t�=�?۾�1��jK�w�0?`S?枾��現�(,>� �V�
=�5+??J2^<��>F�$?9�)���߽�Z>4>��>!#�>�'
>S䮾*ܽ0�?~�T?�z��Y�����>ƽ��qx�r�e=B>�5��S��.^>�q�<����Pp�bގ�}��<�:X?�ȍ>��(�n��q������0=��w?*,?V(�>ak?>IE?a'�<s�����T���� �=�X?�f?W�>8nv���Ͼ0ɦ���6?-,f?P�H>H s�|�8-�h��R?{�n?�? 7򼂞{�����&��>6?'�v?�a^�Oh������V�F5�>1E�>���>�9�v5�>�>?�"�6=�������_4�T?��@ϊ�?�'8<�뵎=�*?�H�>O3O�ƾn��򳵾�r=�>򚧾�=v�y��5�,�o_8?���?���>ܞ�����)ԃ=�����?�Q�?C}��E�=���d�s�������=9�<3�/�r�=�p羾V(��뫾��N|Ǿ����Ȩ�>&@��>�dը>�dN�m��i@տ�g�\������M�>�2�>�J��n��_Z��rv��xC�T�.�������>4%>i��=,���ڪ��%S�yӗ=��>ć��׫�>z��������/��<Ԣ�>�'�>�O>�M��%N�����?�3���ο��������O?2��?���?��?1���E���H�I��1����5?�o?�N?�I�=B�۽����qX?Q��Nc�b�@�5�I�#f>`jC?+�?~Z8�6|̺��=>�
�>�>Z�5W�������JϾߜ�?���?�Xؾn��>��?-%4?0b0�Č������2�"��0n>�$?�ý�^���l˾�_������!?��?<ބ��V�^�_?(�a�K�p���-�n�ƽ�ۡ>�0� f\��M�����Xe����@y����?L^�?h�?Ե�� #�g6%?�>e����8Ǿ��<���>�(�>*N>NH_���u>����:�	i	>���?�~�?Uj?���������U>�}?G��>R6�?$,�=���>���=�����I�!>��=7�;�L?��M?T��>��=d�7��.�LfF��R�9Z�nC�S�>"�a?oL?�mb>�y���90��:!�sϽ�/��5ۼ��@�'�0�<�ܽ�5>h>>�>�D��zҾ��?Mp�8�ؿ j��#p'��54?3��>�?����t�����;_?Tz�>�6��+���%���B�^��?�G�?<�?��׾R̼�>*�>�I�>��Խ����J�����7>%�B?Z��D��p�o�j�>���?	�@�ծ?hi�	?���P���`~�<��m7���=�7?m0�q�z>=��>(�=�nv������s����>�B�?�{�?c��>��l?e�o�w�B�!�1=3N�>��k?Ds?��o�+󾗰B>��?3������"L�f?��
@wu@p�^?~����ꚿ(ӾJ,�ln����<c >�Sɽp>n/U=��>	��b�����>XC,>yRq>�ps>F?�>��p>dQy�7���ÿm���	C��_7��r���!�g�޾��޾����[�������a=ܳ�v5ݻ�3��
����܄�[�=v)p?"�\?�$^?��>Q�0�!\�;rY��мx�#�~*�=T�>��5?��G?P;3?�Yw=�����_�����?����}�(v�>˃>��>���>r��>�ށ��G�=��>���>~U�=����k=䊄=��6>MG�>a�>(a�>�x�=�5<>����
��������w�� �?�����q���b��䙾������q<�<?�-m>�}��,�ʿ2��"�>?j>�����O԰�_�B>�O2?��>?��>�~־���<WՀ>G*Y��s���/>0^�=����T&/�M��>�A?Dhf>Z�t>�3�x8�P�P�Nw��6	|>r36?ض�+�9��u�a�H��Qݾ��L>���>	6?��_�Y����!�1/i��^|=�[:?wt?�m������Ʒu�%!���:R>R�[>�="�=uqM>�b��ƽ��G��6,=�s�=��^>�u?��+>ah�=��>��wpP��C�>�OB>�K->�??�$?�[�k	������g�-�?�v>'D�>�j�>>�hJ�F��=c��>Wb>n�b����8���?�uX>6�|�ц_�A�t���u=qH��g�=���=ґ �'<��8%=�~?���(䈿��e���lD?S+?b �=
�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��N��=}�>
׫>�ξ�L��?��Ž5Ǣ�ɔ	�0)#�jS�?��?��/�Zʋ�<l�~6>�^%?��Ӿ4g�>h���Z��F���u��#=[��>�@H?�q���O�ۻ=��i
?�?�P�գ����ȿ�rv����>��?�?��m��5���@�U�>���?�rY?�Ti>�A۾�aZ�`�>�@?
R?��>cF�{'�F�?5ն??JR%>1��?$�t?��>�Ʀ�)�8�|%��|����o=�)�@>O�s>C����M?�.���@����e�b���=�=�Cb=��>諢��Qľ�#�=�D��FW�����Ɠ�>�}�>�Av>�>�>U �>�J�>�&�>	v�<�-ܽ��J�"���N�K?���?����2n��M�<e��=&�^�`&?YI4?�b[�m�Ͼ֨>�\?Z?�[?�c�>P��>>��@迿�}�����<��K>G4�>�H�>�$���FK>�ԾX5D��p�>aЗ>�����?ھs,��fE��BB�>le!?x��>;Ӯ=�� ?5�#?�j>P9�>+hE��7��S�E����>��>mP?��~?Z�?i���IX3�����ࡿ'�[��7N>(�x?�]?�ϕ>ǎ������ΔI�NJ��Ғ�ҡ�?�mg?:��� ?�(�?}�??B�A?�Gf>Zv�A ؾɰ���Ԁ>P�!?6,���A��k&����|?�1?=�>"i��RFֽ ʼ���̔��S�?�2\?��%?����`��t¾���<�A'���U�Q�;�8L�P�>(4>�爽�˳=�>�G�=�Bm��\5�de< ��=�>�K�=�W7�/ь��=,?ٲG�ۃ�/�=��r��wD�>�>�IL>B����^?k=�h�{�;���x���U��?(��?Tk�?���ڝh��$=?��?�?�#�>OI��|~޾����Mw��|x��w���>`��>�l����n����F����Ž�a�>��>��>��?�ކ>)?Cc��7P��k���#�Y�(�Q��`��6!��?�1��)cD���>V���Eھ7-�>Gy�=N\�>��?{��>�i=��>%�]>4$�>T�~>Ͳs>s0N>�<>Xt>7�>��'�+�%��ZM?!k����&�Fw��Ǿ]4?��j?�?�>�!��4ჿ�y���?�~�?��?�U>G l�V�%�#�?��?����?���=R=)
�<`ɶ��9��;���J�k+~>��32���N���a�^
?A#?��D�]^���^�������s=1J�?
�(?��)��CQ�Cko��W���R�����k��C��o�#�(p�̔�������ك�%�(�l�%=Ќ*?.[�?���G[��ϭ�_�k�|�?��.i>��>�k�>Ǝ�>��K>�		�c1�ia]��Y'�J3��ϕ�>�z?�[�>��E?�D<?J�V?GP?�0~>w�>�ְ��d	?U"�<ۓ>���>O�0?�:?R
4?��?#(?��~>g(Ž`���)�ؾ�?sM?��?m��>�?^�~�����Wx	<��Q<�b���l4�=-�:=������ �=��Q>
�?�.��;I�����{>�f0?T�>?~t㾠r}���}>xۨ>g��>R>�5þ닿��d��>�ȉ?�b��}��d4;>Ѝ�=�����"���s>9L��n��=n�ȃ��q�y�>�8=��W���g�,�>TJ�i��=2u�>3�?���>�C�>l@��� �b���e�=�Y>�S>z>�Eپ�}���$����g�"^y>�w�?�z�?9�f=��=��=�|��cU����������<ˣ?FJ#? XT?H��?i�=?Wj#?Ե>+�\M���^�������?��+?0~�>����ʾ��3���?�?o a�^�:4)���¾ �ҽ�->:H/�,@~��毿´C��W�Q���N��;��?Y��?�a=�
�6�A�]���=T��\OC?/{�>�.�>��>K�)���g�&���:>A~�>{�Q?��>n�}?-Ղ?�E?�h>�9J�q��������̽)�>q�.?6��?䮇?x�s?�4�>`�
>x�����R��=�"��i2.�	�l>f�T>#��>TH�>��N>��ؼ��=�8=Ln��2���>���>�w�>{y�>t�> T�=��g?�	�>���i;Ǿ��ؾ�+�����<��t?,tz?��>��">-MϾ t(�M��Tͭ>���?�;�?�A?x�����>��%�����u����=?��?�b�=�K����=�������>�4?6&�&!��_�D=v=�T:?5!K?�� ���ÿ�n�񗉾Є����ܼՓ�Fe�P�X���M��Ri=1󞾸����`��� |�q��iR{�:윾�򬾝ȓ����>QO�=���=DT�=BG=�˻c΂����=��s�����۔Q�Rg�:�ۼf��ǝH���)��Us���)=���˾��}?�AI?��+?��C?->y>�>�4���>�����?X�V>բN�����`O;�����1����ؾ��׾��c�2���]>%�I�Q�>�3>�=�G�<���=�2t=@f�=��Q��=L��=]��=C_�=�h�=��>rK>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��=��=j?b�:�J�J5L��]c�FN��j�#?�%�D	��`g>!��=��̾b�׾w*�;��>��&=�|�<z���>�T�<Ⱦ��=�=�>�R>ה=.���5��=#c�Zj>��>Qˋ=��;�i= �=�IͽN&&>q�>	?�>x�?-3?�~j?\��>��z�[�־�:¾�>�>�\�>�b1=\K*>,��>yv;?��@?�iI?n��>1V�=<��>��>N����g�i��LO���W=d��?�x�?f��>��=�P.���sr>�A�ؽ�?�7?��?�<�>�U����SY&���.�������>��+=/mr��PU������l������=�p�>)��>�>�Ty>��9>�N>k�>�>V5�<$n�=0ߌ��µ<��約=8�����<�{ż�u���e&���+������;���;��]<��;��
=bT�>.>�V�>���=�����א>�4f�+�S�q�:�ȾDA��g���q�w���3�����=���>��T�/4����>&-�>L~T>��?�wz?��>(��z��S����8���h��"!�B�O�G(���3���c�JUV��㶾�J�>�
�>��>��R>�P.���?���=�NȾ��2�  �>�Ș��\c��:��d��響z����e���=��C?�)��!-�=��?�J?46�?,g�>Y|������=.s|�U�h<hz�r���H�pv?u4"?AB�>Jl���@��˾龽mk�>-�D���P�_����0���0�X���8�>(3��� Ҿ�
2�.��v���Q�A�)�r���>�O?4�?5�_�CP���aO����9��td?�h?>��>!U?�?b������~��m�=&on?j�?���?k)>:��=���
1�>?�?���?Vg�?r�o?)O����>� �<dq>����m�=\�>WD�=*�=�
??�?�����W	���r��ɪf���<®�=.A�>���>'ok>���=H,=��=ȟW>hG�>���>�[>�>���>�^�>51�~�?j>��>��\?o��>�A����򽿳3>�a���O��~������~5ڽ<�ļR>����ӽ�� >
��>z�¿�#�?�}�>ԅ�_*?U�����O�>�3>d���>v�>}G�>g8�>��?�`�>t��=$c�=)FӾ>f��Je!��+C�P�R�־Ѿ2�z>�����&�����z��DI��m���e��j�r.���;=�:ν<�G�?����r�k�L�)�C���	�?h\�>�6?
܌������>I��>
Ǎ>�I������ȍ�g���?1��?�<c>�>n�W?��?�1��3��sZ�i�u��&A��e��`�`፿G�����
������_?��x?xA?א�<�Cz>Ϣ�?��%�dԏ�� �>�!/�Y%;��<=]*�>;+��G�`��Ӿ��þ�4�oNF>C�o?$�?SX?TYV�x����N>JB?3�7?�4m?d�<?�=?��C�_�?�|>���>uc	?�d3?Vi,?z�?Z>2>�N�=g�漶r�=��)������������(���M	=� 4=N(>=-�B=�ž;�E-�(���6���?��9,j�v�;��v=خ>��>��#?#2D?r0?R?��_?�f�<�:���߾J�{?�f�=���	�˽�c��%�]�W�F��\?|}�?&5b?Jc�>]�L���M�95�>���>:3	>�N>��>��b���w�>��=w�<��c�<h%>G��@پh���P�4>�(�>�n�>�|>�`����%>�/���{��h>kWN��
��=�V�H�Z�1���t�IO�>�#K?�d?��=���=u����f���(?Ѽ<?58M?�a�?�{�=O(۾��:�b�K��y�s�>�t�<��
��ܢ��d���8:�)u8�,r>���Y̨��V>��M�Ͼ��z�M1f�����=����Ɗ=�&�D�Ծ<�R�<��>�������w6��j㣿��H?�]r=�4�����(Ⱦ5W�=�>�>,ܐ>{6:�
-��%d��=��Y�=�L�>_�=-��� ���U��m�ꂈ>�;?�Bg?���?i�W�3#f�;���#�d����`;��?�Ip>R�?6�Y>q4>3n�����ut�b�b�>G�>��>���P�r�Ҿ�2߾�����>S�?WZ>۳�>wT[?�>5q^?u�?6�?hY�>8耼SQ���/?"=~?�x*>u#�����H�H�0��>{>?�����]>0j�>+C	?`�@?A
^?�})?�Ɍ>�� ��:V���>�l�>�Q���ǿ�Û=_i]?�>�)g?i��?���>��2�ぬ�R��'�>t��=�Sn?I�0?��2?r��>uK�>�ѾF�>>w�?�~?1�u?�? "�=���> ��=���>ܫ�=_��>��??y)?�=?��t?1�G?�o�>��U=ڥ�e[��E�W�]�q<0d����{;F=�Y��#�\�\����=�0>%t#>t���tн���/�߼kA�B��>qvs>bΕ�q!2>P�þK��� 4D>�u��&���拾<67�i�=S��>�� ?P��>a@%�ә�=�j�>�*�>���&m'?��?�?1l;F�a�{�ܾ��N���>s|B?���=�%l�PV��g(v��}=�n?@�]?N�X�������b?�^?�+�U!=���þ�b�.���O?��
?�sG�S�>(�~?& r?���>*ef��"n����cWb���j����=�P�>#=���d���>�|7?(�>@nc>D�=]۾�w�98��Q?m��?P
�?�?�o*>a�n�-���������b?���>����k7!?\ͼ�a׾�������l�ؾ���q-���C��+���X�����;����Y�=�k?ҭj?��v?p\?
�v�[�I�b��=���dU���,��['=�'�@�Od>�/o��J����X���E:=�k�z�P����?��+?�D]�M[�>����(��lӾ�g>�3���7D��ӽ����Z=��^=z����5½�-���$?{,�>�4�>�@0?�wi�!�$��F�L�B��s���)�=慛>`!�>���>?�N<	�}��t"����q�p�ȥ���le>^?�V?�J?�B���&�Ë���'��½ĩ��f�>��>(��>�ҽ/^ ��x�Gh$�����?��-�����s)>�f?cV7>��k>.��?�ݓ>��	��Ǻ� Z��Y�B�X��_#>�݄?���>���>:����=�1��>C�l?���>$h�>_���;!��|���̽�L�>�>��>��p>�+�u�[��q���i��`9�&��=f�h?�s��Ը`��ԅ>i�Q?�O�9�%C<VM�>rs���!����C'��o>/�?K�=��<>�Bž\�� �{�u����7?��-?�M����>��6�>�L?�o�>9L>��t?7�>��ھ%�޻��?��Z?�}I?]�Y?��!?�g}>��e���&�b�t=���>��s>������q>�(�]���E Ҿ�P�;��z>'f�>Z[�:9F�=��r� ���b���p>qӿ��N��E����ܲ��N��a&�i|�=��4�,њ��ǅ� ��쟾@�
���3=	2�������_�Wm�gG�?�h�?S�������6ב��|��S$�"=�>4n7<�P�hzǾ��_��|���-�2�=�o���+��N�WOX�A�8?�����˿�ȍ��y��1?�0?y;�?Ώ��<D��vH����>���=<=<��A��Q$ƿ�Bb���q?���>S	��9$�Ԙ�>vS�>��?@
G>Cl��Bjٽ�Z8��ve?��>��?�!��ƿ ���1,0=\�?f@�|A?��(�X��Y�U=y��>|�	?B�?>YW1�H�����@U�>s<�?B��?=�M=��W���	�5~e?�<#�F���ݻ��=�?�=�W=���$�J>�S�>Cz��WA��@ܽ߹4>�څ>'r"�У�w^�턾<��]>��ս�D��4Մ?�z\�uf���/��T���U>��T?�*�>%;�=Ų,?P7H�P}Ͽ��\��*a?�0�?��?H�(?�ڿ��ؚ>��ܾ{�M?ED6?��>�d&��t����=y7�^�������&V�u��=��>��>��,����O��G�����=�� �k�ſ~�)�-�9����h�@v������ý�!�ڲ��g�q�C'��ng=PC�=5Q>e�>�7L>:�O>.�Z?�$t?R;�>P@�=����,��44׾M4/=>I�������-�Ǧ����.h;�!����'��"!ƾ�Q:��|x=b�T�����5�/�x���=�ux1?�a,>�����Y�P��(׾�[�����<�񘽧���!�2���f��O�?�<?i�{���:��.�h ƽ'�ʽ"??�[T�~���~����;E>W"d��`���u>�jM�����n?��@���0?$�?Ǉ���쑾�+>.�����=1@+?֏?�x< T�>�%?�(�4��Xe\>�e5>@Ǥ>�J�>��>�����۽�b?��T?3�Ki��QH�>�=��;{�7 V=��>�u3�bjѼ�[>g�<+��Tun����[�<�)W?���>��)���9R����r�==y�x?�?GG�>�ok?��B?���<aY��3�S���5x=��W?�i?X�>�z��Kо�j��z�5?ʙe?�N>�dh�N���.�R��(?&�n?�_?�0���w}�������Im6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������P��=�㧾��?�ԅ?C����R=����;t��W �2S�<V��=朤���
��%��ׁ3��Ͽ�3��u⃾U�N��3�>�h@���}��>�~,��ֿ�O̿��v�E~��犾~q?G5�>��c�n���3�y� Ur��}N��E��!<��L�>6�>��������(�{��s;��X��a�>
�0�>��S�<#��'���1�5<)�>��>%��>�L��H뽾[ę?�^���>ο�������X?bg�?m�?�k?��9<��v�5y{����,G?�s?�Z?��%�&=]�7�R�n?�2im������3�m�9>��+?�w�>��%�����
�>n]?���>��#��)¿����?�+��?��?���?�t�?�7?�WԾR��-.u�����U��9�g?�>>�����f��_�ds�O�?�/L?^='�&�3�^�_?�a�G�p���-�<�ƽ�ۡ>��0�f\�M������Xe����@y����?F^�?h�?{��� #�Z6%?�>Z����8Ǿ��<���>�(�>)*N>�H_�j�u>����:�<i	>���?�~�?Oj?���������U>�}?�>"�?��=6��>0��=� ��*O�	�">��=g�=���?��M?w��>��=�9��.��2F��{R��
�C�J}�>��a?ѵL?42a>�蹽y|/�M� �tϽ�62���A�@���-��x߽��7>-t=>?>Q�D��mӾ��?����|ؿ[���(�X5?Z݃>�?�s��n|�6�ٻ�_?I\�>Z�K1��1���M���ի?z��?):?7־���X;>?T�>k�>9qѽ�������L,9>�oC?��yK��vso�i��>U�?�1@:��?��f��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?tQo���i�B>��?"������L��f?�
@u@a�^?*@�ۿ����eֳ��Kg�{j>%!=Z�{>0�u<�<�c��+�S=�m�<Gc7>Rm�>���>s|�>a�|>��<.p"</�����l,������~B�,�a|����kK���7l��� |���վ(���N��.׶�s�7��ؽ7��Q�=��M?��Z?J?`� ?���vI�=k��:�:0P%�`��= *>'*3?�]>?�/?C�r=�h��
8p��k�����-��/ܴ>Z,r>,��>b��>��>�IH�V�g> �k>�u">J��=R^�<�p=��-=�{o>堼>!^�>�Q�>��8>�>����Ov��� o�͘��`^˽��?uL����F�|���|������i=)8+?���=����<Oп�����J?.ʔ�r{�
/.�1R�=E[3?m	Y?�Q->tG��/���>Z����CX��>}�
�#!��gT.��M>�?�3>�
k>yP8�Ge6���Z�۾�R>,�>?d5���`n��N����X>���>&(<��dI���4z�ܐ>����=�7?9?u���wʾt_��r�����>9�N>*���Jl�=0V>>�V�����}�-#F����;z	A>�M?��+>�~�=&ף>`���QP�D��>�B>v,>�@?�%%?/%��͗������-��w>�Q�>�>9G>mTJ��ݯ=�t�>��a>�8���������?�m�W>�}���_�71u���x=�|���$�=�b�=U� �\=�&=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�<�>R=�JU��$΄���{�X��<�0�>|:L?ո��e���h�r�, ?��?]1뾍b���[ȿ��x�u��>���?�v�?~)n�L.���T=��+�>�
�?�W?	l>��ž�os�;f�>�i??bO?@j�>�) �>�C��[?��?���?��|>���?X�[?'�!=e�4>� ��:���2��� �>�v7�kճ>�Yv>Ϛ��NZ�����\�[��vx���+��P�>
.�<��>]6r��Ծ�F`>��A�^�&j����>)��>��V>d�>҈'?�?���>, U=�;a>��뾶Ѿ��K?���?����2n��a�<���=��^��$? I4?�'[���Ͼ�٨>��\?=?+[?c�>r���>���濿�}��3��<�K>g6�>RC�>�)��tFK>G�Ծc9D�&m�>�З>~�>ھ'*��<���@�>�d!?ϑ�>�î=p  ?]�#?}�o>�I�>*<D��1��܃G�@��>��>V�?*	~?�?;ݻ��4�f����8����\��L>��y?'�?_�>������x�HT��2�����?$h?�D�{�?È?�@?Б??"�Z>[��e�վ���:'�>e�!?Z�n�A��O&����?�N?=��>���8�ս�ּ�������?)\?D&?/��
*a��þH>�<�"�ӧW�E��;�#D��>�>2������=�>5а=aTm�T6���f<C_�=>��>��=['7�,o����+?��E�1&���,�=��r�N�D��~>�M>�q��V�^?�)>�t�{�����xn���/T�T�?-u�?/�?Y:��6Ih���<?�	�?�,?���>����)X޾���1�x�{wx������>��>�j��c�	���e����_��G�Ž?�h��Y�>�Ɂ>�?��?�S�=��?G]=,}_��+.�on��*�{� ���-�6=@��~'�xɒ������.ͽx幾�/���^�>��y��y>s?�Wp>�Xm>�?֊<҉�>'@>�<b>�Ɇ>륍>_�>AH�=C(�<[�H��OR?���Z�'�������	:B?\ld?h3�>�'i�J���/����?@��?Fn�?`�u>�h�t2+��y?f�>��n
?�:="���؉<�c�����=��CA����>Z�ֽ� :�QM�N{f��]
?�-?ȸ���d̾��ֽ�m|�H>F=���?$�?%v)�\�'�-�n�[��<�"�~�J$�O;���u=�C2z��u��3q��ȍ���	��>�?�ҙ?��$�	p�2k��B\��wE�?��>F�?��=>+��>P�u>\���-	5�����0"�p'���W�>��?_ҫ>i�C?Y�*?�QT?��n?l|�>�^�>������>��<Q��=���>shH?�j0?IW?�q@?AyR?S�>Y�ν�������,D?7<?=�?1�>v�>aO����L�{�<kV�=]Ҿr���X[�<�(>��
�kO>\�=߫>~!"?�%:�}�B��,����K>��A?K��>tu�>�Ռ�����EE=.��>�?���>�]�XR���i�8D�>N@�?:����=)�2>��=��`<)N���=��� �O=��{�#�=KA�դ�=iY.=��D�XR<��8<˯�=�2�=�t�>6�?���>�C�>�@��!� �l���e�=�Y>>S>>�Eپ�}���$��x�g��]y>�w�?�z�?i�f=��=U��=}���U�����H���s��<�??J#?XT?X��?y�=?gj#?��>+�fM���^�������?Y!,?튑>�����ʾ���3�Ý?u[?m<a�&���;)��¾&�Խg�>�[/�T/~����&D�X셻���-��#��?忝?GA�\�6��x�տ��\��c�C?�!�>,Y�>s�>`�)�y�g�y%��0;>���>ZR?"�>6�S?G&x?��H?k�d>��2��ٯ�����j��;�O1>�!@?�h�?�N�?$�s?�ڱ>��>�-��N��&񾯆2�ޞ��9g�Z�=�.>��>���>���>a�u=�j۽ī��l>"� j�=R��>^�?���>�O�>:�c>����U?uY?H����V��ۂ���=M�v��$4?X*�?�߂?xO׽<-�Pt��u��7�>�ҹ?�I�?�S?�����|�=���:%y��뉾?���>n��>���M��;4>��>ͩ�>���8�5�*�z��Y?�,B?}w(>�oſ��p���x�	���8T;�ڕ��c����rR��)�=�e��r�)٪���[��G��B��筲����z.}�$g ?B��=p�=�j�="�<jY�3a<��K=g��<|=�����a<<3:���N�����-�a��O<�m/=�-�u�˾VO}?��H?��+?��C?��x>c�>��-�=�>�R��24?�jS>^0Q�(E��X<�W���
��5�ؾm�׾I�c��ş� 5>&�H���>�W3>F��=���<��=eJs=jP�=�IG���=�^�=�=�ԭ=74�=~�>�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>s��=w�2�T��>��J>���K��A����4�?��@��??�ዿТϿ6a/>nr6>�%>ڿR�'=1���\��c��Y�"?�";��}̾Q1�>֌�=�߾	ƾ�b-=�5>:Bc=>�5\���=�y�	�>=<�n=�v�>��B>���=H&���e�=*TK=&4�=��O>�珻�{<��*�K�4=���=�Ta>��%>R��>l�?��0?6�d?)[�>��o�d�Ͼ�pþ���>Hr�=��>�l�=J}E>�r�>�_8?�LD?fsK?�h�>�Jf=���>C��>q-�u�o�m��@w��3�<8��?~�?�+�>T�5<	�:��R�Ư;�����O?�2?/	?�<�>�d��8쿎�$�1� ����4�:T�%>H�2�%j0��e ;p���ĽH�n=�	�>���>G$�>��>$�:> ��=��>:>����!��dƑ�=~�=`;�=�D�=u����>O��==̔��Q��@쪽�W���Kk�z����}=& >l��=�t�>�>�=D#�>�' >=�پ��]>nG&�7�k���:<y*r� �6�rO�%6��V5�;����$>\Xd>���P������>��>��s>ˣ�?-p?���>�O?�.���������$�^�޾'Rk�ߎ>�FW�� ��Q��U^��I��u�>A�>̟�>~�c>O=���K�Ȼ�=ȅ��G�?����>�Fj��==�!���D��(ՠ��1��ΘW�"��=�.H?�t���g>�}?HH?��?wx�>}@`����isl=�撾B�!=.2'������=?�e,?ϩ�>�����i��H̾,���޷>�@I�*�O���T�0���'ͷ���>������оl$3��g�������B�Mr�W��>%�O?��?,:b��W��KUO����w(���q?�|g?N�>�J?�@?�%���y�r���v�=�n?ó�?G=�?�>���=3᾽o��>E?�?h�?u?�x>����>�{;%&>�@�����=��>��=i�=1`?S�
?��	?�*���f
���M����Z����<�V�=�0�>M��>��g>Q��=�Gz=䍯=�}g>Sϝ>T�>k�X>nۢ>���>�ľ6Z��?��[>~�>�X?얔>���=�œ���2�=�˾󢫾s*��
��{�=a#Y���=���;���>��ÿ�ߥ?��>�k��~?��F��pپFЉ>��>'��ў�>�������=���>�>M�M���{>�B9>�r����>�'�8����j���x��f�����>��ܾ�%���X��U5=� H�-�Ǿ;�羱�m�����W�wi�;�D�?�@�#�w��P"��%���)?m�>�@?����w���$>on?��>Ѐ��\�����ܼ���V�?Q��?�;c>��>Z�W?�?�1��3�vZ�-�u�Y(A�e�1�`�፿���	�
�=���_?��x?yA?�T�</:z>Y��?�%�}ӏ��)�>�/�(';��@<=�+�>*��%�`�O�ӾL�þ8�&HF>t�o?,%�?QY?�SV���i�з>�n;?��4?��v?M�1?P�=?u��t_#?[(>{u?^�	?L6?��4?{�?�3>7B�= a};�z!=�ׇ�oϋ���ͽ�ʽ!zڼ��=V�-=ڗ亹�P;��<R|<U:���@%��v�<ӭʼ��|<�i&=�h�=p��=�
�>X�^?���>Zg>�8?'+��3�3/��5�1?�S�=Aᄾ~h��M����7�B:>�m?0�?v[?�V>�QA�	=� �>u4�>�")>�WX>g0�>5���Y�+�I=30>��$>���=UF��l~��B�VW����=�`%>���>�-|>�&��T�'>s����Kz���d>��Q�,ú�b�S���G���1��v��O�>��K?E�?~��=�_�@��9Df��.)?�\<?PM?�?��=w�۾+�9���J��>���>�̪<�������Z#��~�:��:K�s>�0��,{���U>ϵ��"ܾ�t�n�I���޾��V=h�	�@hD=w-�]�Ⱦqm����=��>`s��z�"����x]���O?�KE=�@��`�J�Ȇ��f�#>���>���>Fv2��ϖ�X�?�8d����=0x�>U�A>�:2�q����KM�S
���>p'M?\�B?���?B�h������K��侾�椾l`#��8?G�>sP�>fB�=��'>�y���
��q�r?G����>#��>W���Q���־5¾�^�:�_>�A)?�w�=$o�>`�H?�Y?jJ?��"?��?�6>t��[���T,?y��?\kS=�����M&��95�iH�=\�>�<_?Ei��%ύ>�?��.?��?�\S?��.?35
�ͿF�H�P���>EuG>�p�뷿�N�<x(m?'�>�Vj??b�?�>��n�����<7�>�+>�-P?9�>k��>Pe>���>ס���=Z��>Xnb?4b�?Rt?�Ξ=I��>�4>��>��=X�>-��>7?�RQ?<Jy?�SH?���>���<��ʽ�a��[AT�JTx��/5<w�<,]=S�9����*YҼa�=*z�:����������	=������t<,f�>�s>�I����0>Iži���s�@>>�������Tv��=9�u�=��>��?��>�$�I�=���>}��>�&��\(?r�?�?�d;��b���ھ��K�7]�>I�A?Se�=��l��}�u�eDj=��m?�y^?��X�W�����b?�^?���l\<�J%ľ�"f����uO?�p?�H���>Rm?��q?��>�g�M�m������b��k��ܵ=#P�>��4�c�.�>77?���>fe>	��=6�ܾ\Sw�T��Q�?^ی?��?O�?I�+>T�n���߿�5ܾ
^���,n?�+�>}�׾<�3?A&����z������"�۾DI��c�Ⱦח��Ѿ�!�qޤ�����>+>c{?��L?�5�?�L?�2�{�Y�5����&��1�N��氾G��9�K�� B�ܮ=��"�����_ �xnb�~��=��~�`�A����?h�'?1��1�>����s|�G;�kB>�t��w��i��=o����;=�
Z=��h�Q.�`���u- ?瀹>	-�>b�<?R�[�|>���1�	�7������4>hw�>_�>���>�v�:��.���轸�ɾ�p����ѽT�>d?��$?W�x?�­=$4e��̄���-e��q��Ң�>��>Ǜ>� G�(�&����ͪ��$o� ������p�d�ۼ�|8?��?��=>�u�?�� ?��7��T�� �:��7�kub���>E��?�(?��W>�~��*��]��>�
x?���>Ko�<{����ɾ+o����x&�>��)?���>�Z5��@n�-��9��ǳ���%D�#B�>�<|?��$�GJi���=��F?3-,���uí>���=� ؾF	־��E=���>/>?���=�>���v�þ�)w��<Ѿ�61?~?���;�,��Մ>�7*?���>�>�҈?�ʴ>fTʾ�����?�?V?��C?#M? ��>�:���+Cؽ�7�D�<5<�>;�M>1��<��>��U������Ľa��=���=�S�;s���en�2*>��=�N>��׿�iD�c�㾝���	�B����N�?���BQn����E˾��`��Z��Tc�Ueռ�O��bu��F���TE�}��?*��?H���7��>���p��*�u�>��]��/l��aǾ�2��!���"ݾF����D��X�r(v�;�i���;?���� ̿�l��i�����`?�?P�?&��� ��� ���>l�=a���վ|g��8[¿ ���a?��>�����	�(U�>���>� >Ѯg>�"`������dZ=Ra?�9?s�?�����ϿzԿ��;>4��?$�@'~A?��(�:�쾵�U=b��>J�	??�?>�G1�F�=����Q�>�;�?���?YM=��W���	���e?�<��F�|޻�=�L�=��=U���yJ>�\�>���[jA�I2ܽ��4>�ۅ>?l"����f�^�[G�<x�]>��ս-)��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�򉤻{���&V�}��=[��>c�>,������O��I��U��=dv��u���"4�̧O��UI��� �s>�1��|h���Ѿ� ������>��?ڳ�>P�>���= t�>�U_>FF?��M?&2�>K��=C� �ݝ��
�����=�G�<�0>�ٽ�yB=W���*���HCھ���Q��2A��5�_Gb<Cl\�k���	I��\�t�&��z ?�	=>B��\�i��3�=��0>��o=� ��'C�¢c��ި?f� ?{���o�<�K��t��=�$W��P?l�ӽ��������<�5,���=��>G��=��	���S���l��:6?��?И��Q�����O>�I���D;�?��>G0>�Q�>W�?>|V�[`>���>� ?z��>�L	�Z������I�%?!�Y?�5����̾�)�>=2ƾT0ؾ�4_=��9>�Cս�}���;?>ղ�=�茾�𠽤�Q<�i�<�%W?V��>��)����Q��X��l�<=2�x?]�?�3�>�sk?W�B?��<<k��X�S�� �
w=��W?8/i?ȶ>�U��"
о����ں5?��e?��N>y�h����/�.��O�n?�n?�a?,��j{}�������im6?��v?s^�xs�����N�V�e=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?��;< �X��=�;?l\�>��O��>ƾ�z������-�q=�"�>���ev����R,�f�8?ݠ�?���>������v��=���,�?�݆?2������<��IHj����[��<ޝk=����7޿�����B���ľʱ�З���t�<JI�>�5@i$ ����>�A�r*�>ҿv����ž��M�}?�S�>Y~'�����ށk��j�{�5���6�&3��4I�>h�>Z�� �����{��p;��^����>�����>��S�}������S�5<��>^��>��>򩯽��]Ǚ?Bb��>ο�������X?9_�?�m�?�p?&�7<��v�ަ{��\��*G?��s?:Z?`�%�&g]��s8�;Pm?d �Y�o�W��BJ��4>�I#?���>�-"��7W=!ߙ>Ǭ?��>&?�Ht��b����?���?8��-?�P�?n�%?��E��r�����E��B�I?ϰ�>[��udF�(1�LA���5%?9LB?T��9-�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�>��?,��=�%�>��=��c�]�(�#>0��=�B��R?`N?U��>�=u�8��/�T�E�TQR���ȇC�P��>a?�ZL?9�e>����-�0��: ��4ҽw�1�(�޼�j@���1�R߽7Z9>�?>��>X�F��HӾ��?T}�B�ؿ�d���'��<4?u��>�?=��7�t�&�)G_?��>�;��)�� +���Z����?mI�?�?R�׾<.˼�5>>ܭ>�>�Խ���2�����7>��B?�!�@���o����>���?�@P֮?��h��	?���P��Ua~����7�d��=��7?�0� �z>���>��=�nv�޻��X�s����>�B�?�{�?��> �l?��o�O�B���1=9M�>͜k?�s?}Qo���i�B>��?#������L��f?�
@u@`�^?*wٿ�0��v�Ǿ��ھ]��Z9�<,K�>�왽,���A�h�1��4c}���V>��>}�>���>��k>&4r>ʼ>/�|�����������,�D���JY ���.������YuE���վ�U����>�g�=fb�t
����4�0����=͛U?v�Q?Mp?%?=V����>1�����<Y�"�☊=+A�>��1?%)L?�*?��=�����d��Q��.7��>����=�>��H>���>���>v��>(�:�H>?>�^�>xK >� =4(F���=�(O>���>n �>q��>��d>�3=ӹ�4I��K��j���n��L��?.g�@�J��_��MF_��`���;�=G)?�>�S��Q�տn���-j[?��ž���Z��m?T>&*V?��;?*�~>�5��Jӻ��Ǎ>P�ܽ�Hݽ�ޖ=|�#�R����x���Y>��?��f>Ku>d�3��e8���P�{���g|>Y46?�涾�B9���u���H�cݾ�IM>?ž>��C��k�^�����ui�E�{=�w:?��?�5���᰾�u��C���OR>�;\>�W=Pi�=xWM>�gc�;�ƽ�H�w.=���=ܮ^>)g?�l,>mq�=c��>�����P�:h�>�B>�+>�L@?F#%? �����k��p�,��cx>�#�>%�>$�>3K��=i��>�c>Ь�7Q����
��@���U>aJ���^���u��w=	����=���=���[D<�V$=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�h�>Hz��Z��|��~�u���#=7��>�8H?�V��U�O�:>�Xw
??2_�ѩ����ȿ)|v����>g�?|��?�m�JA��I@�$��>Ģ�?sgY?�ni>�g۾�_Z�;��>��@?�R?��>-:�6�'���?߶?篅?��R>�G�?*Sj?��>��</���J��S����=Q]�=�b�>��<��о��A����z����h��o��>��*=��>�I��b�Ͼ��-=?�8)v�ʐ���>���>��Z>�Њ>Z?U�>�Z�>�.���� �4�a��Љ�V?�̎?���,r����=��&>���u,?:\?}<����<r>�J?�ă?�%^?�U�>�a�LW���з�V����;�>���>$��>-'$=Nq>������'�>6�j>pɼ
� ������A���>D�A?w�?�f>i�"?}�#?7)n>�9�>z�M�����{@�f�a>���>Ȟ#?�x�?��?�,ɾ~�*�r����ţ�I\�6�>Dn?ȁ?�2|>&���k�t��쑼O�k�V�}�4@�?�[]?��Ǿ��?�#�?�wV?v?�9H>(��;
}���N��z�=�"?�P�fA��q&�_����?ڴ?���>�A��@�ӽ ?����8C���)?.(\?h�&?~W�+a�P>þ�:�<�!'����&<�yB�Z>�">k4���=6<>��=�l��c6���P<��=+M�>q�=dg5�ԗ��$=,?2�G��ۃ���=u�r�TxD���>%JL>A����^?jk=���{�����x���	U�� �?��?Ik�?B��a�h��$=?�?H	?�"�>�J���}޾��}Qw�I~x��w�w�>m��>;�l�E�%��������F��
�Ž�k��s[�>�y>�x?D?�)$>��>3)t���T��>����L$e���)�ۀ@��9�I�*�Xؕ�F��.���,��I?��Ͷ>���yZ�>�k ?>��>X�4>���>�P���a3>��@>��t>�9�>2>�bl>A�Խh�<�̻�KR?����%�'����²��g3B?�qd?S1�>ui�;��������?���?Qs�?=v>h��,+��n?�>�>H��Vq
?�T:=Y8�;�<V��t��3��)�1��>�D׽� :��M�Dnf�sj
?�/?�����̾�;׽���Ln�:�D�?��*?�,���G���t��W�bMV��-���u�����2��rt������0~�P���s��	�=(�%?yV�?P�������{��m��-N��7C>���>s��>�۰>��->v��W+�zX���h[;���>�r?E�>��>?9`M?�5O?&:@?�t>��?�T��P�>A��>4��>��>�9?�g?�@?�:<?��`?0N\>�B¾���2j��'T:?H�1?�6?S��>�a&?�o�����=����Kg�/3m�6�
�uW�=��>gP�E���ywE=8�P>�Z?���{�8�H�����j>�7?�|�>���>���6/���<��>"�
?�8�>� ��r�ed�*Y�>Y��?����=W�)>��=.ԅ�M��{k�=�¼7�=�灼�;���<��=|�=Sh~�����kT�: 4�;�X�<���>X�'?�x�>��(>C���e,��F�c1:>��u>|��=��Ւ������ Bp���,>~!v?��?��i>���=�u>�Ǽ�����4�v/y�k�=�W�>L�*?��a?j��?�#?��<?m�N>���*\��#͈��`U�n�?�!,?���>�����ʾ�񨿦�3�ӝ?p[?�<a�9���;)���¾Q�Խq�>�[/�~/~����"D��ׅ����/��,��?뿝?�A�j�6��x�ҿ���[��s�C?'"�>Y�>��>N�)���g�v%�2;>1��>yR?i�>[�O?��y?}_\?�]>�Z:�$��������Bo���>&�A?s�?���? w?�O�>��> )��~�]���kN#�FC�A����Q=��]>Rؐ>���>|��>f�=��Ľ\c��#�?���=mD]>R��>nz�>�3�>��r>N�<�TT?�� ?V������g���_��a5�wI?ᴞ?��2?9�n�0��sF$��z����>��?���?�-?��}��=�/��'Ͻ�@���_�>�\�>5ؙ>LJ�<��=0o>:A�>bP�>�����"%��B�U�QQ?z�<?��<��ſ��h��c��,���7�!�N����M0�Y 0�+�8���=lř�0½�����T��ʢ���&�������OS�0�?���=ڏ�=	�>~D���Q=��<c.=�=�|ν��~=��d�2�?��̨����Y��(-�����,sɾO|?��D?!-?�zH?�8[>�>O*��>=���@?�XT>�H��u����e4�%��C����ݾIپNd_��ř�
k>�pm��g
>50/>A:�=��<���=�Do=m�x=M��;5Y!=Gȶ=ZT�=���=�*�=�C>:e>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>X�6>�w>]dR��y0���W��e���Z� �!?�{;�6#̾��>���=`�߾l�ƾ&�0=�4>�`=H��Z3\�Nm�=��v�|J;=2f=un�>*ZC>���=�I���T�=�]I=���=rP>:7���t;��%���9=�=�=W�a>~f%>ތ�>.�?�[0?[d?*Q�>�Dn�3$Ͼ�0��~8�>��=t_�>s�=�MB>Q��>�7?&�D?`�K?�k�>��=��>��>��,�g�m�od�#ɧ��T�<���?ˆ?0ϸ>BQ<܂A�/��ef>���Ľ$x?oH1?�e?#۞>���޿��&�#�0�lŬ�ѻ�L=Xj��LQ�!���aڽ:�=�7�>�|�>K9�>�&w>+�>>"�P>���>��>64�<J_�=ε�q;�<����r=Nd�D�
=d�
�?�;����m�9�:X��^��\Y9���<�?�;
�j=U�>F}8=�;�>���=��ξJX>�{B�f���y=�6���5��#m��u��;5��WR>�w)>q��ڗ��?��a>l%U>`�?�&v?�5�>H�1�`�������C������8��=�"5>U0��R*���H��I��A�a��>�"h>uB�>{�e>o\)��0H��]�=�뿾%8�}��>�~/��g:���C��x�Ӛ���d����X�Y��<�wG?泍��{7>�x?��A?��?�ٺ>�&^��lξ���=i���"<���_��@o��Z� ?�(?0��>c���\�H̾$h��?�>��H�r�O������0��Z"�z鷾L|�>F��AѾR3��i������zB�\r���>�O?iޮ?��`�b��lO�ǒ�۴���9?2[g?�7�>�@?T.?�?��ō�,a��ل�=��n?��?U:�?9><~�=Ę��S��>�	?p��?O��?��s?��A�4��>랢;5� >ȋ�����=��>�8�=�R�=R
?9x
?�A
?����&�	�rm�C�!^��S�<��=�>"��>�tq>u��=ah=R��=*\>쒞>�~�>��d>��>�S�>���؆��a?��P>�A�>O�'?dz�>��>%<�fj��uA�x�1�o?����D�	rD���ؼ����R�=f*9<�q�>܌ڿ��?O�*>�/�0(?r�*��:==�>��I>�b�~��>�2>�ap>���>�y�>��=��>M>u>33ӾRE>����h!��8C�{mR��Ѿ3�z><���K*&�q��_S��dHI�tb���Z���i��/���G=�v�<]H�?N��o�k�$�)��d���?�X�>6?Rڌ�S���>���>]Ѝ>7T��}����ȍ��Xᾗ�?>��?��w>h1�>^?P�?�@����;�1$z���k���=���G�%�W���:��)��Nk��2@?~U?��K?ls>��h>fŕ?��K�"��HB�>4#��D?�(f�<��>2���LI��ž���>�߽�_f>�J?�sz?h�/?.���ȽCK>y�?�̃?�Rw?��-?�cs?[R��N��>?�r>�g�>S�>٭V?�M?ރ4?��>��?�ݍ=����{Q���������}�<�$���Z=�e=G�ɽ>ʽ��]���B=m�?����BN�=#���4L�;�%P<�i�=�Z >�*�>�\??��>*�y>�6?���.�8��1��#/?"��=�P����������Z���>�l?���?ŃT?rG>�^F�,�F�F�!>���>��$>�r?>;d�>z�	��ep�1��=�y>�#>[͵=�hs�e��*	�ዊ���=d>��>2|>��ݴ'>d{��`,z�z�d>�Q��ɺ���S�!�G�n�1���v�_Y�>��K?l�?Q��=I_龓4���Hf�B/)?>]<?�NM?��?��=M�۾��9���J��;���>Zh�<��������#��r�:����:��s>2��,{���U>ϵ��"ܾ�t�n�I���޾��V=h�	�@hD=w-�]�Ⱦqm����=��>`s��z�"����x]���O?�KE=�@��`�J�Ȇ��f�#>���>���>Fv2��ϖ�X�?�8d����=0x�>U�A>�:2�q����KM�S
���>p'M?\�B?���?B�h������K��侾�椾l`#��8?G�>sP�>fB�=��'>�y���
��q�r?G����>#��>W���Q���־5¾�^�:�_>�A)?�w�=$o�>`�H?�Y?jJ?��"?��?�6>t��[���T,?y��?\kS=�����M&��95�iH�=\�>�<_?Ei��%ύ>�?��.?��?�\S?��.?35
�ͿF�H�P���>EuG>�p�뷿�N�<x(m?'�>�Vj??b�?�>��n�����<7�>�+>�-P?9�>k��>Pe>���>ס���=Z��>Xnb?4b�?Rt?�Ξ=I��>�4>��>��=X�>-��>7?�RQ?<Jy?�SH?���>���<��ʽ�a��[AT�JTx��/5<w�<,]=S�9����*YҼa�=*z�:����������	=������t<,f�>�s>�I����0>Iži���s�@>>�������Tv��=9�u�=��>��?��>�$�I�=���>}��>�&��\(?r�?�?�d;��b���ھ��K�7]�>I�A?Se�=��l��}�u�eDj=��m?�y^?��X�W�����b?�^?���l\<�J%ľ�"f����uO?�p?�H���>Rm?��q?��>�g�M�m������b��k��ܵ=#P�>��4�c�.�>77?���>fe>	��=6�ܾ\Sw�T��Q�?^ی?��?O�?I�+>T�n���߿�5ܾ
^���,n?�+�>}�׾<�3?A&����z������"�۾DI��c�Ⱦח��Ѿ�!�qޤ�����>+>c{?��L?�5�?�L?�2�{�Y�5����&��1�N��氾G��9�K�� B�ܮ=��"�����_ �xnb�~��=��~�`�A����?h�'?1��1�>����s|�G;�kB>�t��w��i��=o����;=�
Z=��h�Q.�`���u- ?瀹>	-�>b�<?R�[�|>���1�	�7������4>hw�>_�>���>�v�:��.���轸�ɾ�p����ѽT�>d?��$?W�x?�­=$4e��̄���-e��q��Ң�>��>Ǜ>� G�(�&����ͪ��$o� ������p�d�ۼ�|8?��?��=>�u�?�� ?��7��T�� �:��7�kub���>E��?�(?��W>�~��*��]��>�
x?���>Ko�<{����ɾ+o����x&�>��)?���>�Z5��@n�-��9��ǳ���%D�#B�>�<|?��$�GJi���=��F?3-,���uí>���=� ؾF	־��E=���>/>?���=�>���v�þ�)w��<Ѿ�61?~?���;�,��Մ>�7*?���>�>�҈?�ʴ>fTʾ�����?�?V?��C?#M? ��>�:���+Cؽ�7�D�<5<�>;�M>1��<��>��U������Ľa��=���=�S�;s���en�2*>��=�N>��׿�iD�c�㾝���	�B����N�?���BQn����E˾��`��Z��Tc�Ueռ�O��bu��F���TE�}��?*��?H���7��>���p��*�u�>��]��/l��aǾ�2��!���"ݾF����D��X�r(v�;�i���;?���� ̿�l��i�����`?�?P�?&��� ��� ���>l�=a���վ|g��8[¿ ���a?��>�����	�(U�>���>� >Ѯg>�"`������dZ=Ra?�9?s�?�����ϿzԿ��;>4��?$�@'~A?��(�:�쾵�U=b��>J�	??�?>�G1�F�=����Q�>�;�?���?YM=��W���	���e?�<��F�|޻�=�L�=��=U���yJ>�\�>���[jA�I2ܽ��4>�ۅ>?l"����f�^�[G�<x�]>��ս-)��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�򉤻{���&V�}��=[��>c�>,������O��I��U��=dv��u���"4�̧O��UI��� �s>�1��|h���Ѿ� ������>��?ڳ�>P�>���= t�>�U_>FF?��M?&2�>K��=C� �ݝ��
�����=�G�<�0>�ٽ�yB=W���*���HCھ���Q��2A��5�_Gb<Cl\�k���	I��\�t�&��z ?�	=>B��\�i��3�=��0>��o=� ��'C�¢c��ި?f� ?{���o�<�K��t��=�$W��P?l�ӽ��������<�5,���=��>G��=��	���S���l��:6?��?И��Q�����O>�I���D;�?��>G0>�Q�>W�?>|V�[`>���>� ?z��>�L	�Z������I�%?!�Y?�5����̾�)�>=2ƾT0ؾ�4_=��9>�Cս�}���;?>ղ�=�茾�𠽤�Q<�i�<�%W?V��>��)����Q��X��l�<=2�x?]�?�3�>�sk?W�B?��<<k��X�S�� �
w=��W?8/i?ȶ>�U��"
о����ں5?��e?��N>y�h����/�.��O�n?�n?�a?,��j{}�������im6?��v?s^�xs�����N�V�e=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?��;< �X��=�;?l\�>��O��>ƾ�z������-�q=�"�>���ev����R,�f�8?ݠ�?���>������v��=���,�?�݆?2������<��IHj����[��<ޝk=����7޿�����B���ľʱ�З���t�<JI�>�5@i$ ����>�A�r*�>ҿv����ž��M�}?�S�>Y~'�����ށk��j�{�5���6�&3��4I�>h�>Z�� �����{��p;��^����>�����>��S�}������S�5<��>^��>��>򩯽��]Ǚ?Bb��>ο�������X?9_�?�m�?�p?&�7<��v�ަ{��\��*G?��s?:Z?`�%�&g]��s8�;Pm?d �Y�o�W��BJ��4>�I#?���>�-"��7W=!ߙ>Ǭ?��>&?�Ht��b����?���?8��-?�P�?n�%?��E��r�����E��B�I?ϰ�>[��udF�(1�LA���5%?9LB?T��9-�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�>��?,��=�%�>��=��c�]�(�#>0��=�B��R?`N?U��>�=u�8��/�T�E�TQR���ȇC�P��>a?�ZL?9�e>����-�0��: ��4ҽw�1�(�޼�j@���1�R߽7Z9>�?>��>X�F��HӾ��?T}�B�ؿ�d���'��<4?u��>�?=��7�t�&�)G_?��>�;��)�� +���Z����?mI�?�?R�׾<.˼�5>>ܭ>�>�Խ���2�����7>��B?�!�@���o����>���?�@P֮?��h��	?���P��Ua~����7�d��=��7?�0� �z>���>��=�nv�޻��X�s����>�B�?�{�?��> �l?��o�O�B���1=9M�>͜k?�s?}Qo���i�B>��?#������L��f?�
@u@`�^?*wٿ�0��v�Ǿ��ھ]��Z9�<,K�>�왽,���A�h�1��4c}���V>��>}�>���>��k>&4r>ʼ>/�|�����������,�D���JY ���.������YuE���վ�U����>�g�=fb�t
����4�0����=͛U?v�Q?Mp?%?=V����>1�����<Y�"�☊=+A�>��1?%)L?�*?��=�����d��Q��.7��>����=�>��H>���>���>v��>(�:�H>?>�^�>xK >� =4(F���=�(O>���>n �>q��>��d>�3=ӹ�4I��K��j���n��L��?.g�@�J��_��MF_��`���;�=G)?�>�S��Q�տn���-j[?��ž���Z��m?T>&*V?��;?*�~>�5��Jӻ��Ǎ>P�ܽ�Hݽ�ޖ=|�#�R����x���Y>��?��f>Ku>d�3��e8���P�{���g|>Y46?�涾�B9���u���H�cݾ�IM>?ž>��C��k�^�����ui�E�{=�w:?��?�5���᰾�u��C���OR>�;\>�W=Pi�=xWM>�gc�;�ƽ�H�w.=���=ܮ^>)g?�l,>mq�=c��>�����P�:h�>�B>�+>�L@?F#%? �����k��p�,��cx>�#�>%�>$�>3K��=i��>�c>Ь�7Q����
��@���U>aJ���^���u��w=	����=���=���[D<�V$=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�h�>Hz��Z��|��~�u���#=7��>�8H?�V��U�O�:>�Xw
??2_�ѩ����ȿ)|v����>g�?|��?�m�JA��I@�$��>Ģ�?sgY?�ni>�g۾�_Z�;��>��@?�R?��>-:�6�'���?߶?篅?��R>�G�?*Sj?��>��</���J��S����=Q]�=�b�>��<��о��A����z����h��o��>��*=��>�I��b�Ͼ��-=?�8)v�ʐ���>���>��Z>�Њ>Z?U�>�Z�>�.���� �4�a��Љ�V?�̎?���,r����=��&>���u,?:\?}<����<r>�J?�ă?�%^?�U�>�a�LW���з�V����;�>���>$��>-'$=Nq>������'�>6�j>pɼ
� ������A���>D�A?w�?�f>i�"?}�#?7)n>�9�>z�M�����{@�f�a>���>Ȟ#?�x�?��?�,ɾ~�*�r����ţ�I\�6�>Dn?ȁ?�2|>&���k�t��쑼O�k�V�}�4@�?�[]?��Ǿ��?�#�?�wV?v?�9H>(��;
}���N��z�=�"?�P�fA��q&�_����?ڴ?���>�A��@�ӽ ?����8C���)?.(\?h�&?~W�+a�P>þ�:�<�!'����&<�yB�Z>�">k4���=6<>��=�l��c6���P<��=+M�>q�=dg5�ԗ��$=,?2�G��ۃ���=u�r�TxD���>%JL>A����^?jk=���{�����x���	U�� �?��?Ik�?B��a�h��$=?�?H	?�"�>�J���}޾��}Qw�I~x��w�w�>m��>;�l�E�%��������F��
�Ž�k��s[�>�y>�x?D?�)$>��>3)t���T��>����L$e���)�ۀ@��9�I�*�Xؕ�F��.���,��I?��Ͷ>���yZ�>�k ?>��>X�4>���>�P���a3>��@>��t>�9�>2>�bl>A�Խh�<�̻�KR?����%�'����²��g3B?�qd?S1�>ui�;��������?���?Qs�?=v>h��,+��n?�>�>H��Vq
?�T:=Y8�;�<V��t��3��)�1��>�D׽� :��M�Dnf�sj
?�/?�����̾�;׽���Ln�:�D�?��*?�,���G���t��W�bMV��-���u�����2��rt������0~�P���s��	�=(�%?yV�?P�������{��m��-N��7C>���>s��>�۰>��->v��W+�zX���h[;���>�r?E�>��>?9`M?�5O?&:@?�t>��?�T��P�>A��>4��>��>�9?�g?�@?�:<?��`?0N\>�B¾���2j��'T:?H�1?�6?S��>�a&?�o�����=����Kg�/3m�6�
�uW�=��>gP�E���ywE=8�P>�Z?���{�8�H�����j>�7?�|�>���>���6/���<��>"�
?�8�>� ��r�ed�*Y�>Y��?����=W�)>��=.ԅ�M��{k�=�¼7�=�灼�;���<��=|�=Sh~�����kT�: 4�;�X�<���>X�'?�x�>��(>C���e,��F�c1:>��u>|��=��Ւ������ Bp���,>~!v?��?��i>���=�u>�Ǽ�����4�v/y�k�=�W�>L�*?��a?j��?�#?��<?m�N>���*\��#͈��`U�n�?�!,?���>�����ʾ�񨿦�3�ӝ?p[?�<a�9���;)���¾Q�Խq�>�[/�~/~����"D��ׅ����/��,��?뿝?�A�j�6��x�ҿ���[��s�C?'"�>Y�>��>N�)���g�v%�2;>1��>yR?i�>[�O?��y?}_\?�]>�Z:�$��������Bo���>&�A?s�?���? w?�O�>��> )��~�]���kN#�FC�A����Q=��]>Rؐ>���>|��>f�=��Ľ\c��#�?���=mD]>R��>nz�>�3�>��r>N�<�TT?�� ?V������g���_��a5�wI?ᴞ?��2?9�n�0��sF$��z����>��?���?�-?��}��=�/��'Ͻ�@���_�>�\�>5ؙ>LJ�<��=0o>:A�>bP�>�����"%��B�U�QQ?z�<?��<��ſ��h��c��,���7�!�N����M0�Y 0�+�8���=lř�0½�����T��ʢ���&�������OS�0�?���=ڏ�=	�>~D���Q=��<c.=�=�|ν��~=��d�2�?��̨����Y��(-�����,sɾO|?��D?!-?�zH?�8[>�>O*��>=���@?�XT>�H��u����e4�%��C����ݾIپNd_��ř�
k>�pm��g
>50/>A:�=��<���=�Do=m�x=M��;5Y!=Gȶ=ZT�=���=�*�=�C>:e>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>X�6>�w>]dR��y0���W��e���Z� �!?�{;�6#̾��>���=`�߾l�ƾ&�0=�4>�`=H��Z3\�Nm�=��v�|J;=2f=un�>*ZC>���=�I���T�=�]I=���=rP>:7���t;��%���9=�=�=W�a>~f%>ތ�>.�?�[0?[d?*Q�>�Dn�3$Ͼ�0��~8�>��=t_�>s�=�MB>Q��>�7?&�D?`�K?�k�>��=��>��>��,�g�m�od�#ɧ��T�<���?ˆ?0ϸ>BQ<܂A�/��ef>���Ľ$x?oH1?�e?#۞>���޿��&�#�0�lŬ�ѻ�L=Xj��LQ�!���aڽ:�=�7�>�|�>K9�>�&w>+�>>"�P>���>��>64�<J_�=ε�q;�<����r=Nd�D�
=d�
�?�;����m�9�:X��^��\Y9���<�?�;
�j=U�>F}8=�;�>���=��ξJX>�{B�f���y=�6���5��#m��u��;5��WR>�w)>q��ڗ��?��a>l%U>`�?�&v?�5�>H�1�`�������C������8��=�"5>U0��R*���H��I��A�a��>�"h>uB�>{�e>o\)��0H��]�=�뿾%8�}��>�~/��g:���C��x�Ӛ���d����X�Y��<�wG?泍��{7>�x?��A?��?�ٺ>�&^��lξ���=i���"<���_��@o��Z� ?�(?0��>c���\�H̾$h��?�>��H�r�O������0��Z"�z鷾L|�>F��AѾR3��i������zB�\r���>�O?iޮ?��`�b��lO�ǒ�۴���9?2[g?�7�>�@?T.?�?��ō�,a��ل�=��n?��?U:�?9><~�=Ę��S��>�	?p��?O��?��s?��A�4��>랢;5� >ȋ�����=��>�8�=�R�=R
?9x
?�A
?����&�	�rm�C�!^��S�<��=�>"��>�tq>u��=ah=R��=*\>쒞>�~�>��d>��>�S�>���؆��a?��P>�A�>O�'?dz�>��>%<�fj��uA�x�1�o?����D�	rD���ؼ����R�=f*9<�q�>܌ڿ��?O�*>�/�0(?r�*��:==�>��I>�b�~��>�2>�ap>���>�y�>��=��>M>u>33ӾRE>����h!��8C�{mR��Ѿ3�z><���K*&�q��_S��dHI�tb���Z���i��/���G=�v�<]H�?N��o�k�$�)��d���?�X�>6?Rڌ�S���>���>]Ѝ>7T��}����ȍ��Xᾗ�?>��?��w>h1�>^?P�?�@����;�1$z���k���=���G�%�W���:��)��Nk��2@?~U?��K?ls>��h>fŕ?��K�"��HB�>4#��D?�(f�<��>2���LI��ž���>�߽�_f>�J?�sz?h�/?.���ȽCK>y�?�̃?�Rw?��-?�cs?[R��N��>?�r>�g�>S�>٭V?�M?ރ4?��>��?�ݍ=����{Q���������}�<�$���Z=�e=G�ɽ>ʽ��]���B=m�?����BN�=#���4L�;�%P<�i�=�Z >�*�>�\??��>*�y>�6?���.�8��1��#/?"��=�P����������Z���>�l?���?ŃT?rG>�^F�,�F�F�!>���>��$>�r?>;d�>z�	��ep�1��=�y>�#>[͵=�hs�e��*	�ዊ���=d>��>2|>��ݴ'>d{��`,z�z�d>�Q��ɺ���S�!�G�n�1���v�_Y�>��K?l�?Q��=I_龓4���Hf�B/)?>]<?�NM?��?��=M�۾��9���J��;���>Zh�<��������#��r�:����:��s>2��9�����1>4�#��%��Jv��Z\��s�=P@>��(.3��6��˾ґr�uм=��6>���=�+�L5���L���Y?fM�������pk���3>uN�>���>$��k8ֽ��J�Ԟ����=W:�>��C>X>�?~�R3V�`���>�bG?�I?9&�?T)���S�.�g���̾�+���$?�=�>uR?�6�=�R�<����-!���j���&���>W>
?ŉ���^�D���۾=\����>��?���=�1?�sk?��!?|�t?�I?3s�>Xg>�Z��I��'B&?|��?�=c�Խ�T�9�F���>΂)?�B���>��? �?��&?�Q?e�?s�>�� ��A@��>�X�> �W��b����_>��J?��>�>Y?lՃ?T�=>+�5�i墾F����u�=�>Z�2?�4#?�?e��>K�>���aU�=���>gc?��?.p?���=��?�.0>�/�>ᮖ=ٟ>)��>d�?��O?��s?��I?�D�>$t�<�G����2hs�G�C���;C�J<�-y=��`lq��v��<<�;�x���Ƈ�����D�6��'�;�_�>��s>�
����0>�ľ�O��,�@>����O��ڊ���:�A޷=0��>��?@��>_X#�$��=���>�H�>?���6(?��?�?�";��b�[�ھM�K���>@	B?q��=��l�����m�u���g=��m?��^?�W�C&���_l?\i?��־��(�ۑ�K���.<���Zu?N�?f����ܢ>�e�?쎍?k�?�A�<��X�/����)p�A���3?]>��=�����i��i���[?�{?k$F>�m�>�����䪿?5��Ƥ$?��?_V�?xa�?x>��h��"ۿ_�߾ܣ���y?v�>���/�2?�r��8Ҿ����FM�5��ͯ������!Q��k�ɾՍ ��x��%�ֽZc�>p�"?��c?~7R?;c?��јc�aYY�{g�$�O�J����V��MW���A���#��Â����r(��V�D�f�=��}�@D�G;�?أ&?R5��l�>�Ι�ȓ�CgϾ�pF>y۠�w��6��=����,=�M=�]j�[9.��W��y�!?찷>@9�>s�=?F�\�Ξ=�Z�1��6�._��r�1>�t�>½�>�d�>���;�+<�K�Ͻ�ľā�����f>"@Z?�9C?y?�ɽ�N5��|��v��2ѽ�,��co>���=�>=[����C��H2��?��q��  �����Az�'QX=g&:?�Ҋ>=pe>Q��?���>���ך��
��SW7�?9=ށ�>��Z?S�>�>v(�b'�F��>s�r?�ɬ>f�G>*SD�N1�IM���jD�fi�>z�>�8?4�=�A3�"6Z������2���oE�=%Q>�
�?m�^v���1u>�.�?����8�!��qr>��>}=j�97����0��>�1�>D�нM�7>nƾ�����"6�l�+?)�3?����!M;�w��>��3?%B�>�\I>|҈?���>��𾫠�=T�?\[?2�A?b�B?��>���i��S;��
�"��=��>��q>�.��S�>񺅾�]��B���w=5M>��=������/����s �=gb�=k��=�0�/�E�
	�ޯ3�	O�Z��#��M�=T�-���I�o?��~���LZ*�o|�ى�<e�ɽo�`�TCY���A���?���?�1޾XC��#��wˁ��
�Y?�@W�]n�#���}������I󾳛��v�
�w�8��.���>�G�*?~�⾮ ˿G�����C�?F�>uǉ?�T��N��FA�h@>��<�3H��ݾ�b���\ѿ�����IO?��?Ug򾏍(���>�>} �>OHc>��ξ{8��M�	>t�?�0?�k�>��Ѿ�ٿ{��O��=~�?�@@}A?��(���쾘V=E��>0�	?�?>$T1��I�v���oT�>q<�?��?I}M=m�W���	�-�e?{<�F�(�ݻ��=<�=�G=�����J>�U�>'��4TA��?ܽj�4>4څ>�}"���ӂ^�`��<��]>��ս|;��5Մ?,{\��f���/��T��U>��T?�*�>V:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�݅�=v6�쉤�z���&V�}��=Z��>b�>Â,������O��I��W��=oh��(ſ�&�X�#�ݿ�<u���>(y��㽰�����T������g�K�׽�9x=s[ >�vY>wj|>b'G>��O>�/Y?��m?���>���=ێ�
���Ⱦ=ެU������������/�'&�������5�A����^U��d�<;Op�˅��-;��r��LS�N�O?�.v>C����)�	2';?��g]��=�=!|ż]'ؾ}t��3O�(ۦ?��+?R��M
#���5r�T@d���Y?.��!������{*�=x�����<Bb�>?������>��T��p0?�?�k��m����*><M ��#=G�+?ș?��g<BЪ>�U%?B*�c?㽐�[>U�3>D��>-j�>��>�5��]}۽V�?�T?2��2�����>�����X{�2`=�r>6 5��g���[>z�<�����US�y����:�<�'W?���>��)��	��T��O���==��x?�?�Q�>�~k?L�B?؟�<�e����S��"�LRw=,�W?�&i?��>�g��y о�v��z�5?!�e?�N>>*h��龋�.�(K�m'?��n?+\?�����v}�
������t6?Mv?�j��ϟ�C���+����;>m)�>�?��:�	-�>]*;?�'��?�������YB�&)�?��?#&�?cv}=���a�=?���>H���7��&\��眩���X=�Y?m���P��P�,�&�Q���3?���?�.?to���x���=ݕ�+[�?&�?4���N�g<2��Ql�zp�����<3ī=���H"�1���7�3�ƾ �
�W����������>�Y@U`轱+�>F8�6�zSϿL��I\о�Tq�4�?v|�>�Ƚ{���r�j��Lu���G�{�H�w���'��>>P�����|�F;����	T�>4H����>�JU�x����ў��RF<B;�>G��>S3�>-��T�����?����.ο�������f�X?�n�?�5�?x?��B<��x�Ai|�}�/0G?��s?g,Z?��$�,�]���:���k?T	��=c�!�4��C��mP>O+?��>sG.����=��>�?�>X��='�2���ÿ�s��RV�.�?�6�?K꾑h�>�_�?��)?����[��%��(�&��R:��B?2�7>eǾ�&�ZL>�='���}??�5?����h�!�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?��>�?V��=��>O��=���1��3#>��=s�?���?߈M?�4�>�B�=t69�1/��PF�"ER� �'�C�۲�>��a?��L?Mwb>�X��X�-��� �Ͻ�>1�`꼽�@�:�+���޽}5>4�=>g>_E�":Ӿ�2?h;:�a8ۿ�>������34?_�^=��?���=Yt�Z��^? �>�)��Q���(���@�5�?I��?N�>v����}=��=g��>o��=bK�9
��DS���>��H?��,ڙ�>!���	>���?Q�@��?�AU��8
?���ݵ����}�� ���6�x��=��7?ͺ�ǁ{>�
�>yH�=��w��謹�Tt��5�>)߯?=��?��>��i?emm��?���:=)�>�4e?��
?F�ݺ���J><�?>�������9�u�d?��
@
?@<�]?M_����ѿ4�������d��RC�=���=;�G>ݽн �1=Y��<6S�<_M�;6>EV�>w�a>�f`>��?>&�3>�>~���e� ����ϲ���?������&r����6ڃ�����ڰ���ž|��� Ow�1&_��U���5�*%��z��=�V?@�R?�o?�?��L��E5>����;�<���1�=��>�13?
@O?Tg,?���=�㎾H�a����H۫����P�>L�d>a<�>�M�>j1�>됀<<[B>�>�Pu>`a>9��<�q��OB(=��N>�.�>F��>T�>E,>��=%����W�y�����ߚ*��]�?��'^�ț��B~��K�����=��/?��y=�����ɿ�����[?�!��K��O}'����=��M?�a?���=��˾����C�Z=��ܽ�F���=uQ�J���:(�$�7>I�?�Gg>�u>�3��Z8�0�P�O��z�|>�(6?Ճ���*9�6�u�B�H�%�ܾ�M>��>,�?��u�����%�%^i�8�{=$P:?]m?蠲�������u�1p��E�R>X�\>0�=�<�=��L>�~c��vƽ�G��a/=���=��^>LV?�+>&��=}ޣ>�X���OP��{�>Q`B>�(,>@?�)%?���Zٗ�������-���v>�H�>

�>S_>�YJ���=f�>\�a>�W��q��.�?��XW>�~�\t_�{au�P�x=(�����=8
�=�� �H=�f�%=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�l�>����[����q�u�!�#=y��>�:H?�Y���P��>��w
?�?�^�ڨ����ȿ�~v����>P�?���?��m�[@��I@�׊�>i��?GaY?�Qi>nf۾�CZ�>׻@?BR?�
�>�@���'�r�?��?߲�?�';>XS�?�g?Y^�>��׼��<��t��
���q@������Ƥ�>J��=$ݳ�|�G��ב�1���y�k�nS!���c>r.2=L�>.	�4~̾���=J�\͌�w:�ڡ�>��i>�Q>㩜>^"?f��>O�>�R�<鸽hc���B��Y�m?�"�?���F(d�ϬK����>cv={��>�w?��>�2�&%�> �d?�̋?�s?|g�>����'W���(��"D�>[04>�1>��8?yz�=��s���ͷ�v��>�C�>�kP�������N�N��Ś>ν/?�t�>D�M>D?��*?�d^>w��>*�4�SՕ�&<����>��>	?�Ņ?P�?񮝾
/-����M_���`��*>	�u? !?��>x�������]U[�oM��ǈ�>b�?�_s?�� �^�?Z��?��M?��V?���>��׽�Ͼ����g�n>�c$?��
�.�@�%%�L�*�Fy?B�	?h��>5]��:ٽ�T��i��Ȇ뾳7?�F^?��%?�L�k�d���˾��<�R���m�TO�;x�K��>]�>����Ő�=X3+>�B�=��}��C��ai<}M�=��>L��=N�8�����&?/�ͽx������<sC���a�l�&>�Bd>!�Ӿ�or?z>�+�w�p>���M��'���b��?�Y�? [�?&W��s0v��I?T�?�v?M��>�~��[g���߾����ZP������Z���>5��;&b��r?��FR���%��5��k����.�>J��>�G?~��>�m1�z��>���]N)�'}��W���Oe��a8�S�R�t4�E��5��ϥ�x=��̾�,a�y�>n_�����>#k?��C>0�>Vq�>����x�>��>dh>l��>�/>�+*>�a>�\۽��F��,T?%�ܳ&�V1辶滾�5A?�f?���>��)�0�����F4 ?,��?6�?Jc�>@vd���,��.�>���>�y���?��	=B4�C�2;5���k:���f˼���>� ��u=���L���]�!?�?Q��WϾ?��{��}*o=�B�?$)?*�)���Q�}�o�	�W�\%S�o���g�0����$�;�p��鏿�b���#��	�(�+=�z*?~�?���^��E ��p'k���>��Yf>���>�>"ھ>�nI>��	��1��]�_7'�󻃾z.�>�>{?��r>�g?�(6?h0?acO?�1�>Ǿ�>����ʼ>�E7>܏>�?�J?oRF?/�/?��??�/?q�=}����o
�΄��3?�Q?�=�>d��>��?���9�Z�r2i����=Z� ��$��
�=tp>�@��Ľ���=��4>�X?>����8�L����k>ʀ7?��>��>n��9-��
�<��>�
?ZF�>d �E~r�c��U�>���?���A�=	�)>T��=w����Ӻ�[�=������=�3��Hz;��^<���=���=�?t�6B�����:i��;l�<l�?g%?��8>�m'<�f�;S¾�G3�i\��Ư?�E�>��p>N<�4G�VR���u��S[>���?�`�?'�P�m�=9�>����B���!����W9>� ,>6�O?��?�/�?��,?dVL?H�k>�±��c����������?x!,?��>�����ʾ��Չ3�ܝ?i[?�<a����;)�ސ¾��Խױ>�[/�g/~����?D�����V��5��?쿝?GA�V�6��x�ۿ���[��|�C?"�>Y�>��>T�)�|�g�q%��1;>���>kR? #�>�O?^<{?C�[?�hT>U�8��0���ә��l3���!>�@?���?��?�y?t�>|�>?�)�p�*T�����HႾ�W= 	Z>���>�(�>��>���=� ȽbZ��|�>��`�=�b>W��>��>��>l�w>cJ�<d�G?��>$���D��n_������?mE��Mu?�n�?�+?T�=���5=F������5�>��?q$�?��*?/JT�EO�=I�Ƽ�ַ��s�$Ѹ>���>���>?�=��P=��>I�>��>'��d���8�BS���?@F?F�=Xƿt�p���o��?��O�o<�ᓾؤb����=�\����=;���������]�l�V��B���1y����z��Z�>Sz�=�M�=���=M�<7|��n��<^bI=�%�<��=�|k��]�<��0��$��9�����]h<�yI=<~�?�ʾ��{?VH?�U-?*C?-l>ޯ>?�8�]�>K=���?��M>b�T�B����FA������&��\۾��Ծ��b��E��\8>��Y���>�>+>&��=��f<V��=$x=��=q�����,=���=a2�=]�=B^�=6�>�.>�6w?X�������4Q��Z罣�:?�8�>h{�=��ƾq@?��>>�2������zb��-?���?�T�??�??ti��d�>K���㎽�q�=P����=2>u��=x�2�S��>��J>���K��D����4�?��@��??�ዿТϿ4a/>�P7>�,>[�R�{1���\���b��<Z���!?VG;��Z̾�@�>1��=�J߾X�ƾc�-=q6>+b=F_�aG\����=�={� �<=b�k=�ى>$D>�/�=�w����=}I=a/�=z"P>+~���G6�!,�r�3=I�=��b>'�%>��>�?�a0?�Xd?�6�>�n��Ͼ,@���H�>N�=�E�>���=�rB>Ґ�>��7?��D?��K?ͅ�>(��=D	�>X�>X�,���m��l�ͧ�Ӎ�<]��?tΆ?�Ѹ>F�Q<�A���1g>��*Ž�v?�R1?pk?x�>�g�:�޿� (�g�1�y���҇���=gp��w�<����� ��0۽���=s��>dT�>�5�>\�h>�')>uD>��>��(>��<��=O�!��bN�[χ�3\�=��<��<Ǚ�~��#/<i#C���@�K<zA�;�*=�;<lr�<S��>��=%�>� ��� �D�.>�3��Z_�>EK>�^���k���x�����_*�M_��>LA�>�~�=5�����!?] �>`w>
e�?��f?���>;����s������eb�S����M0>��=X���.�INm��$S����9��>X�>�>��l>�,�8%?��w=x ⾏d5����>�f��l��3�=q��<������i���ۺ�D?E��d`�=t~?�I?4��?u�>�y��9�ؾW0>�G���=���q�#E��C�?[	'?���>[(�U�D���˾�q½<��>�oH�BP�u���0���%��J�����>*O���%Ѿh�2�&G��N��6HB�R+r�"��>EP?��?N�`��[����N����
��H?�Mg?+��>j ?	�?�j����[����=�#o?��?	5�?p>���=�g���@�>��	?�?��?��s?1B�O��>?�O;/�>}4����=k>���=�G�=��?�
?O�	?����]
����P����]��n�<���=��>%	�>XGr>���=e�W=�Y�=p/\>�A�>zc�>?zd>am�><9�>������b7?�L�=��>̥(?KGg>�M'=�.Q�<e��/t�=�5�
���_W)��+J��)��P���{]=��&=w�?ׅͿ:v�?��>0�M�I?o%��:�l!>30�>
�c����>DԽ>���>��>�Y�>�b�=Q�I>a�>�qѾ�Q>�g�!�ND���Q�$>Ҿ�ʁ>�֜��0���	��k���sG��7���>��sj�t��� [=�z��<ɏ�?���d9k��k)�g�����
?�׫>�4?b���W���s�>�@�>=%�>������s�����" �?��?3ܑ>���=Q<\?5W?F`L�����l��F��9H�F�H�éC�6Й�n����� �s�оC�?�>�?��Z?�W�=!z>z�?�Ay��"辴K�>g�0��fR��]~<S� ?b�Ǿp�r� �������Yn>��b?y��?�F?�
�hq\��N�f?w̅?/~�?�^E?�s�?������r>M�0�/>�-&?b%?��O?��G?���>,Ѱ>�(�0 ��Gν�	ɾ�̽�р��8<5Q[=��3="�<�y�_J=���=��E���b��'Ľ¢�l�o��u�<�={>9��>�]?��>�Ņ>��7?�\� i8�}˯��/?X�E=$��○��������>�j?�߫?٘Z?� d>��A�]_B��2>=�>�E%>#�[>�g�>l����E� ��=�'>�>"�=�DI�f�����	��w�����<5 >���>;�}>�����%>h���+/x��e>lQ�	��L�Q�+�G��1��u�v'�>9L?S?*$�=e꾇����)f���)?�K<?X�L?�/�?��=�'ݾ�9�_zJ����(��>?��<�6	�~���y0���f:�ߩ9;��t>���0:��w!i>�K%��Q���{���M�����p��>1��m;���rd�k幽�O<4Y>�Ѿ�D,������pR?'>�c�����ɽ�����=�h�>W�v>�U�+���	d�RP��j�>g��>ٵ>��G����@V�I��t�t>�qM?ݍJ?<��?x�̽�z���?������E�!��/!?���>, �>�&>���=�d ���)��)f���<v�>c��>���h�u͍��^;���m&�>g�?�$>!l?`_??sb?��#?1��>u�V>�V	�]?���@&?B��?=�=�Խ��T��9��F���>?�)?+�B��Ɨ>ъ?Խ?��&?�Q?��?�>� �"4@���>�S�>E�W�8h��S�_>u�J?���>�DY?.փ?��=>�5��Т�Q��d��=)&>n�2?3-#?��?��>Έ�>J���A>�>� n?�9�?�[?"���v%�>a�<>�?O��> �p>�6�>b��>�\C?Zo�?�$?�I>#<��ƽ���=�#g�0���$_��y�����=t��<.�kp�X�tN��轮!�<����[��e\�=}��<��>��s>���A�0>��ľ)��n�@>�֡��꛾B���[�:��^�=���>n?	��>T#��=�s�>�0�>����6(?��?�?��5;�b�<۾[�K�d�>QB?y�=��l������u�Ng=��m?��^?DW�E����of?=�Z?��۾��P��_��i�q�v�;�
R?�?/��>�R>|h�?��?��,?��^�χS������e���¾	eG>Ы>jW��7I�5����n?�?u��>)-�>u|����������2�J?���?Wb�?�y�?]�=�-]�Rӿ��J���X�?���>G���r�+?Ü�A]ɾ�Wƾ�v��r��:2þھ�Yʌ�����f��m����߽Q">_�?�G\?q�d?'�e?��C�p���k��\z���B���ݾ&0��	a��)>�mT"���k��a ��꾈}Z�È>��{��N�&�?C"?��1��f�>m�������B>Z֓�E�.��>=�ɍ�K�[<b;�<��e�1.�꧞�Ȓ$?���>��>x7@?d�]��cD�?9�s�7��#�G�@>�>�VQ>�l�>
�=��B���׽�rǾ%[f�tZX��O>>Ra?�qA?<{�?�&���)?�����6�<����پ� >�ϗ=��n>��e�Í+�? /�r<H���y����������#�W��<��<?n�>��<>���?�+ ?��^<Ǿ�̇�2��K'�=��>�/g?���>�>�7,����� �>G�W?���>H�>��Ⱦ�Y7�i����p��i4�>Z��>�T3?�10=7u��zP������|���c&�"� >��??�쥾���̡�>�\?�"R>�㪼�y>������P�>?d��䉾�>�0?�{�=5d�>��ɾ��T�� ��c�=���*?&�?����)��)v>в!?6K�>\��>�p�?N��>�`ƾ�f�*�?S�a?f/N?O	B?k��>g�<���s�ѽB����9=�օ>��i>�"I=6��=!�4lb� ��q��=͇�=M�w�ڽ��;b�Z3�<��=�x<>�߿�wR��k ���2�l���F��G���>8BG�~_;��톾j�žg9���ƽ�6�=�l�a���)+��������?�+�?����[���)У�ܛW����I*?��J�Wj��擾=��g�Q��~�:�
���7���3�9�G�1�/?��վָпO؛�Zv�Xt.?��?>��?� ��W9�*�n�\G�>OI>�ǵ�ֻپ���e�ÿI��M4t?J]?N� ��/��p�>�i�>!��>�	>�A�^��Th=�C?�7\?���>�����ؿX��@��=��?H@�|A?��(����V=}��>D�	?��?>FT1��I������T�>q<�?���?�{M=i�W��	�9�e?	<��F�'�ݻ��=<�=�E=z��z�J>SU�>���SA�7?ܽ�4>3څ>�~"�����^�&��<��]>��ս-;���Մ?p\��f���/�S��}f>��T?�.�>���=��,?�6H�zϿv�\�U/a?:1�?Ӥ�?��(?⿾�՚>|�ܾ��M?@6?��>�T&�ؽt�I	�=H`�0֧����KV�� �=}��>GQ>K�,�����tO�Ø�o�=z��g�ƿV%�Ԣ �@1�<�k��g��Kν�����7e��=��]�u�n��7Vt=���=�/O>�+�>�]O>#\>J"Y?gl?�2�>��	>�(��������Ͼ�^<�����P���� �#M�����^�ھ����l������ƾ9C��ɗ=�b�˱����7�{�Q�Jd=���T?Lt6>O�ɾ��,�I��C����z��AΖ=R���J�Ծ���&L��?��Q? ��F4�ȗ�l���^��I?^��(C澺󢾸p�=q��=r����%�>���;�K��=��VT�%G0?f#?b侾�{��*-,>�x ��R
=�-+?��?�=y<4�>.S%?4�(���ླྀ�\>#w5>��>0�>�	>L���_ڽD�?�T?��9���Nk�>A���'�}�W[=-	>�2�VG�8DZ>a=�<����vK�񨎽 ��<(W?ś�>��)�2�Pe��"�<0==�x?A�?o6�>,}k?��B?W��<�g����S� �Yhw=��W?�(i?V�>����о����5?��e?{�N>�Zh���(�.��R�6#?��n?�]?cz���v}��������m6?��{?�Dg�ܚ����������}>���>�?	v:����>�17?�#�Js���	���?7�_��?V�?	��?_DZ=��ӽ��=�J ?���>����'�_�D=�u�����<�Z?cπ�ׂ�����I�6v,?D�?��?�3���	�ʽ�=�_��pw�?a�?�'��3i<È�*�k���t.�<�o�=ŞV���B����8�l�Ǿ��	��>���f,�>ш>��@,�t��>�"=�HL⿿xϿ�1����˾�q���?#�>8�ܽ�L��cNk��o��;C�w6D��0���N�>��>,���}���~�{�,r;��4��u�>a����>��S��!��o����6<��>Ԩ�>��>9���潾�ę?�b���>οs���ϟ�d�X?�g�?�n�?�r?×9<��v��{���Z0G?�s?DZ?;v%�B>]���7��rk?�߭��/a�v�5�XdE���U>؟0?�Y�>�-�t�y=J�>]��>ֲ>�U0�a�ÿ����#M��}|�?}��?i��*L�>���?�*?���yv��^b����&��eܺB�A?|P7>fȾ~�"��A<�1���)�?2/2?ӆ����]�_?*�a�M�p���-���ƽ�ۡ>��0��e\��M�����Xe����@y����?N^�?i�?ٵ�� #�e6%?�>d����8Ǿ��<���>�(�>*N>lH_���u>����:�i	>���?�~�?Qj?���������U>	�}?���>`�?ɚ�=�6�>W(>9��%��j�>$�>o����?�M?�m�>�F�=���� �n~C��7S��v �
GD�S�>`f?��P?7τ>dy��G�6+�L��E=A���; �)�ȼ�=��B>�>#�>$�1�.�ƾP�7?u5�_�ݿ?���L�{��	K?���=5�?���䎾WK��c@y?��X>��3��b��h���K@����?��@�{�>�@��=<�=�H�>�Y=��@�r��<�^|����>�Z?~�l�lP����b���k>#��?��@��?r`x���?P
��y������K�^�$��`�=a�:?�A���_q>,Q�>C��=.!v������s��ˮ>�o�?��?C��>rGd?�Qh��1��V6=j�>��S?|?�Z=���[>�?�	�/x��� ��a?a@p�@+V]?�F���1����������}h>9�=��:> ���#z�i�
��h�������;�3�>Z$z>A�>?��=�z�=� >���-��v򝿕���\�=��T�9�������v@��s�%�t_�����e+���*��%H��a���m;�=wjV?<U?��x?a�?��Z�8�8>Ha �TDO=b���OS=0'�>�K5?mS?�e+?q�=�a��N�_�=�y�N>��ʹ����>^�W>���>ȝ�>js�>�Mk<LM>}�.>̴d>��=ٿ=cB�:�:���G>;�>U��>ӈ�>74>'Z�=�ٴ�8��
t��(������?�Ҟ��jO�8��Z�����z��-=_�1?I</ƒ���ɿBǳ�c�T?K���DQ��2��=��C?��f?�v�=�>��G�"�<�Q
�G�K�N�*>��?�󄮾��!���>�c#?��e>�u>L�3��8�A Q��|����{>>�6?q��I9��;u�:�H��!ܾ"M>�i�>�B�1}�ź��Į~���g���|=�:?��?k���4Q��ʮv��y����P>�=\>��=qv�=glM>�k�}ƽ�I�_?)=���= ^\>qV?��+>b��=�£>�h���PP�1w�>JmB>C,>�@?0.%?���`������5.�K%w>�`�>�"�>�O>:uJ���=|�>��a>�p�b8������?��2W>�J~�`_���u���x=89��[��=S��=|� �U/=���%=�~?���&䈿��Te���lD?Q+?� �=�F<��"�D ���H��C�?q�@m�?��	��V�.�?�@�?$��}��=�|�>�֫>�ξ�L�ȱ?��Ž3Ǣ���	��(#�`S�?��?��/�Xʋ�.l��6>�^%?�Ӿ�,�>0�����������v��l1={D�>�3H?�U����W��SA�m�
?�X?���-���|Nɿ��v�*-�>*{�?�͔?Fzm�������?��c�>�j�?J�W?Re>YW۾�VX�FՍ>gA?U�P?�ʴ>c��J�%�$?I�?g�?ƥ2>""�?��e?=9?�Ma��hB�鎭�l��IQ��j	���z�>���=3���(a:�C銿�4���er��"���>x�X=�^�>�t ��Ƽ�*>f���F����Z�=9�>+�e>�e�>���>Y�>l�>���>�ʀԽ�$_�R�o�3;]?��?Ɵ���K�l���y>�ݼ����>
�}?V>t��EDA>vu?3Ϙ?�%�?��>� )��1���o��$���>��7> ,�>G�?0��[��[�9;T���>1s�>r������v�ƾ�K�����>C}?&E�>�`>>�?b�)?�Kd>���>�0��'����B�tK�>�v�>'��>Ѐ?G?�/����'��d���ע�^�b��m!>�x?6"?Ƥ�>����������q<Ƃ���W�?�wn?Z~�5�?��?RL?�M?�>����n~־����c�C>v�'?:�	�>��F�U�6��h?�7?�x�>�nV<�½ĶȽEh�;�ҾO ?Ii?�{&?]��ʦg� �̾,e�<����ϼ��~<~�_:]W>��=���� ��=HVQ>a�=L����i�s蔼��=s��>�x�= T�ڼs�*?��ӽ�<w��rf<5S}��TZ���>P"�>���{�j?�����������n��#���׉?�r�?���?����v�� I?V��?q?^��>�7˾r r�0��gQ����'�$��X��<D��>F=�վ�;��%B����/]�	���Q.�>l|�>_��>δ�>�QT=�>�C���%��羒��Se�O='��@B���E������^G!�Ҽe��þ:�w��:�>�'b�)�>p�'?�
�=p�=� �>e����>��>n�>W!�>��|>��>�W3=�[v<�O6�wmS?Tּ��o&�K��i���B?ae?B �>?h������H�d�?sՓ?�N�?ۅ�>d��L-�E) ?�C�>�
{�!�?^#)=�5�;�?<ੲ�	���\���̖�9�>��ٽ�w<��M�F�]��?�~?���)̾�ý͞��<G=�L�?��)?��)�ҸP���o��lW��T�y��5e��3��c`%� o��⏿:�������I'��Q=��*?�m�?D�������l��o@�=�d>��>>P�>��>��@>��
�0��B^�"#���}�7q�>\Vz?R>Ph?m�F?��B?�\r?��c>�	�>���h��>��=�>j�	?V�G?s�3?��??n?N?>Ĩ=�y)�� �X����<%?	MP?�?Q�> �&? ����1�������뼸cK��e,���>�JE=�f�@dq=g��=��">�X?�����8�`���%k>��7?d��>��>����,����<��>�
?�F�>5 ��}r��b�~V�>s��?R��h�=��)>���=������ҺY�=������=�3��X{;�a<I��=-��=�rt�J$��S�:΢�;�m�<��?� ?l��=�2p>�CU�?����A�����M?�o?J_�=�������A|����k���>k��?���?ţ3����=]o>����G%��,����J��<�Na>%�4?�v�?>�?_?�WG?,�A>����ɗ�X���R׾��?r!,?"��>�����ʾ��ɉ3�ϝ?g[?}<a�����;)�ɐ¾x�Խ�>�[/�S/~����>D��셻���B��.��?뿝?|A�U�6��x�ۿ���[��p�C?"�>Y�>��>S�)�l�g�p%��1;>��>aR?���>7�O?+7{?	�[?��T>�8�O���̙�ۥ1���!>u�??Ƣ�?��?�y?�t�>m�>	�)��#�4:�������c����*W=��Y>�u�>�>�>���>ȧ�=^!ȽGG����>��V�=�lb>hJ�>ֆ�>/�>�w>�<��F?K��>�����	�BC��w�;╽}p?Qb�?j9%?A��<%�R�K�3���j��>v��?���?�2?��p�:��=(��N���k��6��>n԰>�l�>x�"=��=�Y4>7��>*U�>�;�9i�?�/�T₽~�?GjF?�E�=R�ſ�p��w��C�����;�W���te�K}��qX��e�==T���P!���5\��ǝ����������3���4y�= ?�Y�=�`�=�G�=@|�<����<{�F=�q<�Y=3�w�JIr<�r'���=�
��iĻ�<�B=!Y��r̾1}?��H? �*?UC?E�w>�?>:�,�k6�>1T��%�?�S>�Z�OS����>�9 ���ڔ��ؾoc׾`d�d��pQ	>�G�F�>3}7>U�=��Y<rL�=��n=%��=ݏ�9!�=K�=Nܾ=�X�=<��=[�>rQ>�6w?X�������4Q��Z罟�:?�8�>{�=��ƾr@?��>>�2������|b��-?���?�T�?A�?;ti��d�>G��m㎽�q�=K����=2>���=|�2�P��>��J>���K��?����4�?��@��??�ዿТϿ6a/>��2>';>��S��]2�+Pb�=�d�U�[�$K#?%:���˾/@�>g��=�	ܾ��ƾ@�<=��4>!�S=�;�i8[��S�=�t���:=&��=<�>��=>WŲ=�>���w�=n>H=U�=��N>X��^N��W+�v=e��=��]>L->	��>F?�q0?�e?u��>�m��c;�c���܌>7m�=��>�p�=�D>��>-�7?H{D?��K?���>���=]��>b��>3�,��Mm�"_微,���`�<�;�?OO�?N��>��O<e�@��]��>��ʽ�S?�/2?�w?��>=������	&��&0��wu��I��#��<�K�$$��@�������
�=��>*��>��>l�O>�y>�?T>S�>�H9>$D��Vu<`0P���0<�c�C$>��弘�O<���3��k���+[�19E�<K��C�<*��<{@=Q��>�">X-�>�޻�DF���U�>���Z��o?>�.���5O��oh��-����<�����4Z>�?.>��,=� ��;�?Sh>��+>��?Mj`?�v>_�ｱ朾'������?L�2�=[�\>�h��LxL�2�p�f�Z���ɾ��>@�>��>w�l>=,��#?�Gzw=���^5�:
�>su��z���-�E9q��>��.���&i��sֺ��D?F��
��= ~?~�I?�?ۈ�>�����ؾk$0>�W��|p=�
�Rq��W��y ?�'?���>-$�2�D��CȾU�����>Ų;���O�蓿F<1����������>Ka��a%ھ94��΄���%B�8%q�E��>K*R?��?��K�>5���+H�q}�q�����>�d?F��>��?>�?��������z�<ܘ=��r?4k�?�5�?N>K��=����^��>Yp?�-�?9Q�?&t?;WI���>к)<A�>��x�
{�=VB>��=�s�=��?J?1b?����}�����!𾼩c�9R�<��=(�>��>xe>�}�=��k=���=�6J>*�>Y��>U�t>3�>;J�>�>־I��=?�Y�=�ʌ>q�:?���>�SY=Ya���6������b���t<�L�]��u����u<׎G<�ݽ�&�>�Mտ��?~:>n� �nc5?�o�({����;*�]>}�����>�8+>I>�>F_�>�9k>I>�Q>I>k!Ӿ�+>X���o!��DC�5qR� �Ѿ�"{>j����&���������H��j��CB�D#j�0��GA=���<�L�?����/�k���)�)���u�?~��>��5?�͌�l���4>�#�>&��>���u����ύ�uQ����?���?��>@}�=��[?0�6?j+��)�q�4�|�y-K��`F���E��,&�-������w���оR�v?C�{?�b?�Y|=�g�>���?.�x�]������>�N>�o~5�t��=^�?���8zu�J�������mj����=S.�?|��?} O?Ҝ�q���t>��)?��N?�%�?�A?�|�?��G5�>��>��?��@?��?��0?V��>�	�>�/?�L��^���1�	�'��ێT�qH�ngֽ�##>��=NVD=?n��ꙹ�x�=皞=N5�f��m�����S<c��=�=��}<��>�<]?KZ�>���>��7?�J���8�z𮾂/?��6='��y��� ��r��=�ak?��?�l[?��^>WDA��O@�Ib>��>i$'>�nZ>a��>v��Y~?�XE�=�>�9>f��=w�X�!���
�u����<m>}�?|x�>�;�
/�=���"��S >���)��k��|�D��i.�����^�>�]?j�,?��:v����9O���a���9?�8?�!?C�?s�=�� ���8�@�W�Ե��L&�>1��=�&����b���l#$��=h�h>+K��KŠ��nb>Z���޾sn�p�I�S���<L=�X�p*U=��^־T%�k�=��
>q���,� �W�������#J?�_j=9q���>U��D����>�ۘ>R�>͜9��5u�Lj@�����Ŗ=���>�I;>�Ֆ�����}G�a#�J��>�&E?<_?lG�?k��BEs�ejC��N�������ؼ�?��>�$?W�C>@K�=��������Xd��\F����>m��>1��ΕG�����p��P
%�E��>IW?��>��?bdR?��
?W&a? }*?�??ُ>q��hض�."?� �? �I=dx��?��T/�6Y���>R?d:i���>�(�>?��;?�a?�?2A�=V?�7���s�>�l�>��R��ʭ�~+z>�W?���>^�Q?�\~?2��>!F(�b"��i���s�=�q*>c�$?� ?���>͟�>���>7�����=���>c?|0�?U�o?߁�=��?�<2>��>m��=|��>q��>�?nXO?�s?T�J?���>���<�5��29��wEs���O���;\�H<��y=��z4t��G�o��<��;�l���W����񼰻D�$W��;9�>��>�:���^<�s�k��ܿ�=��6�龎`��Ç��@>�>J��>)=�>>�����>��>.��>�_*���A?~v?��?i	O>�X��"�4lB=��>�8?dD2�4���3���]��ha��6�^?2�V?VJ�=Ԝ����i?j[N?^]��Z�4�_ȾPO�&O��k4Y?&�?�W���V�>�ـ?g�n?y�>�����>w��>��j�U��?���=�̊>B�
��FZ�[��>p6C?V˵>;�n>C:�=�w��=by�Ձ���&?��? �?n��?�(>i{t��^ۿq�������+^?;��>�*���"?�?�d�Ͼ����K����p�����az���˕��s��1�#��Z��ޗս(��={�?��r?�Uq?F�_?F� �*�c��,^����b&V����U���E���D��C�ۊn� N�����qs���dH=�ο��#����?�?Dn���>��������7=:�ɾP�O�������l�=)�>����༅���o5?#X�>�Hs>��+?ZIM�vZ=��PL�����Q��֧_=E�>�.>0�>&/�>;�>Y�=�Xܾ��A��Y>�6v>�xc?�K?�n?�o��*1�膂�s�!�Ĺ/�d���B>�h>��>d�W�H���9&�~Y>���r�E��Zv����	�8�~=��2?�(�>[��>P�?�?^{	�j���kx�1�1�l��<�0�>l i?�@�>D�>�н� �/��>��l?ب�>g�>���(Z!��{�
�ʽr&�>~߭>���>L�o>�,��#\��j��n����9��v�=)�h?�����`�I�>pR?��:J�G<.}�>��v���!�&����'��>_|?o��=m�;>�ž�$���{��7����)?۳?������'��Q�>� ?���>l֧>Kw�??5�>�������3�?|]? �K?��B?UL�>���<{3��ھ�#7'��D=dч>�R>�_+=&�=l���RY�����==�þ="��Ž��;Nu8���<;E�<mG,>hlۿ
@K���پ�	���@
��Ȳ��g��ݹ�vd��F���Yx����'��V��,c�\����l�n��?U;�?���-��k�������������>�q�`��r���&�����c����_!��O�g#i�;�e�G�%?=s��@ȿ�����־ޓ!?�?��y?�X	�k� �8��>X��<�9����㾄w��"jο����5_?0�>���XI��>�ы>5U>-�i>�ȃ��å�V$�<�}?{-?x�?��i��>ɿ�鼿�%{<�M�?.�@F�?�4v����9��>?��>�l>�"��V��U��Ma>6]�?|յ?ɻ�=:�a�~^q�Û�?�o�=V��bB�=��#>�} >�h>�_��Ï?>�%�>XUϾ��Ծ��]�>&�>����ҵ��j�'���g>�ї>��z�7X_�҄?ha\�a�e�Վ/�!J����>-�T?%G�>���=\�,?v$H�wϿ"�\��a?�+�?���?�(?�����>��ܾqM?tP6?�>1g&���t�Y��=���dv���㾑#V�s�=���>E>&�,�i}�iTO�+���ot�=����ſ��#��F����<7���U�o���齒z���,U��ݠ��gr������M=���=�R>3�>�3a>GOU>fhU?t�j??�>GD>q߽� ���dξ��'���}�����#���������|g��ྐ�	������iʾ�6=����=��R�ϣ��l!��fb��FF�P�.?�'>1�ʾ��M�4�<��ʾ���i�3ɠ�i�˾;[1�T�m�w�?�@?.���V����*��L뺽J�W?���������P��=_۱��=ڲ�>�m�=^����2���R�F1?��?OH���Gt��2>a^4�L�=��4?(2?I������>ȉ?O�a��湽.��>���>'p�>��>��6>c慨�Q���&?�I?�(�Tc���!�>o̾�������=�Z�='������$>��k���<������Ax?u��>Y)��e��-����ֽSd�>��~?�?a��>Ki�?��V?���=h��f��?�8�*V?��m?6�>�^��ѾP䆾�
?�(�?�y�>��2�JK��(���NR���#?�un?�u3?���;�r�͗�:��?j�v?�r^�Qs�����:�V��<�>Z[�>���>��9��k�>��>?e#��G��庿�iY4�Þ?��@���?~�;<�#�L��=�;?9\�>�O��>ƾ�|�� ����q=�"�>�����ev�����S,��8?���?���>o��������=ٕ��Z�?N�?��g<"��$l��n��Aj�<}̫=��.H"������7��ƾW�
�㩜��ҿ�ܦ�>Z@�Y�+*�>AC8�6�TϿ����ZоoTq���?���>��Ƚ������j��Ou�ɳG���H�����x��>C�>�L��N͑�_M{�_;�?�{����>��{�"+x>Q�a��|���!����<��>V1�>�y�>����������?2F��2�̿�=�����3
O?���?�ރ?C�"?3n�;�G�+��9�<�M?�s?([N?%b���\���<I�j?�_��bU`���4�iHE��U>Q#3?�C�>�-�e�|=�>)��>�g>�#/�j�Ŀ�ٶ�����4��?ŉ�?�o�I��>M��?Ws+?|i��7��'[��4�*��+��;A?�2>:����!��/=��ђ�¼
?"~0?�|��.�y?�6j�VƄ���0�F��z�> ��h���#e>/Ǐ�E�`�ζ��ǉ��"�?�?๪?�/q��e���:?���>md��۾yԌ=o?���>W�<'��=�� >��������?m�?��?�?����񛿟0n>�?LM�>j"�?Ք>>��?4آ��VԾ�,?>�}>�"�=�w>�b?��=?iu�>���=�1q�E����[��e�����v����> %Z?�Ĉ?�#R>k��8�T]���}�����>:���!����?����=>�>xnn��#��PN��?�q�Ŗؿ_i��/b'��44?���>��?m��԰t��C�*;_?�~�>�4�X+��&���@�Y��?bF�?4�?Ӹ׾�#̼I>��>SG�>E�Խ[��D���[�7>��B?�%C��
�o��
�>���?V�@�Ԯ?Zi��	?���P��Va~����7�b��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>!�l?��o�P�B���1=8M�>Μk?�s?�Po���j�B>��?"������L��f?�
@u@a�^?*�魿t���j���-����蟼�8=��3>�]���>�`�={V�=+Ƽ�9s=e�>�H�>�Ţ>�$>6>�?$>�s�o�#��Y������Q<_�^��9T�����2x�zI���6�m۾Gg��0.R=>v�>g�X���J�w�S=F��=��U?R?p?؋ ?��x�=�>�����#=
t#����=�0�>�b2?�L?;�*?�œ=������d�_��fI�������>�qI>~�>#G�>g�>f 29%�I>v"?>��>R� >=d'=
�i=?�N>�J�>���>bw�>q�9>@�>����F:��8�h�>*v���ʽ_Ǣ?_횾�J�(7�������7��ix�=A�.?ߓ>�ڑ���Ͽcx����G?[q��h���J,�E�>��0?�V?�0>O��ġZ��>ǁ��"j��>Q�����k��b)��2P>Z�?�)�>�]�>/,��>��KH��Z���ɰ>+�9?�t�����n�X��/��վH�e>�^�>0����"�9A���h���َ����=�NA?]w?;d뽊Z�͸@��;s�M;�=�<�>�i����=�g!>�G���n��^�E6B=w��=U'>n?Ss.>	a�="a�>䐘�y-R��a�>�&F>s0>[�>?hf$?љ#����>��.S%��X>���>�x>wG
>�MI��1�=8��>�b>g�������
�Mm>��S>�gq��5`�Wyk���c=3&�����=7ݘ=�b����:�x�=s7L?cķ�B��'���Us>`�B?ck�>��>K��=Vm�ǣ��rC����?IK@�͎?�2 ���W��4?���?��:���=`N?3��>hi��Қ�$.�>~�@�ل
�\�����G���?ot�?�5��CY��������>U7?�O��w�>�y�IX������u�`�#=���>�<H?�C��]?P��=��~
?/?�Z�{����ȿ}v�Z��>X�?��?��m�<���@��w�>���?wfY?d�i>1^۾�Z��m�>�@?�R?  �>h2�O'���?�Զ?���?gI>��?̝s?k�>U3x�e[/��7��Ֆ��j=aAY;2c�>wR>����cF��Փ�Kg����j�L����a>ͤ$=3�>+N�y6��"@�=5ߋ�4E��z�f�|��>�/q>~�I>�T�>D� ?�b�>{��>�\=nr���ှ.�����L?�(�?,���Wn�.��<u�=??V�ކ?}r4?N�J�I�;�/�>��Z?�A�?�Y?4��>�6�/���c���;贾�$�<}O>���>R}�>ᛡ��JK>h�Ҿ��G���>�&�>D����پg���K�M�4��>i� ?���>���=/t-?�I?��\>�0�>W~J��Z��s�(��}�>���>�;?��?!U?�`���$E��Đ��Ù�Q�5�d�> �m?i3?�>����*��p��<�Gռ#B�<Oׁ?`v?+�X5?D�?a�O?-B?��!> ���N��,��ԟ>�76?��:;C7�5����u�3?uJ�>�F?�d->�A��&�=�K����?x�R?Q�?3��{��9}=~� ;��`=ڥs<�u��cp��^�.>׉<K��=�X>#�:=�`)�%���A��ۇ=R�>�2!>�5������*?j�J��9��/ѕ=�r�ƑD��|>�6K>.¾��]?q�?��{�{����G��#�U��͍?��? ��?�����h���<?B��?�y?qh�>`n���j߾@�޾��r���v�Ȉ�Տ >��>x���,���"���ª��l��k�ȽZ�VY�>�\�>�c?Cf�>�->D�>ﳣ�g�&�v�;����;U�x���C�h�+��/���|������c�J���%�\��>����>�?�I>��M>�!�>��D���>G B>2�r>���>�>��=^8�=�*=�Eн��Y?پr�$��?��t��b?g�q?5�>*o)��P��	���f�=?fw�?v�}?���=�`c�U��w�>Ʀ>��M�"?�n<������7�|�E�dJ���g���=&�~>qC(�HM�S[����x�?��?T�,;�I۾��ͽ\����o=�M�?�(?��)���Q���o���W�S����Ch��k��r�$�Ԟp�f돿.Z�����k�(��7*=��*?/�??����e��~"k�R?�-Vf>x�>��>��>rI>3�	�P�1���]�L'�����G�>T{?։�>i�I?� <?evP?:iL?���>`�>�*���o�>���;���>���>��9?��-?;0?�?s+?�c>r\��� ����ؾ�?8�? F??ί?�����ý�ؗ�ǽg���y�ܖ����=K��<O�׽� u�z�T=��S>�M0? �½2J9��@��0O>��V?c�?���>"���d��r�=��>f��>'с>#� ��Mo��7��J�>��^?� ��Fދ=�>3 0=A�!���*�i�u=N��X�d=��=4����ŻZ��<"7�=��<bIE=�L�:֯���hK���>!X?�y�>*��>����H	�*��-��=�I�=]��>��=	�پ����V���%`� ��>���?(�?�D�=<�>L˵=���[d��
�Ϗ�<>�m)?r�1?�\R?���?��*?��<?��=���r��v�p�+�z�ʐ?V(,?~��>�����ʾw쨿�3�q�?#b?-'a�O���3)��¾Zս¿>T/��%~�����$D��w�����������?3ĝ?;A��6�di����e��Q�C?��>�Y�>W�>�)�l�g����;>+��>�R?���>I?6�g?��K?8>c@�N͹�����o��'��<��,?��^?�˅?{��?���>�7,>�kr��|��~���Z��;�젽�Ϙ�� '���z>��>���>��>k�>	����瓽��X�(�=�2y>��>��`>�#�>s�;>��=ȻG?���>����2<�0	�������<��2v?���?�)?YI=06���F��(��u�>4�?�۪?~_%?ݮI����=!}��M���n��T�>�>�%�>��=� =�">kK�>9�>���̮���8�W;�?2�E?莮=(�ȿ�"�B��=xc��S6>�tJ��������� ��������w��2Q���o���+��e꺾H���[�3�[п�P��>�x�_<	>�>�Ʊ=V��׽P=�]*�q=�M����R�:c�=L�=�U�<�@�=� �+�Y<���Z�?o�I?�=j?�?M�X>B�.>�>x�X+E>� <��-?r�Z>������9{\��Ž�=� ���
�H�����uVR��M>���G(>S]u=`!�����=�>~����m�<��9�H�=�7=�`>�[l<�L>�@
>&j=36w?^���$����4Q��]罁�:?�8�>	|�=@�ƾ+@?�>>�2������0b�.?}��?�T�?�?xsi�ad�>~���掽�p�=����>2>%��=��2�r��>��J>���K�����4�?��@y�??�ዿ��Ͽ�a/>��=d�=��H��X/�Y^W�w�x���u��?��<�'*ž2�g>�f=��ھJӾ��~<�A>��=�ބ�.�Y��8>=�=�ai�=b(D=���>��A>�'|=�ĩ�1��=5�B=s�>��9>D}���VĽ	���<�ك<
e>GQ>	��>[�?]:?m�*?���>9�ܽy��/������>?�=���>�);���>yk?,&h?��??��?hP> %�>,��>�ԓ>���K'�}C��`}�o��>=�?���?'��>&�=s6��� ���G�7E����$?b)?��>>�>�U����,Y&���.�����6��+=�mr�"RU�����Wm�C�㽙�=p�>|��>��>4Ty>B�9>��N>x�>��>K7�<�p�=�ጻ���<1��V��=����)�<�vż����w&��+�ۏ��d�;���;��]<[��;� �=�F�>18>I��>���=�Z���d >�����MM��=��%�A��]b��
~�5*.�J*�*'S>�{o>G��o���X]?��b>��:>n�?��r?��>�2���˾����#[���W����=��=�G�~�:��[c�@H���Ҿ���>�>3�>��l>,�H!?�4x=�⾂^5���>�q��!x�R+��5q�y>����i�UuںB�D?�G�����= ~?!�I?�ߏ?q��>T3��D�ؾ�(0>DL��:=G
�+q�t��5�?�'?K��>��P�D���Ⱦ�H�����>�F+���M��d��1(,�峏�f����>.߰�)%Ѿ�'6��͇�KR����:��N�<��>��K?)�?C�^��胿(@O��b���ֽGR?[@k?��>�?�x?R¨�׾�Rz�  �=h�d?y��?���?��
><�=�g��LX�>O-	?W��?Ͱ�?�Zs?G�?��[�>��;�[ >u���l�=�>��=��=Pi?Y|
?��
?W����	�:��/��\�]����<.��=
��>q�>[�r>�;�=g=�l�=<�[>���>4�>ke>��>"0�>�9Ǿ���U-?�)>Q��>�B8?�l�>6�G=�����=����u.L��8��0�#
��$6�;_]���<���C�>#�ƿ��?�S>J�7?I���n	�ɺO>�g>����>ȽX>�>�n�>���>�� >�ʈ>FW>�FӾ�>����d!��,C���R���Ѿ�{z>����.&����Fy���AI�m���f�j�B.���;=���<H�?����k�0�)�����|�?�[�>�6?�ٌ�)
��X�>T��>ȍ>�I�����Yȍ�Jh�\�?��?Ѝ<>��>� a?�?ހ7�M�.���X���u��B�|^U�_�e�,ቿ#Z������F���_?�+y?�A?�8�</�>�2{?��(������k{>:<0�l�2�g��=Q�>����)-��־���>��	�E>K)f?e|?tF? �*��m��'>��:?Ǜ1?�Ot?��1?h�;?h����$?Io3>�F?�q?+N5?��.?�
?)2>�	�=��V�'=�6���l�ѽ�~ʽ1����3=�^{=bM͸��
<ߐ=Z��<w����ټQ�;�$���%�<:=:�=��=X�R>N/K?��?F�>2
?ޥ
�4������3?F'>��Ǿ�n��s�ݾ^��u�=ke?� �?�Y?@�G>�HT��W����.>�D>$�%>H|>3��>cc���7�ll=�
>���=���=������	���-���>�p>���>V/�>�.>OB�>+ן���Ⱦ��I>��
��)���U"��@��� �.w����H>�$G?lWV?��>��
�5̳��Tc��Z�>-�k?��G?�<?�uN>G�侪kS�I�c�ڻ�=Lݨ<"�(>j*�ꦦ�k��X�=��H�=���>	*��kݠ��Vb>w���q޾��n��J����N�L=�����U=k�I�վ)�9��=}7
>{����� ����\Ҫ��0J?T�j=���#RU�gk���>��>��>~�:�w�G�@�ձ���A�=��>�
;>����2ﾹ|G�m3��8�>�E?Y#_?�7�?���#+s�p�B�� ��	���Ἕ�?(�>�{?DeD>��=����>�dUd��]F�o&�>A��>*h�G�Hў����"�$��ʊ>��?p�>��?LR?� ?��`?�a*?n�?Rď>���(��_�#?R�}?�=����Н>�x7���L��i�>�k?������>G?��?��5?@�_?n??D�=��R�'�输>��>NLP�`���Cd>��M?�?�>�b?@��?}�e>��5��޳��н2O�=  &>��)?�I?I�?�h�>��>B�����=C��>c?�/�?��o?��=��?^:2>���>��=���>���>
?XO?D�s?H�J?��>���<�9���/��UBs���O����;b�H<��y=���2t��C�,��<���;�o���E����񼀺D�����N��;��>�F>2��X=.Aľ^����>�mN��c�lK�����M�Q>���>��>�z>:^@=�W�>R�>��<>q�5�^�S?���>��>�]�;IN{�������W��=�>�/?9\��	�� ��Cjs��P�=�LI?خZ?�v=\���*li?�@A?���Q�9�
%ܾ�� >3怾��d?�,?�a�����><�e?�a?���>5j��pq�15����P�߇-��|{=w��>��i�S��R[>Py�>rB�>e@>�TO>��!��5M�I��ō�>��?%_�?��?Ig>r�����n���A��+^?̃�>jE����"?���Z�ϾgT��s��'⾛���&��UK���t��n�$�"ԃ�׽�¼=N�?(s?.Yq?��_?1� ���c��/^�O
���oV��!�� ���E�-$E�+�C�(�n��e��#�������G=E�_��-�B�??	?����˩>�����f��Ⱦ:��=􌣾���i`=aS<�*�=�-:>G�F��B�^��"?�%�>�t�>0�%?U�^���@��7�ɸL�;���G����>�l>�?��V>3
�=�����.�xo����мZ+v>zc?^�K?�n?�l��&1�˄��Ϛ!��/�A^��v�B>�b>巉>߲W���r:&�sZ>���r�?���u���	�`~=��2?
+�>t��>NM�?��?z	�f��1fx���1��Q�<�.�>�i?(@�>��>�Ͻ�� ���>Z�l?D��>�>�����Z!�V�{�͟ʽ-#�>;�>Ҹ�>]�o>��,�� \�j��|���s9��Y�= �h?T�����`��>�R?`��:O�G<Jx�>��v�տ!�~���'�#�>�{?䊪=��;>��ž"%��{��6��A)?5~?Ǜ���>(���>�J?��>`Ʀ>nt�? s�><�þ��ڼh&?�Ga?+�O?�U@?���>-�=y������F&��s"=��>�KV>;_c=�7�=h��N�(��!`@=��=��3eԽ�;�;�~8�?S�<a�<}-)>���8?��;a�*��e��j�vg���=u$��p.���Ⱦ`ѕ�h���28�O�S�R���˚$�Dv{���m�<��?\��?�摾�v�;W��\�e�Q���!�>�;����;�e��S����H����Ǿ�ľ��6�^�Z��<_�M�4��'?�����ǿ򰡿�9ܾk! ?�A ?�y?�m�"��8��� >V�<$�����X�����οe��� �^?w��>0�0����>���>��X>�Dq>����螾�R�<�?�-?��>݋r�ʕɿ���<���?��@�/?����� ��
��?ej�>8��>����^�^�g�ʽo�>�C�?��?6�W=6�i�f�սk��?5&+<����Z�=�ި>R>z�����x=�P�>��q��m��	���g7�>f�>��z�]�����*���c>�hV>�!¾)!���?�_V���d��/,��`z�6�=�Q?ʰ�> K�=��&?XE�N�οc�[��_?��?���?� &?SZ��j6�>p�ھu�H?��9?��>+*�F�q��A>6���}?��Y)׾��U�QH�=��>dk>b�:����po;�ޗ���9�=���qgſ�#���"�z�<kcJ�{yp�чɽa�����E�l���g�p����GL=+A�=��M>	e�>%�T>�S>o�W?��j?TW�>U�>3�ٽӨ��^lѾ�|�:�1��j�(�'������:Ϣ��!���߾��
��n����D�ƾ�FC��h�=
NP�5����!��b� G�!�1?Я,>�˾�M���<�˾Q)��M����߹�݈Ǿ\w/�Z	l�� �?��A?���HQT�_��)���/Z۽��U?п
�:$��l��b)�=:Ъ���=�P�>;@{=��x�2��OM�/�0?�?2�þ/�����(>����)=�V*?μ?�f};���>��?��8�ܯ��pă>u�`>�e�>�}�>@�>$���h�̽Q{"?§P?�h#������>��վ�ރ�p��=QL�=\W+��7C��>>�
ջ5|���<R�U�LA�;�Mh?梈>�X����U���k�J>]	�>�k?[|?�R�>T��?��L?�ɇ=%	��c��]>����=9Ep?TW?�O�=K.��Y\��g�U�Y�?���?5&3>*.��]ھ=I��ڍ�x�4? �q?X�?���^c��1���96�@P?��v?q^�}s������V�O5�>�X�>��>��9��h�>:�>?�	#��F��+���X4��?J�@I��?�v;<�7�*��=�;?z]�>ХO��>ƾW���䀵���q=�&�>+���{ev����Y,�x�8?Ҟ�?0��>��������=3ȕ�{Y�?+�?3}���a<����6l�Wk��\�<8x�=����!����7��ƾ�
�=q��{=��F��>�P@�(��0�>|p8�L*�oIϿ���isо��q���?oA�>�Fǽ%-���yj�h@u���G�a�H��{��q6h>�s%=�@	��s��g{���I�����&�?���=N�?>$���(ؾ+�ԾO�@=Qn�>#?���>�-&=�s����?e�u�ο��?����{J?C��?�rq?�D�>��.�����Z=��Gx	>f�k?"ȏ?� Y?sѽ�y��&�ϽB�j?_���T`���4�=HE�A U>&#3?�D�>ǒ-���|=�>S��>�i>~#/�I�Ŀ�ٶ��������?���?�n����>���?r+?5i�x7��L\��m�*��'�;<A?32>W���ʸ!��.=�{ϒ���
?�|0?/}��.���B?�|]�zq���.���+�g
N>͍�2n=��<<�_�� kf�	#����G�ag�?,��?"%�?3mE����583?���>Ջ�b���e�;4�>���>��h>�
��m�=�>�g[�7ݤ=n��?a�?�*(?�ϛ��𵿈�W=a?~B�>	@�?�-�>G�#?�]N�$ؾlX�=��">�:�=˒>�:
?Ǆ2?��>m�=��z��W$��)P��0d��L��P����>2�E?t�v?�;>�m���@ǽ�5�\���MZ���ͽEo���p�5�6��"X=.�<�pv=��n�������?Op�5�ؿ�i��p'��54?��>�?����t�%���;_?Rz�>�6��+���%���B�^��?�G�??�?��׾kR̼�>:�>�I�>2�Խ����V�����7>.�B?N��D��r�o�o�>���?
�@�ծ?li�\$?F� ���}��E��	C���=��8?߰ᾼ�o>{^�>��=TWx��Ũ�&t��y�>[.�?���?���>7n?��n��MC���^=5��>�xd?�a?���;�_��XE>ma?���t��v
���i?d@@OTa?r����p县"q������������AK>
��8>2��=�ּ�4���i{=�[>%N[>#HX>3u>g�:>]�>�V��t�������^�P���"����C�˽�־Nb�9���ͪ�ZF;58�����ԫ����m@3�U���6�=h�U?�2R?�\p?�U ?��v��>����^�=��"�Ii�=W�>R2?�@L?�K*?��=���&e��P���<��X������>�sH>�a�>���>+̭>g����J>=?>�h�>=- >�j$=Y`��j=�	O>��>r��>�f�>�C<>��>Dϴ��1��k�h��
w��̽1�?y���S�J��1���9��Ԧ���h�=Eb.?|>���?пc����2H?$���w)��+���>z�0?�cW?�>��\�T�4:>9����j�6`>�+ �tl���)��%Q>xl?ALl>P�|>�:1��7��P��d����>,7?����+��Jq���G��m۾��N>.��>�?��	���ܰ~���s����=Z?<?o�?*���ڶ�^5w�Qs���?H>�3a>�L=�ţ=SKH>7xd�6ܽ�/G���8=�y�=��a>e?��.>Sȩ=�>�����
R�d��>0l.>- >8@?�]?C�$���ǽ���)��>�i�>�܀>���=CQ����=g��>��t>����흽 ��"�G� [>K�F�``S�[��c=\���݆�=Lmq=>V��rv+�1=�[?�4��8%�������x>�K?V��>m_9>n�=��辳լ��Zо�8�?6�@vВ?ih#���\���0?�?a���}����� ?;��>��&>� ��Z>����������,o�����?K��?��m���y��*�>ILA?�="��g�>Bx�FZ�������u�6�#=���>�8H?�U����O�=>��v
?�?_�ϩ����ȿ�{v����>-�?���?9�m�_A���@����>��?�fY?�ni>Ig۾^`Z�*��>��@?�R?��>�9�<�'��?�޶?�?.I>��?�s?�{�> Xx��W/��1������_=�&_;)f�>WW>����VeF�|֓�g��8�j���E�a>Ro$=�>�?佀5��).�=�ϋ�hG��Bg� ��>�'q>��I>jN�>�� ?�W�>��>%�=�b��h‾ﶖ�%P?��?k���^��墽��>s�ü�v?mNW?�y�=\sj� �>��A?�k?]�S?L�>����������;u7>�ߞ>SL�>���>q)�� d<>�ž�����>
�R>-��RGپ	�U�����N�>-�%?�W�>P#=
`!?ZN#?��i>��>�E�����@B��l�>̬�>�?�.�?m?�ݹ��54�I����i��gAX��X>QAw?��?S(�>'9���R��+�
��7)�ϊ��͂?f?fX�R�?��?��@?�A?@ia>Ϫ���׾�@����>�"?<�i��m?��_�Vv=A��>1L>�?��=@˂�}�ή�P��M��h2D? u�?kw!?����Y*�d�=,�^=�#����ڼ�Dr����e3O=�P�>c��=
QQ>��]>�ր=�W�w|��Y9F���<��>�f`>;훾.���d)?^+�����o��=��o���F��zx>��;>}�ƾƖ[?%�N��x����������T� �?I[�?�ĕ?��ĽULg��=?���?�A?Ƿ�>(}���ݾ$�ܾ=m��)b�����=�!�>��ռ�E���r먿#�������,5��U�>�>҈?ޠ?���=�:�>+�x3��U������LJ�`���W=�:�-��U�o"8��P��]�仾˷��.��>ɏ����>'?a!>^
�>��>�u=��>�>4*W>Pڲ>ٗ >�e>d?�=�Eu=�6�;F�S?�þ��$�:�����"�G?u�]?�u�>�uq�bV��U�Ծ�*?�Ǝ?r)�?�CL>�cV���&�R�>���>�1��}4?'�˼����]��<�ؾ�*Q�t����)=��>���ڒL��K�eH�I�?��?|��;	̾�J�<���6 m= �?�5(?g�)�T�Q��;p��W���R�6��F�h��%��a�$�qp��揿T���~��m�(��S2=Z�*?RĈ?�6����p¬�Ҫj���?�ۀd>���>��>r�>��H>��	�B|1��^�n�&�M���D�>��{?L��>[�I?6�;?�uP?ojL?$��>\^�>5��e�>���;z��>%��>��9?��-?�70?�y?ts+?^7c>3n�� ��T�ؾ0?��?kI?5?��?Cڅ�;jý�,��|�f���y�a����=*�<\�׽*Au��T=�T>(�%?����'�z��RB>��h?�?�	�>pbH���оJ#�=���>ۡ?�^E>3P�i����(��S�>�Ȋ?h/4�&��<_ �=�%R=v]��==t�:��=��!>w%[�zX��ͽ"T�=���=��=渂<I��fj�8���F�?��	?��?a�>P�������$5�|}�|�g>�?^+>�Qɾ�=��!����ZD��C�>+�?
m�?C�F�%�o>	�N>F��W'�� �B����W@>*�O?^J?��K?���? E?��K?��a>�
�����fF?��0m��?!,?)��>~���ʾ���3���?]?m2a����46)�ϐ¾��Խ��>MX/�x(~����dD�^������Y�����?g��?�A��6��y�龘�
d���C?��>_W�>w�>4�)�d�g�C%�/;>ǌ�>6R?dw�>�]>?\T?�?O?u�D>z�D�Gɪ�������leýW&-?"W?L��?�)�?<�?e�/>���췟�����H8;0Ž.�Ⱦҋ�=yZt>Tq�>�ͯ>o�>���=����ʬ��K��R��=�ʔ>�z�>Lb[>ǹ�><�f>uu�= �G?���>!M���{�褾�����8��ku?*z�?�+?�=ڜ���E�d���|�>�T�?\׫?�"*?��R�&�=��ּ�����Yr�$ҷ>"ʹ>ܖ�>@Ñ=\�C=��>9�>���>@��YH��m8���N���?F?Ԟ�=��Ͽ�m�bRk�f�����t|��EYr�Y:��Tc �O��=➾�T �«����m��+��|�����ؕ��t,���| ?$v�=�3�=M��=ے=&'����=��Q;B=�������<�wN���������%��I
;� ==?~�^��z<�?'�w?�n�?;��>ʒ�>��=�Ӳ���=�>O�3?���2�RJ�!$��3{߾�g����^�ɰ����c�!���]s�|w�tЕ>NI�>��|�@��<��>5hx�|�=U���̒�]�<�1�=,�=`�*>�VY>�@>Y0w?ܚ��5����3Q�o~�i�:?T2�>���=�rƾ/@?w�>>�2�����\��+?=��?�S�?#�?�`i��o�>���"���b�=����M2>�>�=2�2����>V�J>݂��H���;��/6�?2�@'�??�⋿�Ͽ\/>�|>m)>�V�p*���N��N���h�.�?�LA���I�'>�p�=p޾�ؾ��<[}E>6�>������W�*�=������=�^�=P��>V�N>d�=�䃽���=���=̟>]x!>�jd�o���E��[1{���a="{d>��<>_�>ǟ?L�(?�`?7�>ޭu��dھ'�þ�X�>�`�=t��>޶+=&�I>u
�>�d@?�A?aEA?7=�>�=�!�>:p�>�)�C-m��,ܾn����(�<UT�?姇?c�>�)����V�����}9�(V���?�
-?�?	�>C.�*߿��$���1�Y峽@�7�2\=�db��.�X�Լ(�����y�=�@�>�>�>g�><�>�7>.�G>�[�>?�>�ڷ<�w=��0�%��<r��㟛=����MT<D; ���U;, ��}~-��Ǽ�F��@��:�)U<��;��=���>��>��>�k�=U���(>슙��KM�T^�=J����A�sc�jC~���.���2�X)K>_c]>UX��}���?��`>��F>w��?9�t?Pa>�C
�/&Ӿ�ڛ�
�Y�'�R��=�u>�dB���;���_�C L�r�;���>h��>��>f�l>�,�N#?���w=�⾼a5�^�>�{��n��)�29q��?������<i��FӺ?�D?�F�����=K"~?�I?$�?��>���m�ؾ�50>�H����=���)q��i���?'?ݖ�>]��D�w�����a�>�6��J����������=���=@:>������ǾE�E��w�3P����.�e�d�J:�>�Mu?#$�?�˞�)s`�d�����f��Dt?�F?n��>�v?��>�O��y�9�	�&�>M��?�(�?�l�?�t�=�k�=�b��D �>-%	?_��?l��?&s?��?����>��;+� >GW��=��={7>�^�=�#�=�n?��
?X�
?Ü��	����~<�m^�2��<!��=5S�>ω>��q>X��=��h=4�=#]>��>�K�>��d>{/�>���>�h��f���"?\�=i�>?>?6f>��l:��$��u�=!
u�`�߽a�T���u*��Y�=Z�=&+=>T�k<�i�>tռ��>�?��=�����?|�p�Ž'��>�=�9�����>(RN>}d�>���>5�>D��=���>Ă}>|����=�p��@�{�B��P�#{���>��_�8ċ�����˽C.u��r��R�+���\}v��T5�\o�=�?Y����I�cf�y���w�?�͆=�?�&��3�����#>Յ�>0�B>��۾<9��3z����b�l?��?�c>��>�Z?��?+�1���1�ֈV�d�w���A�܊_���`�Dċ�]w��w���-���`?U$x?"B?�X�<�wx>�G~?��Շ��I�>\�.��&9�w�<p�>A߰�F�Y��ξ����}����I>xAj?e�?��?�*R��n��+'>��:?9�1?�Qt?h2?<�;?<��:�$?Jp3>�H?g?wH5?_�.?�
?�2>���=O���3�'=7?����'�ѽ�pʽc��3=q*{=l��7�y<jd=�x�<�z�Q�ؼ��;�=���Z�<�T:=��=S��=�o�>�:L?�T�>pl�>��$?G��?[&�� ܾ�e?���=�2��Q����۾��'��=Y\h?�U�?��W?B ,>I�� �c`>��>&�">ֹB>~u�>P��J��jx�=w_6>�=>�D=��ƽ������V傾�+{=��>���>�>9hV=<�">�`���ƕ��T�>�}��������2���:�!�6�^�վ�.b>��;?��T?�>�������EW���?�^g?��V?rH*?�J�=8���zQ��o���[=��=>(>B�&�=e���ߞ��z*���=N��>7���kݠ��Vb>w���q޾��n��J����N�L=�����U=k�I�վ)�9��=}7
>{����� ����\Ҫ��0J?T�j=���#RU�gk���>��>��>~�:�w�G�@�ձ���A�=��>�
;>����2ﾹ|G�m3��8�>�E?Y#_?�7�?���#+s�p�B�� ��	���Ἕ�?(�>�{?DeD>��=����>�dUd��]F�o&�>A��>*h�G�Hў����"�$��ʊ>��?p�>��?LR?� ?��`?�a*?n�?Rď>���(��_�#?R�}?�=����Н>�x7���L��i�>�k?������>G?��?��5?@�_?n??D�=��R�'�输>��>NLP�`���Cd>��M?�?�>�b?@��?}�e>��5��޳��н2O�=  &>��)?�I?I�?�h�>��>B�����=C��>c?�/�?��o?��=��?^:2>���>��=���>���>
?XO?D�s?H�J?��>���<�9���/��UBs���O����;b�H<��y=���2t��C�,��<���;�o���E����񼀺D�����N��;��>�F>2��X=.Aľ^����>�mN��c�lK�����M�Q>���>��>�z>:^@=�W�>R�>��<>q�5�^�S?���>��>�]�;IN{�������W��=�>�/?9\��	�� ��Cjs��P�=�LI?خZ?�v=\���*li?�@A?���Q�9�
%ܾ�� >3怾��d?�,?�a�����><�e?�a?���>5j��pq�15����P�߇-��|{=w��>��i�S��R[>Py�>rB�>e@>�TO>��!��5M�I��ō�>��?%_�?��?Ig>r�����n���A��+^?̃�>jE����"?���Z�ϾgT��s��'⾛���&��UK���t��n�$�"ԃ�׽�¼=N�?(s?.Yq?��_?1� ���c��/^�O
���oV��!�� ���E�-$E�+�C�(�n��e��#�������G=E�_��-�B�??	?����˩>�����f��Ⱦ:��=􌣾���i`=aS<�*�=�-:>G�F��B�^��"?�%�>�t�>0�%?U�^���@��7�ɸL�;���G����>�l>�?��V>3
�=�����.�xo����мZ+v>zc?^�K?�n?�l��&1�˄��Ϛ!��/�A^��v�B>�b>巉>߲W���r:&�sZ>���r�?���u���	�`~=��2?
+�>t��>NM�?��?z	�f��1fx���1��Q�<�.�>�i?(@�>��>�Ͻ�� ���>Z�l?D��>�>�����Z!�V�{�͟ʽ-#�>;�>Ҹ�>]�o>��,�� \�j��|���s9��Y�= �h?T�����`��>�R?`��:O�G<Jx�>��v�տ!�~���'�#�>�{?䊪=��;>��ž"%��{��6��A)?5~?Ǜ���>(���>�J?��>`Ʀ>nt�? s�><�þ��ڼh&?�Ga?+�O?�U@?���>-�=y������F&��s"=��>�KV>;_c=�7�=h��N�(��!`@=��=��3eԽ�;�;�~8�?S�<a�<}-)>���8?��;a�*��e��j�vg���=u$��p.���Ⱦ`ѕ�h���28�O�S�R���˚$�Dv{���m�<��?\��?�摾�v�;W��\�e�Q���!�>�;����;�e��S����H����Ǿ�ľ��6�^�Z��<_�M�4��'?�����ǿ򰡿�9ܾk! ?�A ?�y?�m�"��8��� >V�<$�����X�����οe��� �^?w��>0�0����>���>��X>�Dq>����螾�R�<�?�-?��>݋r�ʕɿ���<���?��@�/?����� ��
��?ej�>8��>����^�^�g�ʽo�>�C�?��?6�W=6�i�f�սk��?5&+<����Z�=�ި>R>z�����x=�P�>��q��m��	���g7�>f�>��z�]�����*���c>�hV>�!¾)!���?�_V���d��/,��`z�6�=�Q?ʰ�> K�=��&?XE�N�οc�[��_?��?���?� &?SZ��j6�>p�ھu�H?��9?��>+*�F�q��A>6���}?��Y)׾��U�QH�=��>dk>b�:����po;�ޗ���9�=���qgſ�#���"�z�<kcJ�{yp�чɽa�����E�l���g�p����GL=+A�=��M>	e�>%�T>�S>o�W?��j?TW�>U�>3�ٽӨ��^lѾ�|�:�1��j�(�'������:Ϣ��!���߾��
��n����D�ƾ�FC��h�=
NP�5����!��b� G�!�1?Я,>�˾�M���<�˾Q)��M����߹�݈Ǿ\w/�Z	l�� �?��A?���HQT�_��)���/Z۽��U?п
�:$��l��b)�=:Ъ���=�P�>;@{=��x�2��OM�/�0?�?2�þ/�����(>����)=�V*?μ?�f};���>��?��8�ܯ��pă>u�`>�e�>�}�>@�>$���h�̽Q{"?§P?�h#������>��վ�ރ�p��=QL�=\W+��7C��>>�
ջ5|���<R�U�LA�;�Mh?梈>�X����U���k�J>]	�>�k?[|?�R�>T��?��L?�ɇ=%	��c��]>����=9Ep?TW?�O�=K.��Y\��g�U�Y�?���?5&3>*.��]ھ=I��ڍ�x�4? �q?X�?���^c��1���96�@P?��v?q^�}s������V�O5�>�X�>��>��9��h�>:�>?�	#��F��+���X4��?J�@I��?�v;<�7�*��=�;?z]�>ХO��>ƾW���䀵���q=�&�>+���{ev����Y,�x�8?Ҟ�?0��>��������=3ȕ�{Y�?+�?3}���a<����6l�Wk��\�<8x�=����!����7��ƾ�
�=q��{=��F��>�P@�(��0�>|p8�L*�oIϿ���isо��q���?oA�>�Fǽ%-���yj�h@u���G�a�H��{��q6h>�s%=�@	��s��g{���I�����&�?���=N�?>$���(ؾ+�ԾO�@=Qn�>#?���>�-&=�s����?e�u�ο��?����{J?C��?�rq?�D�>��.�����Z=��Gx	>f�k?"ȏ?� Y?sѽ�y��&�ϽB�j?_���T`���4�=HE�A U>&#3?�D�>ǒ-���|=�>S��>�i>~#/�I�Ŀ�ٶ��������?���?�n����>���?r+?5i�x7��L\��m�*��'�;<A?32>W���ʸ!��.=�{ϒ���
?�|0?/}��.���B?�|]�zq���.���+�g
N>͍�2n=��<<�_�� kf�	#����G�ag�?,��?"%�?3mE����583?���>Ջ�b���e�;4�>���>��h>�
��m�=�>�g[�7ݤ=n��?a�?�*(?�ϛ��𵿈�W=a?~B�>	@�?�-�>G�#?�]N�$ؾlX�=��">�:�=˒>�:
?Ǆ2?��>m�=��z��W$��)P��0d��L��P����>2�E?t�v?�;>�m���@ǽ�5�\���MZ���ͽEo���p�5�6��"X=.�<�pv=��n�������?Op�5�ؿ�i��p'��54?��>�?����t�%���;_?Rz�>�6��+���%���B�^��?�G�??�?��׾kR̼�>:�>�I�>2�Խ����V�����7>.�B?N��D��r�o�o�>���?
�@�ծ?li�\$?F� ���}��E��	C���=��8?߰ᾼ�o>{^�>��=TWx��Ũ�&t��y�>[.�?���?���>7n?��n��MC���^=5��>�xd?�a?���;�_��XE>ma?���t��v
���i?d@@OTa?r����p县"q������������AK>
��8>2��=�ּ�4���i{=�[>%N[>#HX>3u>g�:>]�>�V��t�������^�P���"����C�˽�־Nb�9���ͪ�ZF;58�����ԫ����m@3�U���6�=h�U?�2R?�\p?�U ?��v��>����^�=��"�Ii�=W�>R2?�@L?�K*?��=���&e��P���<��X������>�sH>�a�>���>+̭>g����J>=?>�h�>=- >�j$=Y`��j=�	O>��>r��>�f�>�C<>��>Dϴ��1��k�h��
w��̽1�?y���S�J��1���9��Ԧ���h�=Eb.?|>���?пc����2H?$���w)��+���>z�0?�cW?�>��\�T�4:>9����j�6`>�+ �tl���)��%Q>xl?ALl>P�|>�:1��7��P��d����>,7?����+��Jq���G��m۾��N>.��>�?��	���ܰ~���s����=Z?<?o�?*���ڶ�^5w�Qs���?H>�3a>�L=�ţ=SKH>7xd�6ܽ�/G���8=�y�=��a>e?��.>Sȩ=�>�����
R�d��>0l.>- >8@?�]?C�$���ǽ���)��>�i�>�܀>���=CQ����=g��>��t>����흽 ��"�G� [>K�F�``S�[��c=\���݆�=Lmq=>V��rv+�1=�[?�4��8%�������x>�K?V��>m_9>n�=��辳լ��Zо�8�?6�@vВ?ih#���\���0?�?a���}����� ?;��>��&>� ��Z>����������,o�����?K��?��m���y��*�>ILA?�="��g�>Bx�FZ�������u�6�#=���>�8H?�U����O�=>��v
?�?_�ϩ����ȿ�{v����>-�?���?9�m�_A���@����>��?�fY?�ni>Ig۾^`Z�*��>��@?�R?��>�9�<�'��?�޶?�?.I>��?�s?�{�> Xx��W/��1������_=�&_;)f�>WW>����VeF�|֓�g��8�j���E�a>Ro$=�>�?佀5��).�=�ϋ�hG��Bg� ��>�'q>��I>jN�>�� ?�W�>��>%�=�b��h‾ﶖ�%P?��?k���^��墽��>s�ü�v?mNW?�y�=\sj� �>��A?�k?]�S?L�>����������;u7>�ߞ>SL�>���>q)�� d<>�ž�����>
�R>-��RGپ	�U�����N�>-�%?�W�>P#=
`!?ZN#?��i>��>�E�����@B��l�>̬�>�?�.�?m?�ݹ��54�I����i��gAX��X>QAw?��?S(�>'9���R��+�
��7)�ϊ��͂?f?fX�R�?��?��@?�A?@ia>Ϫ���׾�@����>�"?<�i��m?��_�Vv=A��>1L>�?��=@˂�}�ή�P��M��h2D? u�?kw!?����Y*�d�=,�^=�#����ڼ�Dr����e3O=�P�>c��=
QQ>��]>�ր=�W�w|��Y9F���<��>�f`>;훾.���d)?^+�����o��=��o���F��zx>��;>}�ƾƖ[?%�N��x����������T� �?I[�?�ĕ?��ĽULg��=?���?�A?Ƿ�>(}���ݾ$�ܾ=m��)b�����=�!�>��ռ�E���r먿#�������,5��U�>�>҈?ޠ?���=�:�>+�x3��U������LJ�`���W=�:�-��U�o"8��P��]�仾˷��.��>ɏ����>'?a!>^
�>��>�u=��>�>4*W>Pڲ>ٗ >�e>d?�=�Eu=�6�;F�S?�þ��$�:�����"�G?u�]?�u�>�uq�bV��U�Ծ�*?�Ǝ?r)�?�CL>�cV���&�R�>���>�1��}4?'�˼����]��<�ؾ�*Q�t����)=��>���ڒL��K�eH�I�?��?|��;	̾�J�<���6 m= �?�5(?g�)�T�Q��;p��W���R�6��F�h��%��a�$�qp��揿T���~��m�(��S2=Z�*?RĈ?�6����p¬�Ҫj���?�ۀd>���>��>r�>��H>��	�B|1��^�n�&�M���D�>��{?L��>[�I?6�;?�uP?ojL?$��>\^�>5��e�>���;z��>%��>��9?��-?�70?�y?ts+?^7c>3n�� ��T�ؾ0?��?kI?5?��?Cڅ�;jý�,��|�f���y�a����=*�<\�׽*Au��T=�T>(�%?����'�z��RB>��h?�?�	�>pbH���оJ#�=���>ۡ?�^E>3P�i����(��S�>�Ȋ?h/4�&��<_ �=�%R=v]��==t�:��=��!>w%[�zX��ͽ"T�=���=��=渂<I��fj�8���F�?��	?��?a�>P�������$5�|}�|�g>�?^+>�Qɾ�=��!����ZD��C�>+�?
m�?C�F�%�o>	�N>F��W'�� �B����W@>*�O?^J?��K?���? E?��K?��a>�
�����fF?��0m��?!,?)��>~���ʾ���3���?]?m2a����46)�ϐ¾��Խ��>MX/�x(~����dD�^������Y�����?g��?�A��6��y�龘�
d���C?��>_W�>w�>4�)�d�g�C%�/;>ǌ�>6R?dw�>�]>?\T?�?O?u�D>z�D�Gɪ�������leýW&-?"W?L��?�)�?<�?e�/>���췟�����H8;0Ž.�Ⱦҋ�=yZt>Tq�>�ͯ>o�>���=����ʬ��K��R��=�ʔ>�z�>Lb[>ǹ�><�f>uu�= �G?���>!M���{�褾�����8��ku?*z�?�+?�=ڜ���E�d���|�>�T�?\׫?�"*?��R�&�=��ּ�����Yr�$ҷ>"ʹ>ܖ�>@Ñ=\�C=��>9�>���>@��YH��m8���N���?F?Ԟ�=��Ͽ�m�bRk�f�����t|��EYr�Y:��Tc �O��=➾�T �«����m��+��|�����ؕ��t,���| ?$v�=�3�=M��=ے=&'����=��Q;B=�������<�wN���������%��I
;� ==?~�^��z<�?'�w?�n�?;��>ʒ�>��=�Ӳ���=�>O�3?���2�RJ�!$��3{߾�g����^�ɰ����c�!���]s�|w�tЕ>NI�>��|�@��<��>5hx�|�=U���̒�]�<�1�=,�=`�*>�VY>�@>Y0w?ܚ��5����3Q�o~�i�:?T2�>���=�rƾ/@?w�>>�2�����\��+?=��?�S�?#�?�`i��o�>���"���b�=����M2>�>�=2�2����>V�J>݂��H���;��/6�?2�@'�??�⋿�Ͽ\/>�|>m)>�V�p*���N��N���h�.�?�LA���I�'>�p�=p޾�ؾ��<[}E>6�>������W�*�=������=�^�=P��>V�N>d�=�䃽���=���=̟>]x!>�jd�o���E��[1{���a="{d>��<>_�>ǟ?L�(?�`?7�>ޭu��dھ'�þ�X�>�`�=t��>޶+=&�I>u
�>�d@?�A?aEA?7=�>�=�!�>:p�>�)�C-m��,ܾn����(�<UT�?姇?c�>�)����V�����}9�(V���?�
-?�?	�>C.�*߿��$���1�Y峽@�7�2\=�db��.�X�Լ(�����y�=�@�>�>�>g�><�>�7>.�G>�[�>?�>�ڷ<�w=��0�%��<r��㟛=����MT<D; ���U;, ��}~-��Ǽ�F��@��:�)U<��;��=���>��>��>�k�=U���(>슙��KM�T^�=J����A�sc�jC~���.���2�X)K>_c]>UX��}���?��`>��F>w��?9�t?Pa>�C
�/&Ӿ�ڛ�
�Y�'�R��=�u>�dB���;���_�C L�r�;���>h��>��>f�l>�,�N#?���w=�⾼a5�^�>�{��n��)�29q��?������<i��FӺ?�D?�F�����=K"~?�I?$�?��>���m�ؾ�50>�H����=���)q��i���?'?ݖ�>]��D�w�����a�>�6��J����������=���=@:>������ǾE�E��w�3P����.�e�d�J:�>�Mu?#$�?�˞�)s`�d�����f��Dt?�F?n��>�v?��>�O��y�9�	�&�>M��?�(�?�l�?�t�=�k�=�b��D �>-%	?_��?l��?&s?��?����>��;+� >GW��=��={7>�^�=�#�=�n?��
?X�
?Ü��	����~<�m^�2��<!��=5S�>ω>��q>X��=��h=4�=#]>��>�K�>��d>{/�>���>�h��f���"?\�=i�>?>?6f>��l:��$��u�=!
u�`�߽a�T���u*��Y�=Z�=&+=>T�k<�i�>tռ��>�?��=�����?|�p�Ž'��>�=�9�����>(RN>}d�>���>5�>D��=���>Ă}>|����=�p��@�{�B��P�#{���>��_�8ċ�����˽C.u��r��R�+���\}v��T5�\o�=�?Y����I�cf�y���w�?�͆=�?�&��3�����#>Յ�>0�B>��۾<9��3z����b�l?��?�c>��>�Z?��?+�1���1�ֈV�d�w���A�܊_���`�Dċ�]w��w���-���`?U$x?"B?�X�<�wx>�G~?��Շ��I�>\�.��&9�w�<p�>A߰�F�Y��ξ����}����I>xAj?e�?��?�*R��n��+'>��:?9�1?�Qt?h2?<�;?<��:�$?Jp3>�H?g?wH5?_�.?�
?�2>���=O���3�'=7?����'�ѽ�pʽc��3=q*{=l��7�y<jd=�x�<�z�Q�ؼ��;�=���Z�<�T:=��=S��=�o�>�:L?�T�>pl�>��$?G��?[&�� ܾ�e?���=�2��Q����۾��'��=Y\h?�U�?��W?B ,>I�� �c`>��>&�">ֹB>~u�>P��J��jx�=w_6>�=>�D=��ƽ������V傾�+{=��>���>�>9hV=<�">�`���ƕ��T�>�}��������2���:�!�6�^�վ�.b>��;?��T?�>�������EW���?�^g?��V?rH*?�J�=8���zQ��o���[=��=>(>B�&�=e���ߞ��z*���=N��>7����ǫ�5�b>���G���Nk�2�J�]�վ�i�=+�L��=r~�h�;�t���%�=*�>�з�����֔�Z����J?��=H���\(M�����)�=Rkr>L��>�����zQ�^�;�G����Xw=�f�>/>��ܼ2���yB����І>��D?#Q_?n��?�4��7nr�cC�5��X��a���?J)�>��?�D>�ֵ=�Q���:��b��"E��>�>i!�>S���fG�����gZ��`�$��Ë>�:?�>��?��P??m�b?)U,?0b?��>� ��?k���?X$?�d=�/�"�o�06�F�Z�Cb�>��?-���g+|>���>0�$?@�R?^�q?Ii�>;�8��Ⱦ�3�<M�>�[�>ˬT�������>��G?��>n�@?�Q�?�_�>t�-�	�����	S�=��4>��?M�?�a�>{��>;��>9���H �=��>=c?a0�?w�o?���=<�?82>��>E��=���>}��>�?XO?��s?��J?#��>伍<�:��_;���Cs�)�O�f��;�pH<l�y=d��/1t��J�
��<+ѳ;�y���H��Y�񼂺D������;�n�>�)9>��M��:>��߾��i��w�=I�k��m���-��!ᠾ]
%>䢯>�G�>��>*ꈽ�H>9_�>��>��2��[?)��>�j�>$�_=��k��E���0�a�>�,?�;�ޜ���8���	c� ��=��Y?Z�K?D��=�t�hTm?=�6?q$�z�)�[ܾ�=?���X??*'?e՛����>лt?VP?]��>Ƞ�!�{�Yq��|gi�9�S�w=R��>�����8���>+u?�>��>]Lo>�ۺ���[��|��I۸>C��?&z�?�a�?�uk>�p���꿿O��7���^?���>e����"?�$��?�Ͼ�*�������p�����D(���z���$��ԃ���׽d�=��?�s??]q?��_?ܢ ��c�?^�����aV�)����E��E� �C�^�n��_�!�����I]H=0�~�2�@�ri�?p�'?��0��r�>����W�񾍤;��B>*tz�sS�=�@���#<=��Z=�e�K,�@%��?�?j��> ��>dH<?�r[��#>���1�Y�7�������2>���>{,�>�y�>���;��)��ὡNȾ�t��I нAv>�|c?�K?��n?_���#1�����!�sV/��d����B>*�>#��>g�W� ���:&�>^>���r�J������E�	�L�~=/�2?��>
��>�H�?\�?Xt	��z���Gx�}1�^�<m#�>6i?o3�>}چ>�Ͻ�� �̨�>�l?�c�>)l�>����!�}({�#wҽ���>��>�x�>�o>�/-��d\��A��s��p8�ĵ�=s�g?0R��-�a�n�>��Q?�z;[�<zK�>d;z��k!�	��J#��r>��?4g�=6�9>�ž�r�%�{����i�!?��?!۝���0����>�B?c�>�^�>�t|?��M>Rƾ�h���	?�j?��e?M;?u׼>�4V���=̕���nJ�2lZ���o>"j.>T�K=��=�9��:�8�����:=U�=$����R�e��;U�P=0О=sy���-$>Kg޿G�=��F�� >��N־M�⾇0����ݵ�A�$=��d� �t���W�o�P����X8���|u����?���?)�پ������2���7ӾE��>U��`y�W0��dɽ�Œ�DMa� ���_�:�,�	�]�i�?��b'?����ǿn���#ܾ��?q ?��y?� ��l"�(u8��!>�n�<P����T����ο����G�^?U��>v�v���P�>u˂>_X>3p>���U������<\�?��-?<J�>�s���ɿ~���&�<e��?t�@�H?} t����1�=� ?�.?�ʹ>Vo�� �4������c>�*�?ι?ϯE=�KC��G���K�?Q��=��l��^�<�m>�"d>��˻�����>�>M����p�^CL����>:��>3����쎾��.�+8>���>b���
aA��΄?0_\��f��/��>��!�>W�T?�>j��=��,?yH��xϿi�\�� a?0/�?��?��(?j�����>�ܾJwM?�U6?Q:�>�&�2�t�_��=ڀ޼0ⶻBW㾉V�-��=ln�> 0>��,��{�&TO�މ��v��=���"�ƿYV"�8����=7�0=? m��/��D����;�����c��ｮ�<
��=�Ie>k}>�`\>&�1>�j]?g�n?��>��c=�s��ٕ��-ʾ�O�r�����r�j���H����ྜྷOԾ���n,
��e� ���q@��^�=��Y��Η�����`��~7��'0?/��=-���nE�w�@<0�̾C��Gz��t���Pľa0�>[k�F4�?�D?��{�J�S����V&��ĥ�&ya?��ҽ�������݂>^��5�p=��>�S�=8L�/��gR��0?4?}h��C���v6>2��>(B=]�(?��?^�<�y�>u?,v0�H����2b>�P>�>g��>�� >����cyƽ2�"?_NV?8���ѣ�p�>U#���N���׵=�=;B8�A5���H>[崺�g��� M��h�x�<�zb?e�>�d)�N�'�^Ǿ�˪=r��>�Z?�@?�Ǐ>S_�?]�G?�#=�\��j��D��R�=�nV?Ǿl?��>���2����a.?���?� N>��G�Q�*a���о�x!?/�m?�?Ď��p��F��MD���D?��v?s^�{s�����S�V�S=�>�[�>���>��9��k�>�>?�#��G������lY4�*Þ?��@���?��;<�����=�;?U\�>y�O�I>ƾ�z��ȃ����q=�"�>ጧ��ev����wQ,���8?۠�?���>Q��������={ٕ��Z�?_�?���AFg<��l�Gn��{�<;Ϋ=6�V@"�I��}�7��ƾ4�
�煮�迼=��>#Z@T�w*�>�C8�&6�TϿ#��b[оQTq�E�?:��>3�Ƚ����B�j��Ou�r�G���H�������>?�>L7X�5߈�r�z�-T>��n�I�>rs��J]�>�0b�M���I���[�w��`�>�#�>|ߑ>�y�����{�?�a��$7п1���U�q�T?��?��?И&?&	;B�C���]�keL���D?�n?(�M?�I>��JT�~jX�S�j?	_��WU`�Ɏ4��HE��U>r#3?�A�>�-��|=H!>���>oh>�#/�p�Ŀ�ٶ�$������?Ӊ�?�n�e��>ʀ�?Ss+?�h�V7���Z���*��%+��;A?*	2>�����!�/=��В���
?�|0?��=.���J?5�[��P�7�����=�X�>�nɾuV���V��Al�E.�V��͇����?lu�?��?(4?�����&?Vm�>9���CB��k
L=� &?^	�>��ļ�?v>E�=n#(���6�W֟<^��?0�?f$?#��ѩ��?�=�׊?�ߠ>t �?0+�>K�?���+���5��=�`��+�^>��<���>"�??J�>�o�=+؃�K���E��xr�ǐ��6R��A�>��T?��`?��R>�C���H�?�L��0�������l= ��v�-=�*e��8>B��<H�=0=���ž0�?�o���ؿ�i��	o'��34?̶�>��?���6�t�����;_?Xx�>�6��+���%��eE���?bG�?��?�׾QT̼c>��>�I�>��Խj���䀇���7>��B?_��D����o���>���?�@֮?�i�U��>Ǭ�%N���:|���6����]<T�E?}Õ�~ �>�D�><�
>5/��NO��)�r�}�>�9�?�$�?�>qB�?S���*rT�\�ko�>�?�O1?���4˵���=}�
?��*�ĭ���Q�1g{?��	@x@&�_?�R��]�ؿ�ԕ�ݚ����
0>۴�=>�Ǩ�]��=u�<���<����5 >&�x>K8;>��F>�W>�2�>)	>=����"�%e���?����>��	�J�ﾬ齒���]`�uB�����@���i�����گ��|JE� �����Vc�=	V?![R?�ip?�G�>\x��F >=����
=��$����=K>�1?�L?��)?�:�=���>5e��w��my��x
��ڄ�>c�H>�R�>��>+ǭ>2Y�:��I>��=>鲀>�� >p+%=E�̺8+=�N>��>C��>*��>$<>;�>�δ��5��ڙh� &w�̽��?����>�J��-��2��e���&��=�\.?){>����;п�����0H?}�����+���>^�0?�OW?j�>������T�i4>�����j�'_>k6 ���l�(�)�\&Q>�i?��,>�>�/���P��hN���־��>�*G?%���0'�3*X�>(%���C��>C��>���<��!�e\���7|���^����=-K?d�?X�j� ���Ͼ�i���>�v�>��^<���=��=�Я���-�2�f��*��	%>h��>_�?�3>n=�='Q�>e?����P�&�>� A>d.9>e�A?ό!?X!�ס�'�y���2��g|>��>�5r>�R�==-T����=���>�o>2������C���%Q�k�G>��X�2�^�E��Ux]=�������=׬�=5
���<8� mE=	�q?� �����˃Ӿ씑><{P?�˽>!�=>t²<|�,����}ɾ[��?Ws@���?x�$�2�M�<g0?���?�5�^,�=;a�>���>� ������%?olg��ޥ���h������?�p�?U�������܀�U*�>��$?M���l�>^k��V����3�u��#=!��>�:H?UN��O���=��u
?�?2m�h�����ȿ�ov����>`�?1��?z�m�fB��Y@��~�>V��?kdY?�Wi>�?۾;�Z�-��>]�@?kR?��>f9�Ǻ'���?nܶ?��?zH> X�?
Bs?���>p&x�n�.�C泿e���vuz=^�;�~�>V>������F�!����r��LGj�)����a>_�%=��>�{ὓ�����=�׈����K�h��ɶ>�	p>�FJ>p��>V� ?���>y�>Xb=�È��/���[��#.P?=�?Q���_�����8?>�����?��Q?�1�;����74�>��A?�~?��=?K�>F�����5���	��� �==�>`��>���>��k�Bi<>��	&o��o�>O$2>�̙��ѾA�U��g�!r�>s?@}�>oU�=�s%?�?�=V>��>��K�� ��X^.��T�>5 �>v�?9m�?�S?֏��9f>�������v�B�Tn>�>r?u�?�Æ>Ԥ���ן�L�˺�<*=�W㼏�s?�x?u�;�:�.?�܍?��B?�)<?*�A>$ur�z��=�i��Ɍ>Eg?ci<�:��+��Y>2��>�
�>h��>#�>�`��{����4�S�����.?��? +?مݾ2&o�����I=.u̽����,�=��<�p�i���M<"�뼹5=��R>[ݿ=/u-�,3��������3=���>��o>����[�3��,?��A�Dd����=%�r�wiD��%>�FL>�;����^?�i>���{�����9v���U����?n��?
h�?[X����h�l=?��??1A�>O<���m޾iD��w��w��s� �>g��>�|��a徦|��pv������[Ž &���>�G�>`�?L��>$@>A8�>�?վ%: �fr�Y
��(C�t���bE�q�0���(�����\3�����.���X��t�>�㰼fב>]�?0��=8�3>g��>Y.���#�>�F/>t�[>�6�>��S>B;.>ZX�=�m��It�<nQ?�Mʾ���t�Ѿ����o�<?�S?�4�>�x���ʂ�ߐ��T5+?�5�?�l�?l�>��X�ë��{�>&}�>�����"?�d�=�ۀ�D�NR���NN�x�+��J�=�(�>w"��oG���W�}�*�<�?��?u_���'��5�>�㏠��o=�J�?K�(?��)�l�Q�Y�o�w�W�)S��^��1h��`��w�$��p�x쏿H^���%��j�(���*=|�*?�?1������%k��?�
[f>J�>0$�>Tܾ>[wI>:�	� �1��^��J'�f����Z�>^{?��> �I?��;?�[P?�|L?���>�:�>�-��
a�>��;��>���>��9?+.?NM0?kl?{W+?�2c>���������wؾ�?;�?�I??i�?�� �½�ȕ��h��y��⁽���=h\�<l�׽�>t�QS=]�S>�(?7 ��9��.���u�=�M?��?5ۡ>l�$��V����->���>�h	?��1>��䅿�u&�*��>ڡ�?T�޼����p>5o>��V<JA=	3�=��=WF�= U:��b?���ϼf̱=M!�=i�=�&=Z�ڽN7�蘟��#�>��?�>ݓ�>� ��$�$��ܾ�pZ>�`E�v��>ڜ��2�J@��롿bd���>�D�?��?e>O��>��L=�+���'��&%�bǙ�ub�>���>��Y?�l?���?f�V?�:?�
 >�)����O0i���]����>_�+?_ؑ>~��h ˾�ը��3�ð?C�?�k`�����(�$����׽l�>?/��|}��ٯ�D��������E����?�͝?�K?���6��\龒���A���qC?���>47�>��>��)�6�g�*&�Nx:>E��>.R?&��>�K?e�k?7[M?���>(N<��ﳿ�I��8O^��'ü�2?�\?��?�ƈ?�� ?7�>Rd}��u��p)����,����i����!��D�>@�>=�>E�>��>:�y��ֽK�Y���=+�~>�K�> �>�v�>A,j>��e=e�G?<��>�T��8i�_	���U���VF�N'u?LQ�?��*?�Y=�����E�s�����>,��?$̫?H^)?ɚQ�ҩ�=��ռd���{o��^�>�v�>�/�>�W�=�r==�t>��>1+�>�Y�^p���8���K���?�F?^��=;/ƿq�o.u�Ů���M<P-��S�_�����^�\��,�=���7���ũ�e�Z� ������$���Û�1�}�� ?��=�)�=��=���<����<j_`=��<�=+m���<�@��ј��74%�	4<�:=�.�m9�,��?��?��n?Z�>�n<>/�o>���E(�>醛���;?��>D.�g����c���˾a�3T/��oB�p���-�c�|�=>���*��>��a>t�=�
2>j�Q=�g�W�>�'���AP��n�=��>H(�==N�=(�+>�5�=t�n?����c����Y��7��M>4?��>�	�=�i�A�@?s�{>L�z�Eu��?�&m?��?�Q�?}�?���`��>�y��ݙ���0�=��>"�>#h=�e����n>cb0>�K��I���{�=���?X:@�.?uX��.9Կ�4>y�7>�i>	�R��{1�P\��c�>�Z��e!?h);��S̾��>���=�߾�{ƾ 0=Ҵ6>~�c=� ��\�gz�=Պz�O�<=Q�m=f��>=�C>��=!d���~�=)J=�:�=��O>Fꦻ-:�S�.���2=a�=�xb>s�%>���>�?mI/?xRb?���>�p�p�Ѿ�����L�>W��=Q��>�Ij=�bE>ڟ�>;9?ڃC?#yI?~��>��=ͥ�>��>�i,�5�m�;��������<C��?�Z�?gt�>��<�E����6�=��Sý�W?M�0?l9?��>�����ۿ`H���	��ו��I>K&>���]�=?�`=���8����=lb>6��>�>�>�79>�+�>bs>;��>!�=h����Ź0�ͼOw�=�e;=s=��ļ�9>��(=�@�闑�H�����<l��=�I�@���s��%��=�X�>T8>�0�>Oc�=Pֵ�g%,>O���J�%^�=������?��>b��~���.���;�`YG>gIf>������� ?,�V>.dH>E��?�t? �>(��cԾ[���R�
_J��N�=B��=�E���<�aa�$tM�R�˾4��>��>��>#�l>�,�� ?��/x=:��U5���>Ox��1��6�?0q�j=�����i����f�D?VG�����=!~?��I?Lߏ?���>1����ؾ�0>�]���#=���q�������?$'?���>3�ؽD��KؾRI���ۈ>dw��|�2�Ɋ���=O���&>�_���K�>R@��WG��ZH��{������h5@������[�>�oQ?��?�gʾ�&n���(��?�������>��:?�~�>w��>��>н���䘺�PY==xKr?c��?��?�f>��=3���Z�>�b?��?�[�?��r?O[@��9�>a��:�1>~��j�=��>���=�7�=~�?�3
?�C?作���	��%�L�]�,9�<��=W�>J��>Tvs>�S�=��e=�&�=�Z>�͞>#��>��f> �>N&�>輥�G�
��&?�O�=kӋ>��1?�{>��-==β�=Y�<�7[�#�=�:�-�q<ƽ����<�J��F}i=ec�����>�nƿ���?�7Q>;A��y?����?��O>0S>;Iڽ���>��F>р�>�ı>���>(�>��>�,>���ѻ)>��&J7��&1�U�r�*���P�>�ϊ��Rh���B�޼(��rb��K	��w`�7�+�/�K��<,�?�~3� �D���޾�� ���>���=-$?*-��n�˷�=^ ?�F+>��� ��������99�?�T�?�z3>� �>��b?��?��n�qi&�ad��:s���L���7�=�\�q��na`�����E���R? n{?_�??V�>Ajw>L�U?'"쾐�����i>�k;�j�2��8=��9>���Nl1�����}2;��l�=��>ܾr?�g_?b� ?����z�m�� '>r�:?~�1?�Ot?��1?�;?�����$?�m3>LF?Cq?�M5?��.?V�
?�2>��=�����'=�6��*���D�ѽ�~ʽ��{�3=�_{=�+Ѹ�<�=C��<����ټ|;�$��|*�<�:=��=��=�+u>�J?]�#?y�>?��p�9j>��Ei���>��<>�R�[̾�����%����;�9c?�;�?�fc?��>�0U�����0>5R�>*��>l��=��><��&͑��">$�=-�>��<ƨO�:Ⱦ�O���s����=\��=NV�>d;�>��=��>A����1���w	=��佂v̾y���Z�.��F�����.>�>��=?��G?(`F>����e =Uh^�!�?^|?!�u?a.?���=����I�ž�h�}c�>`�\=��
�E���`���̭���(����=|$�>�S�I�����J>�I!���$v��V��挾]�F>+���tf=����
i��̬o��[N>�*>�C���L��������e�D?1<���э��ھJJ8>ᘔ>���>k��R$A���K������-B=&J�>s8->9���� ��]�D����<�>:PE?:Y_?rk�?�!���s���B�����j��;qǼ��?\t�>�g?�B>�=���� ���d��G�$�>��>����G�<���-��k�$����>�;?�>l�?��R?��
?D�`?�*? C?&$�>���o��� %?n�?�-�=l�޽wUL��`9��mH���>�'?��N��)�>X�?�?��%?U�T?�2?&s>]� ��;�;'�>�s�>�DX��r��ɼ_>��I?�ɰ>ȐX?ۃ?�f>>V4�����t������=-�#>�2?�� ?�?��>8��>����׀=Xz�>c?^!�?��o?,��=��?��1>���>˕=�H�>�_�>�'?�qO?��s?��J?M��>��<xc���j��s�
&K�]�{;�wH<MC{=B)��Xt�����
�<�r�;z����o���B��B��?�;���>b�.>q憾�"D>�8��š���J=�V��)?��B���`���J><�>ɣ?'�>�۽k�p>9� ?�[�>^C�/�m?�l�>:?�Ƚ=�?m��Z�+]^=���>1?�m����\.���a��$>y�J?�J?_!��!Tw���p?��I?e#���;�Ɍ����!��	���9U?�`?$kI��A�>T,}?��f?�Y�>�n���|�G���(R�6���f�=�i>� � �`���b>tK?��?�^>��H>����\z�6d?ԍ?Y�?TR�?{�=��`�xi�<��wG��^?φ�>�9��m�"?V� ���ϾWX��� ��Z�E�����qD��!v����$��΃���ֽ���=c�?�s?�Zq?��_?�� �� d�U.^��� iV�h%��!���E�%E��C��n�F]��*��*����G=r݀�2�=����?E�*?�
1�;�>a���L����ھ��f>n���כ�규=P{ԽH�<^ZB=�"e��7��ᦾ�!?$@�>R��>U�:?��X���<��.��%3�zt��+	:>ݠ>{q�>��>�![;Bs0������;v���گ�m6v>yc?p�K?ҹn?{p�-+1�r����!�Q�/��c����B>�k>��>n�W�ϝ�&:&�mY>���r�t���w����	�ҧ~=T�2?�'�>[��>�O�?�?�{	�Il���jx��1�;��<�0�>T i?�@�>��>�н6� ���>
�l?���>�K�>�����g!��{��V˽���>EL�>�0�>ؐo>&�,�J\��l��{���9����=F�h?����`���>R?u��:DE<�y�>�3v�¶!�:��߽'�D>��?pn�=UW;>��ž�3���{�;����*?��?(Γ��>*��w>/�"?���>�m�>��?I��>Z�����:!�?�S^?4�H?|zA?��>��<���E�Ƚ�X�l�1=^q�>5�a>�:=?�=V�"<`�����N=B�=�f��N䲽���;2������<��=a9>;mۿ�BK�g�پ�D�s?
��爾����d��Ų��a��-��OXx�����'�mV�17c�𢌾��l�Ǉ�?�=�?����0�����7����������>z�q�������)��c)��ǖ�L���Kd!���O��&i�u�e���>O���9jǿ�A���*�� ?�D8?�^s?�0���jT=�ƨ\>E;�;��E=���r|���t˿oq�qzR??��>�$ξ�Q<���>w��>��=C�K=1y����~f=}�?�~)?� �>�u����ǿ������Q��?�@�SL?խ{����Y�
�f��>֭V?��s>�����ZS�����U�>���?�?O�L>�P��0����m?#ʿ=�~S�d��=|�>�>���<fܾ��B=A�f>@��'�%�
����>o?ý&�Á��A=V�*z.>��c>�|�=SM�Մ??z\��f�^�/�WT���S>��T?2)�>d:�=��,?�6H�Z}Ͽ|�\��)a?�0�?��?��(?ۿ��ٚ>:�ܾȉM?�C6?���>�c&���t�b��=��8������%V�<��="��>�>!�,����^�O�hC����=&�ܵƿ9�$�.x�H�=��ںg�[����j��|�T�)���]o���Gh=bu�=qQ>�w�>�EW>�CZ>:gW?�k?�U�>�g>8e�I���kξ ���K�����������磾/?��߾�u	����<��U�ɾ�D����=�GT�U��`#���e��>;�w�3?�>7�ƾ�,H�NxB< �ƾ6���DU�򅗽�p̾R�0�R�s�yÚ?�F9?·���
[�����@��S���IU?e�����_���O�=1����P=0G�>]��=��q'4��U���D?hY?�α�RV���Q >��Q��^>�_G?�|?4?%>@�>t�!?�"l�*<j=��>��>��>L��>S��=\�־+@�<|J.?�1O?�ʼ/ �k��>c�־T��Q�c>}I=�:�}^�P>��;5���F�=���=�Ŋ=�\?�Ӌ>'�����|��,���=�Dy?�?u.�>�p?�OB?v��<.;�o%S�k{���<��Q?�8k?��>�8ýb�5촾��*?Y�k?�~>ad��Xվ,/9��Q
�׏?�i?u�!?��k<�v�ɏ�������)?~�u?�h^�aM����vEZ�G��>��>p,�>��8� i�>,~>?��"�(d�������@4��Ş?�e@׈�?X�M<f��S
�=�?���>iP��3þ�h��oY����r=Sg�>B���� w������(���9?Ỹ?��>�>���*��=ڕ��Z�?\�?����&Gg<���Kl�Ep����<�˫=���:"������7���ƾ�
�M����꿼(��>Z@�P��*�>�D8�16⿬SϿ���Zо�Qq���?ހ�>ٟȽ����{�j��Ou�`�G�y�H������R�>�\
>�?��V���|��:�7�F���>Hw��#,�>QmG��ڲ�㠾8��:���>�Z�>+��>{���-���Y�?����K&ͿZ���&�8)[?J�?Ǖ�?n�?�g��qG}��(~��� �y�H?զu?�wY?��6�/j�C�f��j?�_��zU`���4�pHE��U>�"3?�B�>H�-���|=�>���>�f>�#/�x�Ŀ�ٶ�M���W��?��?�o���>o��?ss+?�i�8���[����*�y�+��<A?	2> ���O�!�M0=�dҒ�ļ
?\~0?�z�L.�"�U?����Z��D�1�r�=�g
?�(���-^���`<�`��~�J��\���ߏ��ê?��?� �?�c��� �� ?��>(ؾH�ľG��=�R&?IY�>��=�Խ=o4=7���Y�3�4
n=���?��?�j?J���Ө��E�>ٙh?�p�>%4�?�o>��?�l�=���ͣ=��B>�W>�=��>�iB?���>=.�=E�R�a�D�)�Y�c�`�@m]��=�>i
c?��|?!Z�=I��ֽ�(/��J���޾3_Ǽ�zĽm��=b��9�>�>�Z�t�־��征��>��ّϿ`љ�2D���>[uI>�?6�׾	��@��=yL\?0�>�A�Fn��P}��-�c����?JN�?H�?:��p�}=��S>�p�>�Q>����Nj��.&��>Q�O?�������]��$^2>t�?m�@�ΰ?�tB�Ѝ�>v�
�}>��Y�y�Xd�����a/_=�9?����r��>�^?(o�=���E����{�b7�>¡?ZG�?rr?8nh?2s��N%����=7�>5�r?/$?�������N>���>��*��و�uվ��?�	@�@��$?�Ȥ�
¿Jty�뜮�{�Ծ`�I=�p�E̟>�Mu=��=JO9=s��=+�<��>��>�3>��g>��$>W�*>f�0<�~�g����˩��k`��7�뮾�:=d/ ��Z�[�&���*�����<�'&���0���Q��+d��C��=��U?]R?�p?*� ?&�x���>���}=�#�=�=�6�>�b2?1�L?P�*?��=3����d��_���G���������>�kI>hy�>�L�>h�>?!,9��I>�
?>���>.� >Lb'=�K��]=��N>yD�>S��>xo�>�==ܕ�=����K���FMx�8Z���B=y��?HR��e6�X#���q�M����V@>�O?���=����)ǿX���Q_?�Ե�-p�5����=]6?)�E?5�<=� ��N�i�o�S=A:��u�Y�e|�=��/�����X,���t>61?7Q|>�<s>�L3��7�p�Q�������>`8?���+�;�Bp���C��׾��R>���>'-Ѻ@��=T��ߗ~�6yf��g�=+�7?�� ??���hϸ�� ��Zw����J>�l>	�?=Z��=�A>�<S�/ս�?�f+|=���=L�j>!-?�0>�9�=��>����{@T�G~�>�I>�1>K�@?�h$?�<�g�����.�(wt>-��>�}>c�>J�P�dg�=;��>l�k>F�������u�^KD�bN>��n��`��Xv��|t=����7�=�y�=�3��v�;���'=�oo?�ۺ��A����Ӿ0DV>+�`?�J�>��>��������d����ྔ��?�
@�q�?e��_�M���6?HH�?+�ɼ��=�+�>0 �>����`�k�i�"?-I������+M����?�]�?1����蘿��˾>qy.?M��35�>~��!1��	���zw��%=���>�H?]��&RB��,���
?̷?���-����Hɿx�
��>�s�?g�?��n�6����zA��s�>���?�C\?4�f>Z�Ӿ�m�֨�>M&A?eP?�4�>R��д%�u�?��?���?��H>˄�?��s?K��>_�x��e/�t#��d���{�|=��;b�>�>����Q�F��ٓ�a��4�j�����a>�|$=5�>�[㽼���<�=u+���1���f�%��>^q>�I>�^�>�� ?R�>���>��=G��g‾���!�]?��?���Pbc�Ɓ2�� >��"��?�[V?��!�u���Dɯ>�.M?�ey?��C?�
�>7��8��_v�����x�=�V>{X�>�I?�q��� >Ų���b���(�>��>�z: O�\�C���;��>	�2?\��>n)>ml1?�P?�z�>	��>-�J����ka��G�>Y�_>� K?ܘ�?�l�>�Un�8bE�N��������M��yN>�:�?�qS?�cS>�M���m��g2�pu�=	�<���?o��?"�ӾS@F?���?�J?.�o?�C�>�8�����O���T>��+?sӭ�?9�o�!���.��?G6�>���>Z?�=ؖC�ѹ��w���|?�d?�9?����dd��쩾B
~=�|q=@Q��t�<>7�<��=IE�=@��B!�=$�>�g>��j��|���:��<J��>��P>'A�C���y?=B(=�Z���:o>�Y���>�O	x>��
>@Q��gy?�Z���_|����8
��-
�����?���?Y��?r�Ͻ�`�[/?}.�?K??���>>�þ��W�pR*�q���`>BR@��6p>��?�B��P/���������]�TPc<	c��6�>�M�>y�?~>�>p��=-v�>W�Ծ�?@�����c��}�Q��p
���S�,3� *��f�VwI����<O����ފ���>�ԫ��v�>��?aa�>�>�>��<oJ�>��q>��>�D�>�:>�>	�=r� ��ϻjFw?f뾥��꾞���c?�Ҍ?Q?��N>����J��e�5?���?���?/w>p�M�QU�䭠>�!�= -G���?����=)�=�4e�p���>�����>FH7>�\�-���+��l	�~��>eOB?珖=Ծ���������=�8�?�9?R$��MV��X��gU��f�ߐ�=�����V��1�����X���v}��6�@��y�=j|/?�%�?M5��Jkﾒ<��H_���6� ��>e�>�~�>���>O}c>�龏��@U��$��c��n��>�nx?�y�>5�I?�;?&sP?�eL?4��>�J�>N<��t_�>8�;g�>���>�9?��-?O50?.u?lx+?�Tc>g���
��zuؾ�	?k�?�J?�?�?�݅�˖ýR����~e�$�y�c������=P]�< �׽*Ku���T=�T>!Y?�����8�����.k>��7?P��>���>���4-����<��>�
?,G�>* ��}r� c�V�>k��?�����=��)>`��=N���kGӺ0Y�=������=�0��]y;��d<���=���=KYt��M��i��:P��;�o�<o��>4�?2X�>��>p���s� ��V�r�=C�U>K�U>��>,ھCo���@����g�-�y>a�?vH�?ƽg=���=�c�=(+���ܽ���wƽ�|8�<�Y?<`"?S�T?�2�?M�=?��#?F�>	p�e.��4Y�����3�?��+?���>~���#ʾK⨿(�3���?�#?�_a��5�}n)���¾�vս�%>k/�8~��诿�C��z�����֐����?���?� A���6�f+�(���杬�.�C?)��>l�>}��>d�)���g�t8�2 :>`�>�R?��>�O?/�z?�+[?�QU>��8��N��DΙ���6�L�>s�??Je�?\Ŏ?��x?5��>�>D)��#�����vt��#�@���V=k�Y>��>��>,��>��=ȋƽ����h?�;�=�|b>g��>̥>�|�>yjv>��<#�<?���>����r����|����'=9?�|?$$�>$��=[>�=a����?e�?a��?��?+3���S>:���&p��f2�3־>6݇>� a>��>:I�=� >���>u��> 5���`�5�~�ν^�?&�2?������Z�`� �J��B��Rp�=&��t{t�Μ��ޕ�O��=빡��[��ۡ�vs�d���ͤ�3ш���F���=��?$�!=�+>�8.=����X��'w=�=b *��U����|�<�����tJ=��(�& �=��
=��<�=)K��?}?�߉?�i�?�mD?<Ǧ>����K~B����>E�羴(B?�>�O9�C��d��ؾ*'޾��2��I �Cfh�z�ƾ��=�@��V>2r�>^=�ǋ���
�;��=\��=��սPoF=���=9��<eQ=�(>�'�>g�D>g�_?|[�������R�o�x��q,?j��>��=�郾�A?�<>����K���>q�H�r?1��?W �?���>�,9�.��>&F �k���=)�>u&�>o�w��N�>��>�1�Ko���$`��q�?m@32?�a��:T߿5U�=R�7>��>C�R�%k1�W�[���b�t�Z��$!?;�l̾b �>���=;�߾0�ƾ��5=�#8>Pg=�B���[����=��{�Kc;=%l=��>ߔC>L7�=<G���w�=�J=���=VsO>ɇ��F;���.�;2=���=��b>'X%>���>ɏ?ܲ?��E?'F�>��p�af澰�ھ��u>q R<m��>~~����=)<�>6�U?h_?�H?꣒>o�$>��>��>�d!��,U��lվ �����=⛁?��?C��>��T=)K�ͭ&��:�IC��?��7?#l�>��k>�U���� Y&���.�����=-3��+=	nr��SU�����wm��㽌�=np�>g��>��>�Ty>��9>�N>��>��>9�<�o�=kꌻT��<h �����=$���z�<�vż�����r&���+�w������;���;}�]<���;3�=C��>L�>���>N��=���*	.>h嗾YM�o�=���B�|�c�Զ~�?�.��G6���C>��Z>ʂ�2��t|?D�]>��A>F��?x3t?m` >b� �־�I��DMe���Q�m �=>�(?��;�X`��XM�c�о�n�>�ݎ>3У>I`n>+�+��>?��Fz=�l��5��^�>X����3 ��?�ܴq�Y<���͟���h��W��~D?�,���-�=�Y~?̶I?ζ�?���>f闽&�ؾ�/>l\��q�=`����n�)���(�?@�&?�g�>/�뾄5D���ƾ�����>����5M�r��&D)����ʾdr�>������Ͼ��+�N���\����?��/u���>dfR?`��?�z[��n��o-S��'�Svx����>��r?T߳>� �>?vg�i1��S��:�= �c?\5�?�Ǽ?�o>���=�����>��?���?��?��r?lnA���>���;y�>����=�>
>��=|��=Σ?�
?��
?�Ú�M�	����)�Ky^�\!�<��=Ƥ�>͌�>�fq>�c�=�g=��=��\>���> a�>�Ae>���>�>4쫾ƈ	�rj%? �=���>�/?�u>��<�e�S�
=
}�4:�wq)���н����8�;�G�<#��=��&��>��ÿH�?�?>���?1)�D*�݌?>�AB>ŋ޽���>�OD>�~�>�V�>��>+>ut�>��1>®ݾ���=�x��,��5L��M���(�>�ʓ�&��.��Mӽ�C�y�����2�f����uf<�����ي�?���=b���mU����?ƌ�>I�)?�m��o���Uw>۱�>���>:6 �qϔ��������?� �?��=^��>��E?�6�>���Z<���c�@���[�U���f�QqK��N���]U�J���>1�f?y0y?w�8?�8�>e=�>ۂ?�<+��̾�z�>�4��L�Sv�=���>����:�^M��)���u�)�Ϭ?e��?�.?Lis>t.!��}�|`'>�3;?��1? Yt?U2?��:?/�h�$?��1>��?�?�4?oW.?$>
?�v0>N�=�����-=C푽�݊��Yӽ=ͽ
i�� 6=X�=	��9\��;O=_ �<3����)ӼWN;Im��Y�<0W<=䮤=���=e�n>+&M?.�>a�>��:?#z��Lb��>��z��>Z�vvH�,�0���_�Q��>�v?5�?�C6?��>`�#�N�3��E>
�>Y�E=eYu>��>v���򳾀��>�`>��=�ޚ�nL�)'ݾ�����u�92�=��<&��>/с>r��G�(>ˇ��������;>�Ad�yB����Q�2M�Ο1��r� ;>s{K?��?�9�=o�Ѿ�O����f��V*?89?`J?eG|?}x~=KZپ>�1��"G�`{����>���C�;G���#��2V:���;_pp>ȸ��=��T��=�FQ�P�žIg���H�@�����R>����>e�Ծ��B��iɾ(�i>�@=W��b������Y��>[?��p<�vI����ﾐ�>"�>c��>�lT=��}>�OZ��o� $����>��>>R=fʾ��[��N-�Y��>�5E?h`?τ?z����r�ڞC��>��OI��M[����??K�>�D?:>���=GZ��D���c�WE��
�>s��>���c�G�+���=����"�f��>��?�| >�?�mS?K�
?|�`?�)?s�?�D�>I���h����B&?���?�=��Խc�T���8�ZF�V�>/�)?��B�մ�>�?��?1�&?U�Q?�?��>0� ��D@�ޑ�>�X�>��W��a���`>n�J?���>q;Y?�ԃ?z�=>D�5�4좾%䩽�P�=�>��2?�5#?��?몸>g��>C�����=c��>y
c?0�?f�o?el�=�? 82>Y��>��= ��>Ո�>�?�WO?�s?��J?���>X��<�3���1���!s��rP��5�;A�H<��y=�~��5t��\�~O�<DȲ;�?��B:�����t�D���޺�;���>P2s>�ڕ� :/>^�žޭ���B>����������K=����=?��>�?[��>(�"�2C�=�G�>}��>cQ��(?��?��?�_E;�b��~۾'"M�@��>�B?z)�=U�l�����!v�Z�_=jwm?��^?��V�����>�m?O�J?�aȾ�E���ܾ$���\N�4E�?�I1?�^�}@a><�?C,�?�:?pǤ�cl�o����O:��w�^��=�Y>�\N�+Da�_9�>�=[?�I�>5<�=mi�>e����Ɉ�/��>�fm?�Ƭ?R�?��z=�I|�X5����Y��Ǜ\?2;�>X}����E?�Tw�Uf��鮉��"����]Aʾ�����o��2��U���L���0�ӏ=�?т?X��?�oN?����t���z��_���,����Q�C-Z��I���D�c�r��t�ٴ�����᏾=����?���?R'?�>-��y�>�l�������;L�M>ә�:���t�= ��m�U=fPf=e�q��9�O<��?系>s��>�6;?h�\���<��G5�U�5��&��*>x��>���>��>�`����/�h��m4ǾD~�I�Ƚ��t>D}c?��L?��o?������0�a!��8���gQ�Gg����H>�
>��>}z_��"��M(��S>���p�(����Lm
�	`�=�_3?�h�>���>0�?N>?G��G��� #v�|Z0���X<� �>ӄh?���>(�>��׽�l �(��>St{?mC?K�u>L���j�O+���\;���>�@�=#�?��I>���Sk����������?2�s�>�|?q����HȾ�S>�8�?W�1�xhk��,�>؞*>S�Z��Y_�[�^=��z>�3�>�h�=c�>���}��+2k�)D[��O)?nK?>蒾 �*�5~>%"?ŀ�><-�>+1�?+�>~pþ�D�б?��^?+BJ?qTA?aI�>-�=���G=Ƚ��&���,=ه�>d�Z>� m=]z�=����q\�gw���D=�p�=T�μO����<!�����J<���<_�3>L�ؿ��>�����pP��Ҽ�����u��!������tǘ�Jw�/����x������2��cu�*�?��ֈ�#^��p�?{y�?}����T��g��-rk�wG��1�?R����Q���@�v�!��O�����X�ľ��0��"N���b��d���'?������ǿ����=ܾ� ?�A ?��y?��Ý"�U�8� � >�/�<w8�����њ����ο���'�^?���>F�{.��Z��>c��>z�X>Cq>���h鞾��<��?H�-?���>ǔr�g�ɿꊻ�a��<���?=�@u|A?��(������U=��>@�	?��?>�B1�	A�(�c�>D;�?���?��M="�W�Z�	��e?�<��F�%�⻄�=w^�==���ƓJ>`�>V��AjA���۽9�4>)�>�"�f����^���<��]>�ս(���؄?��a�
�c�A/���|�Z�L>7yY?�?�>V_�=s/-?3�Q�L�ο�O�o�h?*6�?mv�?� ?IpǾ�O�>��پ݃R?��5?���>�h"�ci�{�>%����==D��@	Z���>^��>(�H>o9!�������O}��p�=F:���ÿ���n���<=�Qż�ڈ����ͱ��`�oe��D!o��@ĽT�=5�=6�U>�E�>fuh>��u>%]?�"q?�Ӛ>��>}-��ݙ�����=PҊ������f��:�_����J��߾;���~����4Ӿ�?��y\=�k�71�����&�d�R)�K1?g*=�1��
%���`=)sž�Rv��f}�*�$�[�����%���[���?�h.?7x����8���$��y���S��t>_?Kw��Դ�������J>	μ�=�G�>�:�=,�������V���3?�r?���{��'k>�����nH=��)?��	?�(��:�>o0,?���w*��;�>�p>�E�>�z�>5<нl;��^ٽ��?4�l?�SȽzZ��?��>Ό�ʬž��o>�a0>�񪽟`�=��=>�Þ�־�f�Y>'���>�(W?}��>��)��aa��v��dY==��x?��?&.�>q{k?��B?�֤<h��}�S����bw= �W?'*i?_�>���{	о3���A�5?�e?��N>�bh� ��.�.�ZU��$?�n?-_?]~��#w}�w��n���n6?��x?��~�#���뻾x���w�>V��>YK�>#C�?`>?,\Z�sD��X뺿3�;�5H�?��	@9K�?�-�=�D�i��	?�b�>'u������x�����5q=uX�>�A�Vss�e�B���j��Ib?a��??*K����"��q�=�K��I�?��?�����|�<���@l�������<9��=n;"�Î'��h��7�9�ƾ��
�[ݜ��6��]��>�R@o�߽���>��8�(E��bϿܵ��:UϾ#�s��?Ù�>�˽ki����j��t���F�J�G�������>��>����c&���{���<��j�����>����y�>��M��(���t��5<���>�j�>ߨ�>h5��F���"�?Y����hο\���k��-�X?�?�Q�?� ?��;%S}��s���vFG?Ӗs?��Y?�T5���Z�M	Q�%�j?�_��xU`��4�sHE��U>�"3?�B�>T�-��|=�>���>g>�#/�y�Ŀ�ٶ�9���Z��?��?�o���>r��?ts+?�i�8���[����*�J�+��<A?�2>���I�!�D0=�QҒ�ż
?X~0?{�f.��d?�zy���i���1��.���>�@���!������+<a�x��(���P\����?2�@���?`"ֽ��&��6#?�Ɗ>�i��,����=6�>���>�w�>@�=���>�s�6�Z���>��?���?R�?<?���[���d�=X�y?���>!��?M��=�X�>�=)��������!>\6�=`;&��?,jN?���>݉�=��:�^j-���B��bQ����D�\%�>%da?�LN?�8c>a����.1��#���нc>/��-�`j6�i�N�e5>��;>'->�G���ʾ3$?D93��ӿS]��p�ݽG�3?��>�� ?^���̴�f6>��M?�1�>�&���k�����i��*�?�|�?\�?�� �<�9>�?���>��u��A��~�?�o>4�;?r��F\�@�[�CR�>z^�?��@.��?�T�9N?��n_���k��Iܾڷ{>)K6?W�����>�
?���=y@e��6���Q{�}W�>�'�?���?�?g#f?@t�M�/��Z�=��>�e?��
?O�@<R���X>�d�>??�����D� �i?�@ה@F�]?�!���kֿ�����L������j�=���=�~2>%ڽn@�=I�7=��8��s��]��=?�>��d>N q>�8O>\p;>q�)>�����!�.n������� D�u�����Z�}���Hv��x��5��6���x6��2ý)�����P��4&��`����=�GU?RjQ?��q?p<�>�TY�L�$>]�� O=��#��q�=j�>��2?��K?��)?9��=�1���c��N���Ϩ�����q��>�F>0=�>n��>H�>��!;ݗL>k�:>��~>�+�=�Y4=Q;9�=0�K>Bϧ>���>���>HA<>w�>.д��.��נh��w�
̽ �?����ѴJ��/���/��'���r��=T^.?s>���a>пi���w2H?]���@$�q�+���>P�0?�cW?X�>d���fT� >ֺ��j��h>^ ��|l�n�)��Q>9e?��g>�V>:�F��o ��-t�DLȾᥝ>ou=?���M���mL|�Z�%�e����T�>�S�>]�t�@���� y���w�G>��E?��?��ּ߽ܾ�2!�������M>�t>���&�=V�y>�Ɲ��y�2R���D;��=v�>K3?Ę0>�m�=C(�>�4��$�Z��i�>��?>�,>�3@?_0&?�¼&�s�̂���0��Dw>k)�>�{>:�>��U����=�z�>�yq>�X��qW���KO�/�Q>�)s��c�gF�c��=����=r��=+����	@�v�m=�
?�.���|��N���=.�J�]?�0?�~<�6�=y�#�ĳ�Iվ<b�?v@�۬?dϾ��a��1�>��?�K%��_�>Q�?��t>��%���l�?ƀz��57�-7�ʵ;��ܲ?�S�?ɀ&<�]����o���=�~$?ȶ�3��>�^�ч��U+l�Z;��9uh�c�>�>?%d�Z�=Y����	?�>����笿�MǿN�g����>���?I��?�Ǒ��3����F��~$?� �? �B?�U>+㺾�$�V$�>�/?�W?���>"�)���׫?�K�?���?�y=>S��?�?���>�먻�@,�$B���j��ZT'��=��>Ȩ�=V�¾ZIR�g��ʏ��@ib�D"��	}>t��=���>��=��ð=���l���RC�;��>��>]�T>Cw�>���>q@�>�W�>OZ�<lk!�����&%���aY?�y?�n��.���2G>k><\�E�J!L?�o�?�叾�(ɾA�?>�a?�^?l�Q?�?�g5�w\���ȿ�fؾ��e=�a>���>���>0v����;�A\��AA�>��?�!s�2���ң�d�(���>�(E?n��>��[��t?1N!?���>���>F��������?���?�n[>��>�`�?�k)?¤=����n(��+ײ�|�O��f3>�Vx?,M?DT>Ip��$���h�y��`��>j�?�J�?�������>֘?O�q?�
x?��>�A��i����Iq�opH>�!?� �P�A��C&��l��q?#P?���>b��Jս��׼�������?�\?�4&?&���9a�Bþ���<�� �x>H��e<�G�M�>��>�D��Gܴ=�>>�#�=Am�)6�7li<Bʼ= h�>���=�K7�����0=,?��G�}ۃ���=��r�?xD���>�IL>����^?kl=��{�����x��	U� �? ��?Zk�?b��@�h��$=?�?S	?m"�>�J���}޾6�྿Pw�~x��w�\�>���>*�l���K���ڙ���F��Z�ŽH�5����>�^�>Kq?�-?��>[��>����9�F�t��]D޾�}b�h�3�d�.����z��pоAԣ�(�ܽ52׾i}����>�rN���y>�_?Y�T>Q�y>�>�i=I��>n��>ڌ�>C�>&�C>Z�L>��=0�׼P2׽��R?Z��F '�n��深���A?z;e?m#�>Ib9��Å�ޘ���?�ݒ?䡜?3�~>�Tf���,��W?J�>Y{����
?cC.=k�L��<������r��E=�#�>�9ڽ+h9�Z�M��h��?�m?	�R���;�H��`���r=4Y�?�*)?��)���Q���o�A�W��S�A���g�-�����$��p�KƏ��\��Q��ht(�{,=�h*?�?*�1��	���$dk�!?��5g>g��>�W�>ZY�>}H>A�	���1��^�F'�oƂ����>P{?��>�K?�",?�h?A�B?V�>W�><���S!�>��;=ӈ�>��+?	�c?J�?>�>	?��,?7�=���<P��u��U?U-?9��>�-.?@]�>�CվVg<�&޽K���G�|D��=��=i���.�ʊ5=Vy�>�X?�����8�����`k>z�7?��>Y��>���-���<f�>�
?G�>> �~r�c��V�>���?}���=��)>���=F�����Һ�Y�=H���*�=d5��z;�+d<���=s��=QIt�f;��W0�:g��;�n�<���>%f5?:��>�d>�������m0�=d��>Y3 >���=����#`~�{#���@r��RH>���?�d�?�d�=U��=�E�=�
k��Vξ���r���$��,0?�^?�V5?lK�?��V?��#?TI�=>2�츎�xm��
���J&?5\?�֎>���ٜ��̵���K���?ٌ?�U�*��<�94�}̆�����O>ޠ��󀿩��1�Y��o�|y��X����?mΓ?�Z��EC� � �>ɕ��S����&?g��>�>���>��H�
�i��n&�N,>��?��{?v!�>}�O?�={?��[?(qT>c�8�G0���љ��4���!>"@?}��?a�?8y?p�>y�>6�)���L�������߂�)W=|Z>i��>�*�>��>���=t�ǽX����>�gV�=�b>o��>�> �>~~w>�,�<�G?��>>W��0��@褾Ƀ��<=���u?Λ�?��+?�T=ԁ���E�fI���D�>�n�?S��?q4*?��S�m��=`�ּ`߶���q�%�>fӹ>@4�>p��=�VF=.n>��>{��>�$�a��q8��pM���?eF?n��=��ÿ�6n�ep��4U���SO������\�%Si�@lg�!�=`Տ��,
����� FM��^���%�����$���OC����?�|]=0X�=��=xA������x^<�MT=b�<���=~��ݴ<wX�D���b#��ؕ�;�ӧ<w)0=Oܼ0*���7q?��:?Q�@?0E?��>��Q>�x �.�Y>�L���,?�<(>���Rm��=7�����ȟ����Ծ�艾w'����>�<K�!B�=K#0>�9�=e�9=�0�=3eK=�s�=z��<�U=��>��=�.�=u�=/Q>e>0|?���� X��1�E�.� �WmF?�>�>��>fl���W?3&>ۀ�?�Ŀ����?4h�?���?�?Aꎾ��J>��l�v����?�}|b��*>>=>��B���>��`=�!+�pc��RW���{�?�@h�*?�˔�2�ֿ�� >��7>s>��R�܄1���\�8�b��oZ�A�!?�I;�7̾�3�>w2�=B7߾�~ƾ�Y.=8x6>iub=���T`\��,�=��z�(<=�"l=���>n�C>���={'��^�=�{J=[f�=6�O>�����k7�7�+���3=���=�~b>��%>"��>P�?�b0?�Wd?5�>�n� Ͼ+@��J�>�=2C�>�υ=�nB>ዸ>��7?�D?i�K?a��>/��=��>��>��,��m�5k�!Χ�ꁬ<��?oΆ?�Ѹ>$�Q<��A�#��!h>�a2Žxv?yS1?pl?V�>B/�Wտ@K?>��霼�T��[�⽏�پ�t�67��s�U�>�g���<%��>	T�>2��>�y�>�2�>M��>�[�>g�=o�Ƽ�c��#�������>,�ɶ>������N<Q�����SA�<��n����.�y�����9-��'=�4�=��>ds>���>��(>���6�B>ƣ���N�"��=tH����K���f��py��$�:�+�#�>�m(>�Vr����H��>�S>α�>�
�?I�r?I�>���;�쾧���>����W���0=�m@=	���x!7��]���P������>�ߎ>t�>Z�l>(,�.#?���w=b�lb5�S�>|�����)��9q��?������+i�Z�Һ��D?�F�����="~?R�I?C�?Ӎ�>����ؾ�70>eH��g�=��*q�Hk��_�?~'?���>��!�D�&2̾�6��^��>8�H�8(P�T����^0�a���K��\�>L���о�*3��;��e4�B�NBr�y��>�wO?���?!Md�
^���*O�*��s����?3?g?���>�D?eW?N����?��R��T�=�wn?�s�?�1�?b�>��=H����H�>)�
?�!�?]-�?�Ps?ۻW��w�>�
�<��%>�����Y�=�>��='��=;�?.�?�?}u��;�ơ����tq��I=VD�=��>�[�>�ށ>���=��=ƹ�="h>���>ᔔ>��b>�9�>��>)���v �΄?�P>�R�>�R?�i�>���nR�Q�	>��<�Y]���f`b��k���=t���c摽ln�W��>㷿$��?��>tc��?����_��Ԏ>ftd>�<��)]�>�~>���>�i�>�A�>��=�l�>}�%>&Ǿ�?>�L����<�d�%�o�
ȵ���>@z��Q$�����t��^���хľğ	��z�Yt�n�=�ϻ==��?I���[�]^$��H4���?�*&>��?�ݝ�-����>��>]�">"�}��������nϾ�ؘ?�4�?A&%>H�>R,u?�?�W��YͽNQy�+n�����d��S��x��x�y	�yZ���@?�I[?�oH?\����T>�x�?�B�3׾#�>@�S�R.J����=���>rB��/Ͼ�D�dX����ž>�=�G]?�8�?�RN?X����q��U�>�,4?��~?q�S?R�+?^|B?�R���EA?���=Ģ?P�?W�@?�O%?��>��>��9=�n���O=&lb�횾nt@�5fl�P�?���p=��=6}7�	g!<UD{=4�r=�.��=н�0�=M�L<��:�O2�'�9=y �<\��>��u?�l?�P�=d/?R�G�"=d�]=۾�(;?�O�iw��g���͹�=�3����ٓL?��?��?DP>�w*�.W���=RR�=z�>��>X�}>�\���w;�z>_�[>���>m�>d�ؽA��V�ı��@E=�|�>��>�H>6����hc�����������>�2վ�����!�0ꉿo4��o.�]�?�g?�Q?����ѾQi�=�v����F?��?�J?{}�?� �&\��C��p�=�;P�>��0�ڃ?��6��.׬��<#�Ԕ�=��.>R���c���]�~>�+1��B��s�}����Mɾ�Y>������> �V)��򣕾�S(>NZ1>�+�����W�H/��.v^?��X<?���5Q�Y)��%�0>�Y�=l8>l5�	d<i�?��_�+��>B��=ؽ&�����%I�n
��"�>�x>?u?I��?�C��y�p���N��<��(q߾ZUY=,'?��>r�?E�->"���R�վK���j�_�-���>���><��8�M�lK��Ϩ���?���>�?U1>>Vu�>؇<?,u�>�s?�*?fL?�Ƃ>Vl�~�ɾ\�+?C=?��x=�7���s���5���5�ot?��5?�׆��`&>e�?@@%??�3?��V?@�?�="��XN��g�>C��>�m��E��-��>zML?F��>j�M?{��?�{>%z=�%����ӽ��=�9O>w�=?� ?�y?p+�>���>�"��N�|=��>��b?�M�?~p?��=�x?>�4>F�>}�=}�>(�>�f?�|O?as?��I?���>h��< ���ٰ��,x�{f��\�;���;��x=/����{���n�<�'�;导�񉼔��[sB�����<t��>�Ӕ>fi{�g=>'᷾G=���}�>A�:���������\+)��vP>���>	?)��>t<0���>@�>t&�>�G4�
t0?7�?�G,?J0P��iG��̾�H���K�>��L?�s4=�fe��ȑ��+l�Y�=�Rq?}2\?ɞ��kV�>c?]?mA�,�=� �ƾZrg�7>��}R?=?;UQ�'v�>��|?A�r?WF?��[��nl�����P�b���x����=�ݛ>w��?rg���>�8?�g�>�d>��=����z������?�Ë?8�?�}�?��)>B�k�X߿A���샿�YP?�G�>����:?�`��	��k毾M�X��~��Do;�P�L쬾������KN��66!�1�_<"�
?�'a?ֵ�?@�F?�u��[�}�����q�;9M�r���G���5�zeB��B�]����%�>���]�/��=>�|�eW?�S��?TM'?QU*��%�>yp��@r���qо��F>Q������v=G����W=��v=�Ik��4�L���z�?��>���>��9?@f]�{=�P�7���6����X�">7D�>���>���>t ��xyA����d�ɾb���PȽ$l>qX?-�z?r�?:���05��W���*���_D�ټ����>��6>Ck�>�l�����J�D��7��d��)��ǆ����<�=�"?�:>�c�>pG�?,)�>�$A��y3���Óf��8 ����>;4=?T)�>kY�>;ƾa ���>ՙ?��4?J��<n�Խ�=���� �<T�'?q��>DJ?���>ojh>t����`���]����q�m�(>�;h??K.�6_Ǿ��>��r?N=��Ƚ;���]�>M�"�+54����h��>��>��h>mN>�����R4v��f��j1)?�D?���a�*��,�>�)"?�7�>Tʣ>~��?
��>C�¾���8�&?�J^?3J?�JA?���>zC=>��f0ʽؾ&���1=Jj�>A�Y>�n=�}�=�j�5�]�DO!���N=m��=��ʼ�⸽Q��;���"Q<	
=[R6>;�̿e$-��a����1j(�yXA���ٽ�>���drS�۸���X�2<����&^:Y}2�\�V�#�X�w�5�r�?a��?I���XX<w�� ���2�����?,����=dMf�z/�ܨ�o�Ѿ(7I�k���A%�3�>�g	a�7�'?�����ǿ����	;ܾ
! ?zA ?:�y?O�	�"���8��� >bG�<�(�����˚���οB���
�^?���>;�1��1��>��>O�X>$Hq>����螾�/�<��?��-?���>Ǝr��ɿ:���ͤ<���?3�@}A?��(����a�U=`��>ێ	?r�?>UJ1��F����U�>Q<�?���?0�M=�W�Q�	�~e?�<I�F��B߻��=�E�=�r=T��a�J>�Y�>���YA�?ܽ~�4>�څ>�n"�Ū���^��R�<�]>�ս$��G��?"l��VK�ԝ1�Ve��'ϲ>k�V?B�>kv>(?HY���Կ&�v���1?p@���?W6?�þMd�>G��eMl?t/?��c>(�T��~�|>�>/LW���>�U׾V�~��}�=�'�>���<�T�H)����2I&=�Ri>*��dſ1�#�9�"��kC<�G��d��c����;<���k���h����sf�=�o�=�dM>2f�>v�Q>3�]>�W?}k?��>�E>�G�h���Qƾ��<xy� J��W�����j.��]&��ܾ����t��*�W�ɾ�z=�..�=w?U��̍��%�� j���>���2?� )>~ȾN�I�P�P<�/Ǿ����A�@=���dƾ�l-���j����?��D?�����5L�_Q�eu�M�ͽ�2V?N������f��:��=���@��<%�>X��=o^۾Ϥ1���U�ގ6?&?%����P�G&�><�9ܸ=��-?u�?�ž� �>3�B?�gg={ژ=(/>G|�=�Ď>K?��;�D��Q
��F?��_?�it��Ȩ��?��龉W��b6ý=�>)ռE�0>{��>8X��jѾ��2=L��k<�>�'W?
��>��)�,��_�����L==�x?��?�/�>6|k?k�B?7�<�g��R�S�u ��Mw=��W?�)i?'�>.����о����?�5?k�e?P�N>�`h���龁�.�?T�%?��n?^?�~��ov}�$�����o6?䙀?dt��dj��갢���K<W��>!��>���>��B� ?L�8?Dl�����绿 ==�?�?�[
@<��?4���=b9L�1T?���>~�a�XǸ���=�#���&E>��>�ξ~Og��0����Ќe?y�?i?�,��(����=�֒� ��?
=�?����"�<[��mm�y���Y�<���=$�E�U��X�� �7� Tž�j�{���������>'O@�d��c��>��J��kῥ�Ͽ���`�ʾ�w}��d?Y��>�]������Ln���u�.XC��-A�������>��?>��=�Ns�ڛ��N�7!���"? �ýSEp>�,������o��fI>��[>��}>A<>������?�ѾZ��-���a`����A?ç?�Z�?��l?FX���-���ٽC�>�)d?l|�?��n?���0q��\V��$�j?�_��vU`��4�lHE��U>�"3?�B�>T�-��|=�>���>,g>�#/�v�Ŀ�ٶ�,���X��?��?�o���>q��?ws+?�i�8���[����*�x�+��<A?�2>���H�!�D0=�PҒ�ȼ
?]~0?*{�f.�h�_?B�a�:�p���-�w�ƽ�ۡ>��0��e\��M�����tXe����Ay����?P^�?s�?״�� #�46%?��>����8Ǿ?�<��>�(�>c*N>hH_���u>����:�jh	>���?�~�?ij?䕏�����U>�}?�G�>J��?��=,��>B��=O���>g�=�V>��=����>�5X?$h ?�y>n 6��,��i1��BG�IN��pO�U��>�Nb?`V?-G1>�������45�� Ľj!ɽ�v��i?��v�����->o)R>IE>�M����þ�&'?>q6���ۿl4�� 3��R�C?�Z >�H	?�Z(����ǁ�=UOB?Wd�>�Y��4(���ד����?�c�?az?�Y�� �=���=���>�`Z>�ˡ��F	�)�2���>
\V?��@���Ds���}>��?Ǻ@pY�?f�x���?�d�b#����s��C�i4	��B�=�t7?EB�$��>��?�@�=�m�����vz����>��?b��?і�>Aj?��t�t-����=f=�>"�Z?;?�v�h��%�i>�?	U��f������_?G�@�@0yZ?ꦿ�hֿ����\N��v�����=���=��2>Aڽ\�=��7=s�8��I��U��=��>�d>�q>�'O>�_;>t�)>����!��q�������C���"���Z�9���Vv� z�l2�����I@���0ý�v���Q�Q1&�GF`�?B�=�T?��N?a�p?8?]J�c�.>^ �r�
=����o=��>��-?}H?�+?�=�띾��d�7r���ר�<Ն�K��>2�D>�v�>���>y$�>�%�;5PG>�X@>
��>ql�=L�1=�i8;�=��T>��>�,�>ٺ>L<>��>Ĵ����ԥh��}x�g̽��?�;���J��1��y��|���Sߠ=ob.?">����1п����<H?�0���6���+��J>1�0?pW?�>�����V�<:>���;�j�/>Ѐ �E�l�*�)���P>_?� f>��t>�3�p�7���O�+����s~>�Q5?m궾w^6�:Su��H��޾�LK>͝�>�_ ��1��ؖ��	��*i��`x=ú:?��?+�����ņy����O>!Z>*�!=s�=WQL>0�`�3�ȽդG�`2/=���=Qx_>�?��+>C��=�>[>��S�I�8�>��=>�*>�f@?Tg$?ϸ�2��:Z����(�f5z>C�>9�~>>c>&)J��=�=�	�>��^>\v��~�#���k?�('S>�����Z��큽.�r=✕�J5�=��=�,��P�:�z+/=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ��>Ygf�� ���\���i�:��=�ތ>X�P?�D-�����cq��� ?X ?+��k���5ͿZ.���?@��?�6�?h���OW��w�M���'?c>�?\0:?�f%>���wL>�1'�>1?(e?��>�I'�=h��h?^=�?x�?r�/>���?�;w?��n>�"���c��W��gJ|���>�_�>�C�>��2�:�J�ԫW�f��?�����a�ج��<�>�>=<��>��齨�
>��N�����<�3�>w��>`x>�&�>#�
?�b�>m��>r���xC�������&��V?tǄ?1������)>�]<k�z�5?@wZ?�~\�Z)�Zo�>;M?F�}?T.P?��>2b�C��t�ƿ�T¾�/�=���==Y�>�?��2=[�<����|��Ä>��?hJ�=���˾&& �+ܞ>#r?j?:��=��?�l%?�6>�t�>�D�2��4	G���>Z �>�?-�?��?�S��7=4��\�������Y�2�W>�zw?��?�+�>�c�����G����y�?�w��G�?Wi?ҳ��ʧ?(I�?X�@?��C?�d>�A��t߾^}��7|>�=?��
�B�@�"��   �*�?k5?P�>p��������<�=
������R?	^?L9'?
����`�;|ʾF�<�s���8'u>��?����$>x >�gv��=��>��=a�s���/�`D�<|8�=�6�>I��=a�+�v�n�3=,?boH��ۃ�И=��r��tD���>�:L>+���[�^?Q�=���{�����u����T���?6��?�g�?����h�l(=?��?�?�0�>�M��σ޾��qtw��mx��w���>&��>F�m�9�ݐ��:����C��+ƽ�7 ����>�>S?&?���>�0?\���E��]���,���Y�A���L�n|��nھG�� ȡ��b�����e�9���r> {�a�x>���>]�>��>x��>�c�=��>Q��>NS>���>��>��V>��>|E�.�νODR?Z���ا'����΀��B?!d?�(�>2oi������B�?���?�q�?�	v>-sh��
+��d?+.�>�i��f
?h�;=����<�?��m!��/��{���Ԏ>��׽v :���L�`[f�T
??������̾^�ֽ?$����=^��?s
*?��3�O�'�dOt�X�_��T�g�K�V��^`��A<��o{�S��� �u�fz{�J���<��?X��?�鬾��վ1ľGjv��QN�Z
o>��>X�<>��>Ӊ=>�{վR�F�Pi�K$&�% ��N?jx?��\>��a?��3?�]y?��P?�b~>I*?]�w#?���}>3�?֬5?�0:?v�?�r?	�(?t��=�Z�<�����@�?�G	?�,?�A
?�ѻ>����pۚ;,N�=(K���b[��/ݽKH�=#z�=�L��P�O�5y�=��>�X?m����8������k>k�7?��>d��>���-����<|�>�
?�F�>; �~r��b��V�>���?����=��)>���=ߎ��i�ҺZ�=������=�6��\y;��d<���=E��=Qt��%��8�:��;�o�<�>��0?��>�cZ>������ݾ(Y ��`P���>��p>ϧ�>��	���n��T��w�m���=�v?r2�?>�>��y=k�=>�(�����8Nھ�"ƾ�5�=�D�>YW)?���?�#�?�?\?�h~>|P�Z��_�A]<�Q,?^!,?��>d��j�ʾ�񨿉�3��?.[?v<a�Q��Q;)�J�¾��Խ"�>�[/�%/~����D�������~��-��?ؿ�?�A�2�6��x�޿��\��?�C?�!�>�X�>1�>:�)�v�g�j%�2;><��>HR?��>��O?!�{?��[?hsS>��8�_?���7����r���">�J@?T�?�?^hx?X��>��>��)��$��=����]���������Q=]�X>�Б>���>S�>���=����kή���@�s�=�?d>O�>I{�>���>��u>���<s�G?���>�]�����褾�Ã�M=�q�u?���?g�+?�X=׀�&�E��E��}J�>o�?���?�3*?��S����=��ּ8඾V�q��$�>�ڹ>�0�>]��=�jF=�]>}�>��>(��`�\q8�[M���?�F?l��=tdƿ�tp��Vw�%���Z�k��[���``��Ɠ��pW��I_=暾0U	��/����A�{����[��lE������Zk�?*��=몳=��=��<����=��=���<�%=$��ܨ;1a*��T����� ���t�;��P=���v�ʾ�x|?A�G?m�+?��C?D�~>0� >W:H��>ϧj� �?7T>��d�/�����4��٥�{��i�پ^%پ��d��ԟ�v>�iR�"!>��4>���=-��<��=��s=���=����wU=/&�=��=��=�)�=�>p>'�?Å��1Y���:��э=��O?�:�>W&>SW���Y?�b.>͇������Z�2ʂ?�c�?��?�x�>�?�'j>����=�O���Y��U�>]d�9�𽃟�>p/�����7��_%����?���?�W'?�}���@Ͽ�/
>!�7>��>�R��~1�K[�k�a���Y��i!?!�:��̾s�>�l�=�!߾�uƾ�%1=�7>
�a=V7��t\���=@L{��==�Kl=Ǒ�>D>�ѹ=<���~�= �F=��=��O>䍻�S7�b�,�v�2=tT�=?�c>W�&>���>��?qb0?�Wd??1�>�n��Ͼ�B���E�>��=�E�>aυ=�eB>=��>~�7?��D?��K?Ӈ�>ξ�=��>��>�,�P�m�^h��Χ�?n�<ߖ�?�͆?�и>�Q<��A���zg>�G0Ž�t?5S1?�m?e�>%������T�i'<�ݚ��U�=v�������w�����q��n���kӅ= ��>Ͽ�>"}�>�?5>�[6=?��>a^�>�7>kJr��V��-�ɽ:�l�P^�=��j>-,�<����C��[�=�ǽ)����������(2��@=��'����=��>y��=9��>�>薆���E>e,˾��Q�7�>ިྙO���m�^����#�����j
>��'>xB������?�B>ll>�?b }?��0>p�R�(�C���dY�Q9���=]�4=
a�P\>���k��M��Gؾ���>��>��>��l>�
,��"?��w=⾾a5�	�>�u�������6q��>��5����i��g׺�D?nF��4��=� ~?d�I?�ߏ?��>9���ؾ*30>�@����={�z/q��g����?d'?d��>�쾜�D��;̾�׾�	 �>YI���O�ʽ����0�����䷾:��>�֪�D�о�3��f��������B�G@r��Ӻ>n�O?��?ab��T���UO����逆�Ds?"yg?�!�>�G?�7?�K��dg�g\��K��=��n?���?�9�?��
>Q��=ԝ��k�>�/?%�?]x�?��z?Yg����>:wi=8�>I���#�i=֪�=J��=�>�� ?ί�>���>�����M	��@�B.�J�g�L=S=?��<��>�n>Ϗc>�>�R�<9x�=�l>��>J��>�T{>p}�>�q�>Ԏ�������?j>Sj�>ң;?>�>���;e�ʽB]�=H�_�T�gU� 1�A�S���=��,�o,�<�����>�S��F�?rT.>
�-�?���4�=��&>�p>ٌo�E�>5�(>j^|>sē>M��>͖>;6�>I�=>a����>f�#�]���R�|\j�� ־���>�缾�齘j����Fmh�u/�����dp�@|��>�<��眽�?���_^��j$��k���PF?d+�>��"?C�ʾ�r+����=�?�߼>Ps��󘟿o��h�$�?��?�ZX>>S�>�^]?�?�z]�;P�7\a��v��^<��`��RO��B��!:��qM����JR?s�l?-DC?�e�<�D]>gJ�?t�������)�>ʶ4��}5�<�=f8�>�E����S�ݢؾ>P���Q�ʢ3>�|a?�b�?%�$?��'�?Ŷ>m~.?ڢ>?�9�?�'?�/W?X̜��u0?Q��{�>ԽV?��#?��T?��>��>��b="�<���><n�� - �!*�Όн�B/�>�};\���>H=��I�����<k���'��WIW=T��	>I�<!�0=@�=p��>��]?BS�>�u�>U�7?��x8�|ͮ�t/?}�8=-v��� ��Ѣ��R�l�>��j?�?�gZ?$d>�B�ׁB�+><�>��&>b�[>@Z�> Cｈ�E�#C�=�>k�>�k�=,M��ā�A�	��k��30�<�>���>�>`p�*f>*ܾB�G�1s�>iٟ�����⽟M}�زG�3�־�V�>y!T?�.?7��=9/оD��ㇿ�U<?+?f�X?��?l6�=���Cv�2^x��ˍ����>�J=G���f��<��,�X��P%��0>�c޾B��2{'>'�S������|��;�-��j��Vڭ=+�d5�=~���O#��̾v@�>���<�qľ>�ξ�o���@���^M?�|�=yą�;�ǽպ��ߑ�=��>���>�_�<��>F�F��S��� �<��>��>�;z��4��ͯN�3f�؝�>ԏE?k@`?[��?'7����r�NC�:��٣�R-żY ?���>Br?4<>F��=����~8�%tc��E�>��>�,�>���v�G�y}������$�m�>��?'>��?ExR?��	?��`?a\)?d�?f?�>b"��	����A&?9��?�=}�Խz�T�� 9�F�O��>��)?��B�乗>l�?�? �&?��Q?ߵ?@�>� ��C@����>�Y�>��W��b����_>��J?隳>N=Y?�ԃ?O�=>O�5�ꢾ�֩�UV�=�>��2?�5#?H�?���>\��>�����=ў�>�c?�0�?�o?��=/�?�:2>I��>%��=���>b��>�?OXO?$�s?��J?Ǒ�>���<�7��78���Ds���O�qт;�sH<��y=���3t��I�>��<b�;1g��-I��y��f�D�v������;�`�>��s>�����0>��ľ�S��	�@>����UK���Պ��:��=���>��?ҭ�>tO#�Ľ�=;��>�B�>����6(?��?�?+!;��b�W�ھH�K���>�B?���=.�l�:�����u�-�g=��m?k�^?��W�� ��q�h? B?�C��W5R�G�Ⱦ��(��c����?lL?�$�Njs>��?Ӗ?w�?
�f�̀�;U����3�A��� �">��>V�#���W�L��>��n?�C'?�	>���>�9��炿����9??o�?�M�?�Q�?���=!�c���տx�������`?u��>�R��:gH?��r�I���z릾��w�"誾�����þW痾W���T�ֽH��Ry�@
U=b>?xPn?X?�?p�S?zh�	3R��n��-_���B�{����j�K��cE��%W� *e����A̾6�
f>���y@����?-�'?�(-��J�>��� ��}ξ�0C>����e�����=u�����:=�pf=�l��2�����k�?0^�>�i�>Gk<?7\�/0<�s03�~�6������'.>��>�܏>�5�>�a)1�݋�)�Ǿ�~�x�ƽ	�k>7:f?n�M?b*w?����+�3�C���F_�84b�k����\_>��>��s>xT}�!t;��%�g�<��lk��J�-a���)��A�=bT2?�s>���>�I�?\?������P�X�&�/��.�Id�>Ae?�0�>���>*�ͽ ��*�>�}?�?�>?�M�%�'��E��t�̽�5�>�g>��>d�)>��%�'u��NQ����p�J��\|>�X?;���q�g���>b5i?�����+<@��>k�>)1����/��=���>��>p�>�:>�U��n��p:���k��O)?�K?B蒾��*�7~>x$"?���>..�>f1�?[*�>�pþp�C���?��^?hBJ?TA?�H�>�=���>Ƚ��&�J�,=�>��Z>�m=�|�=��Ps\��u���D=�q�=�μgP��z�<*~���K<��<��3>��ҿ�G8�
^�IO�:�ǾY���J������w�����!K�
y_�������E0�G���b��ݑ�6瀾0�?��?����'������׃����9�>ay~��� �s���/�˥��7���\Ǿ/&%��/��7U���c�G�'?3�����ǿ����Cܾ� ?? ? �y?�� �"�c�8��� >9��< {�����^�����ο������^?G��>y�4��.��>���>�X>_?q>C��Ꞿ���<��?��-?
��>��r��ɿ���h<�<I��?�@q|A?�(����oV= ��>��	?��?>�Q1�_I�;���>V�>-<�?���?~�M=��W�8�	��e?�=<Y�F���ݻ��=�=�=aX=����J>U�>���RA�i9ܽ��4>�م>�}"�?��S^��~�<��]>��ս�B��w��?�Zh�B�U��7�{$���K�>��p?���>5|�=G%? �|���ǿ�H3��w?�@ݵ�?T�?�vӾ:�>���}^?�V)?��>��6�ȫo���:>�u���=�" ���^�� �>���>jB�>���R9��B��`B'<�H>'� �_	�� ��"�S��;x�q=�Z�Z��P���8뽽R���U��"�;�=x��=�W> w>��A>��s>��^?-fz?���>)�,>��k������о��H=��x� *�f�*����"Ͼ�;ƾ�%˾&Y�=��4/������=�O��=�:Y�����W��2b�t�A���)?�&
>$վ��=��_�<2�ξ�B���R鼝~���ƾX7/��@k���?�9=?�K��FJ�]��f@��*����T?���`��F���N�>@�PRf=��>�up="�Ӿ��/��O�Ë3?8h"?ʔ��	���.�>�z��[o�=�D0?��?ӷ�=�Z�>�`#?^���k?���z>��[>e�>���>(�<awپ��꽡�?�p?�LD�Z溾��k>	d����2z8>��#>:!��5��=���">��N�=oR)���=)W?+��>��)��	��d���@�V�==��x?ϒ?(�>vwk?K�B?�ߥ<�Z���S��&��v=<�W?t+i?��>%����о�����5?��e?WO>LUh�Q��X�.�2]��$?��n?�d?��gm}�:����5i6?�Ez?HB~��ϗ�*uȾ���J$�>���>N��>��<���?ӦF?!"C����S����8���?�P@��?]���6���m6=R?���>�uW��+��Ny���;�����=A�>��Ⱦ��v���:��PH�J^[?��?Fg?IK�����5��=kԕ�`Z�?.�?���)�i<���dl�Xr���i�<�٫=�R��"�,����7��ƾۼ
����(ῼ䦆>_Y@"�&�>Q8�5�XSϿ����UоD^q���?m�>o�Ƚ������j��Hu��G�d�H������@�>�>/s��] ��"�{��r;�"\��>,�><~��ӈ>�\S��޵�����,�;<>
d�>=��>�9��Nֽ��Ǚ?�f���7ο������X?	k�?�f�?�l?a�:<>'w�5.{�Ui�m-G?�vs?�Z?�/%�kT]��f8�R�j?^f���U`��4�EE�0U>� 3?�C�>�-�[�|=2(>K��>gi> #/�8�Ŀ�ض��������?܈�?Nl�J��>j��?[s+?�g�67��1Y����*�ʗ+��=A?F2>*�����!�1=�[ϒ���
?�0?�v��0���`?Mf���l�ĝ-��O��ֵ>Ŀ�!�L���z�Խ�hj��f��-�y�׾�?�� @�ų?�	�M(#��' ?A��>�����ľ�C:;�:�>���>��t>�6̽�>_����G���>��?���?"<?k������=��=e�z?�
�>G �?>r�?�ey>|D�E�����=���=/c;��?�Y?�L�>���=]�%��S�!U'���K����L���>�oH?��d?���>�1y�n�a��8�	�p��Ⲿ>rѽ������<���
>C�+>al!=R�!�gͳ�~�)?��G���пY���Є�'zH?�}Q>�)?gU�����K>�y8?���>����������7�P�ev�?�a�?k@?x%���>���=c��>�-r>`N�s������>�J?�;���)�N�3[>�r�?9�	@p�?'g}�۹?����?)s����^&�D��=b6?�I��w��>4+?��=�j����Ÿw�L��>>i�?.'�?/5�>$f?�rm�*l/��L�=�Ӡ>�]?�a	?;����a>��?-�ʑ�I5	�t�a?��@��@�W?���8ڿ&횿{����j��`��=RO
=ð#>]�����=�=�����:>P�>$`g>�݁>��O>%�>f#1>��V�&�Я��e󑿳�<�v���b�nb����~����b��ɾ)`žv~�,UC�hc����O�i����OL�=��Z?:O@?��?�?l߽�H>Ű���=�Z�2Z�=h�>�K+?u{??>�?�/�=�̟��pZ���s��L��x�`���>b<">���>Q��>K�>* �H)�>�=��j>[��='Wm=�#�=ǬP=@kI>љ>EK�>P�>�@<>h�>�ϴ�51��M�h�Fw�;̽� �?v�����J��0���7��ʧ��`r�=�`.?�x>%��q>п����3H?�����)���+���>�0?9cW?�>���g�T��8>g���j��`>4- �4l�D�)��"Q>kk?i[>Ѡh>��N�����v�h�оぜ>�3?3���1��ll��H'��������>�O�>��߽������z���z�X�=&Q?%Z�>�4��SeԾ���}U��o	>ma>|���o�;���>��4�`ĽYي��S��.��=��>�g?̏2>�Е=(T�>R����b�̱�>!p?>T�(>�B?�]'?4̼����� ���)�ٳv>���>�&y>Ri�=�kV����=Y�>fz>3׼>c���S�[�ՊJ>�퉽P�g�1�@� ��=�̥�]��=䲌=c�.
=�ڰ$=~?4`��ұ���쾤n���rD?�?�=X�_<�t"��F��W���}��?�@	˚?���zV�'P?��?��2��=�>'��>aξCXO��1?3�̽ۿ����	�mx"��i�?7��?Ƙ2�{΋��#l��K>�O%? Ӿ�a�>�����w���E���u��V>���>JvV? �(�at��\���?(�/?Q����ɡ�irԿTˈ���>"��?��?������_�E�a�%?��?��G?G�=���R�u�>��>p�?�O?���>7��B�O�>�޴?s�?�~A>�A�?�6w?��>��m���/�۲�
����=�����>uF�=L�ȾxUI�Ѵ��䈿�3e���0�d>��F=Ab�>@뜽�����Qw=���g+���e!���>�0�>\[>�b�>h��>���>}v�>��o/D��sl�򨏾s�[?�-�?��̾B������>�	�=h��F?ԏ?,�M�M����?�>;�^?V�m?��x?#��>��2�s`��kM���%ľ�y�=QI{>Z;�>���>�Ѿ�A�<�K�2Ξ�b<?�P�>7Dg��G�>��i��կ>��A?���>*��=}f?c>(?�5�>�A�>\;P�����mK��?q��>���>BO�?�A?�оAn!�Aό�ӧ��9D�x#z>��m?�=?�@�<]����¶�����;�$�X>Q��?��s?|v��q��>`~�?�g?w�f?�P>�m�� ��Ӽ6ϙ>v�!?���=B���%�.�O?hS?ڿ�>�ؓ��ӽbPӼk�^���d"?��[?��%?�K�[a���þ�y�<��ir$��	 <�-P���>��>�������=��>:]�=n��5�?�e<�=&�>�V�=�!8�����=,?��G�wڃ���= �r��xD��>�HL>��� �^?xg=���{���Fx���U�� �?Ѡ�?�j�?\����h��$=?��?�
?�"�>>I��s~޾��ྶRw�x��w�[�>W��>��l���ߏ��s���@F����Ž�(����>Np�>�?�C,?K+�>6*�>
��J>�tO���R��Yh��%�@�0�=��f��yiӾ�i��$�ӽ�rξ4Rq��Ћ>dH�/��>
��>�Z>&��>���>-d�=M��>޸w>ŋ>@,�>�|$>�
>�d=�R���+�=3]?�������	��-���gP?�Ձ?��?�;N>*����
���9?�$�?ܴ�?4P�>i�U�\�N����>AЭ>^"i�#?j-�=t��J3>�o��8N��P�f�=�>�>i�L��b-���]�6or�<�(?��:?��M����������=���?=�*?�8)�O�Q�p�=�U�,S�d��]�ݐ���Y%�.�p�Ǫ��@w��\���G'�M1=��*?_��?���Pﾼ����Vj��!>��up>���>�#�>���>��J>�z	��x/��r\�N=(�ҫ����>Bdz?�я>o+M?�P5?=�S?/nR?�@>�>W�����>`�!=���>?4?��"?Q�$?�O?dO)?�@2>*���	��I���	?4�%?*?��?HC�>K*��9���,m���=��q�6�l۟��Ii=V��:�Zǽ�í�\�b=�0R>�X?���Ŭ8�z���xk>n�7?��>Z��>���-��@�<_�>�
?�F�>E �~r�c��V�>���?����=��)>���=������Һ1Z�=�����=+5���y;��f<���=x��=-It�e���1�:��;�m�<���><?���>:>ЖƽD����Q���9�4��>i�> ���r�"�*x��橿:q�f�U>�^�?�W�?le<=o� >�=�ϳ��F��R�ž�T����_=�>���>Y�;?P�?��S?8!?�`(>��� ���"r�j(;x�'?�%?�!�>��f��������9�k�?��?!^��A��"�'�Ao���,�N�>�`'���j��8LM� ����I������8�?\��?	Tݼ�0-��?��g�����.:?�'�>�n�>+x?�B6��<l�����>�
?�d?��><�O?y!{?��[?�CU>{�8����4̙��/�`!>�@?��?��?��x?�Q�>~�>#�)�\��M���� ��!�͂�[W={}Y>!��>V�>-��>���=�ɽbȰ���>���=Pc>�w�>⁥>e��>�w>�u�<Y�G?���>�<��՜�Ƥ��胾�&=�әu?E��?��+?��=�|���E�}<��G�>l�?#��?q/*?��S�	q�=L�ּFٶ���q�P�>��>�'�>��=��D=g�>0�>f��>�3�;_��t8�L4N�T?0F?ѻ=�_��\Tf�~����2���GA�Vc��sjS�Is�06{�wK~=�kg�#���UĹ��<��𪾺�����������^���|�?�q=A��=�>�Z���R!<�?=�Ns=�@<<�=e����*R=������\C��|E;��:=�;%<��'�|�ž�r?e&8?�+?{�M?�Ӊ>C>�q��\>� ���Y
?��'>��������x� ��vy���������q2l��菉>tA>/ˎ��z=�\>Y��=SW�<�>7�==,�>��=n?=�C>� �=�c�=qI�=�s >��>�)|?č�:+����8�q����I?|��>��>I)ľ��i?� >����4}������C�?�a�?���?���>/�����^>�p3���˼��������>Me>�0V��a�>iL�=ԆN��ݜ�.=�����?�;@�d)?�'���7ٿ�I>n	6>L{>�U�.Y/��4g���a��V�H� ?e7;���ȾNv�>��=[o�fD����=��2>{4r=A���\��=�4s�-�9=.Et=�̈́>azE>1w�=6���	p�=th=bD�=C�M>��ƻ$�9�i��ԩ2=��=�1Y>D�>���>��?)e0?l[d?�0�>�n�u"Ͼ�:��A�>�=�L�>L؅=C`B>ޅ�>��7?�D?��K?��>>ŉ=$�>��>��,��m�ar復ϧ�p�<#��?�͆?w׸>1�Q<p�A�F���b>��,Žq?R1?m?b�>k)�#�ѿ �31$��>K����
�?ʾ+m��#�E�)���6->5��>�Э>C�>�ڑ>�>0?�7�>��=�1���=���4>8�=�0�=f��і�*Z��
�=�x=c��+p���r��j㼒�T=���<z��=yk�>c�>���> ��=�/��:U2>IK��r�L����=,c���]C���d�Y�z�C|)�ܤ+�*>>��G>��������W ?�[E>�e>�c�?|�t?��>&+���־����l^�(._���=���=v\��7�a�`���J�ǣо^��>�ߎ>P�>?�l>W,��#?�R�w=}�*b5���>�{������(��9q��?�������i���Һ��D?�F�����="~?m�I??�?���>;����ؾ�90>'I����=���)q�Yi����?�'?Y��>��d�D��̾M��y{�>oCG���O�㵕�9�0���������>�����о53�fb����4�B���q���>#�O?-�?��b��:���eO������cL?��g?�+�>��?&A?�R��U����;O�=^Fn?)��?S�?;U>Dq�=�ڴ�
*�>z*	?���?}��?w~s?��?��M�>���;� >�����=�>-��=�\�=?^?�s
?�
?������	����X��:^���<���=N��>&p�>�r>���=*h=���=�L\>�ٞ>O�>P�d>r�>H�>Vc��r���!?!�>�b�>e.C?�"�>���	���F=�"�;@
U�+�@�<t��"��Os�=��X������j�����>-8����?+ra>3���!?w.��u���C>BS>�Fn�Ʋ�>j�>F`7>��>O��>!N	>ŉ�>:�D>˼���	>���u��K�^��1T��þ��>�r����/�	8��PLF��i�o����!z�Rnq��B���;�{�?U��9�A��g�7�E�?k�e>S�9?m���7�G>���>,T�>uM�O���]��X���d�?rA@�->v$�>�u�?oJ?��J��]�zt���f��w,�d�Q��V�[��sL���W3�ų���c?��X?�xP?�<z�N>���?����&��k\>;�i�	�M��vi>n�?g�����O�(�i'��	���6�=sy]?'��?�h?:*���/o��>E�/?�gD?��m?8)?�L?�����3?n��<� ?�v ?�=?W�.?���>Q�q>s�>��V���<Ͻ��v��l/��O������R>J�>^���q��=.+�=~^b;Y��^޴��<��|!�:��=w��=�Pm=���=���>2�e?A3?A^W>N�,?Q\��Y�{@��B�9?I�n=����=㾢���� �u=�<dd?�?*<�?<(>_�,�G�&��H�=6�K>76Q>�o.>��>�v�݃н��>�5>��[>���=�����	��z���h���&=50->�3�>#�.>пW�%oབOо*����>Г�iO��w�`�X����($�(Θ����>��p?g?w�y=��ܾ�2����$�N?D�?��_?�7�?�da=,L��AH���h��J����>p)��=���ⰿ�ư��I*�!�=R&>訌�=��T��=�FQ�P�žIg���H�@�����R>����>e�Ծ��B��iɾ(�i>�@=W��b������Y��>[?��p<�vI����ﾐ�>"�>c��>�lT=��}>�OZ��o� $����>��>>R=fʾ��[��N-�Y��>�5E?h`?τ?z����r�ڞC��>��OI��M[����??K�>�D?:>���=GZ��D���c�WE��
�>s��>���c�G�+���=����"�f��>��?�| >�?�mS?K�
?|�`?�)?s�?�D�>I���h����B&?���?�=��Խc�T���8�ZF�V�>/�)?��B�մ�>�?��?1�&?U�Q?�?��>0� ��D@�ޑ�>�X�>��W��a���`>n�J?���>q;Y?�ԃ?z�=>D�5�4좾%䩽�P�=�>��2?�5#?��?몸>g��>C�����=c��>y
c?0�?f�o?el�=�? 82>Y��>��= ��>Ո�>�?�WO?�s?��J?���>X��<�3���1���!s��rP��5�;A�H<��y=�~��5t��\�~O�<DȲ;�?��B:�����t�D���޺�;���>P2s>�ڕ� :/>^�žޭ���B>����������K=����=?��>�?[��>(�"�2C�=�G�>}��>cQ��(?��?��?�_E;�b��~۾'"M�@��>�B?z)�=U�l�����!v�Z�_=jwm?��^?��V�����>�m?O�J?�aȾ�E���ܾ$���\N�4E�?�I1?�^�}@a><�?C,�?�:?pǤ�cl�o����O:��w�^��=�Y>�\N�+Da�_9�>�=[?�I�>5<�=mi�>e����Ɉ�/��>�fm?�Ƭ?R�?��z=�I|�X5����Y��Ǜ\?2;�>X}����E?�Tw�Uf��鮉��"����]Aʾ�����o��2��U���L���0�ӏ=�?т?X��?�oN?����t���z��_���,����Q�C-Z��I���D�c�r��t�ٴ�����᏾=����?���?R'?�>-��y�>�l�������;L�M>ә�:���t�= ��m�U=fPf=e�q��9�O<��?系>s��>�6;?h�\���<��G5�U�5��&��*>x��>���>��>�`����/�h��m4ǾD~�I�Ƚ��t>D}c?��L?��o?������0�a!��8���gQ�Gg����H>�
>��>}z_��"��M(��S>���p�(����Lm
�	`�=�_3?�h�>���>0�?N>?G��G��� #v�|Z0���X<� �>ӄh?���>(�>��׽�l �(��>St{?mC?K�u>L���j�O+���\;���>�@�=#�?��I>���Sk����������?2�s�>�|?q����HȾ�S>�8�?W�1�xhk��,�>؞*>S�Z��Y_�[�^=��z>�3�>�h�=c�>���}��+2k�)D[��O)?nK?>蒾 �*�5~>%"?ŀ�><-�>+1�?+�>~pþ�D�б?��^?+BJ?qTA?aI�>-�=���G=Ƚ��&���,=ه�>d�Z>� m=]z�=����q\�gw���D=�p�=T�μO����<!�����J<���<_�3>L�ؿ��>�����pP��Ҽ�����u��!������tǘ�Jw�/����x������2��cu�*�?��ֈ�#^��p�?{y�?}����T��g��-rk�wG��1�?R����Q���@�v�!��O�����X�ľ��0��"N���b��d���'?������ǿ����=ܾ� ?�A ?��y?��Ý"�U�8� � >�/�<w8�����њ����ο���'�^?���>F�{.��Z��>c��>z�X>Cq>���h鞾��<��?H�-?���>ǔr�g�ɿꊻ�a��<���?=�@u|A?��(������U=��>@�	?��?>�B1�	A�(�c�>D;�?���?��M="�W�Z�	��e?�<��F�%�⻄�=w^�==���ƓJ>`�>V��AjA���۽9�4>)�>�"�f����^���<��]>�ս(���؄?��a�
�c�A/���|�Z�L>7yY?�?�>V_�=s/-?3�Q�L�ο�O�o�h?*6�?mv�?� ?IpǾ�O�>��پ݃R?��5?���>�h"�ci�{�>%����==D��@	Z���>^��>(�H>o9!�������O}��p�=F:���ÿ���n���<=�Qż�ڈ����ͱ��`�oe��D!o��@ĽT�=5�=6�U>�E�>fuh>��u>%]?�"q?�Ӛ>��>}-��ݙ�����=PҊ������f��:�_����J��߾;���~����4Ӿ�?��y\=�k�71�����&�d�R)�K1?g*=�1��
%���`=)sž�Rv��f}�*�$�[�����%���[���?�h.?7x����8���$��y���S��t>_?Kw��Դ�������J>	μ�=�G�>�:�=,�������V���3?�r?���{��'k>�����nH=��)?��	?�(��:�>o0,?���w*��;�>�p>�E�>�z�>5<нl;��^ٽ��?4�l?�SȽzZ��?��>Ό�ʬž��o>�a0>�񪽟`�=��=>�Þ�־�f�Y>'���>�(W?}��>��)��aa��v��dY==��x?��?&.�>q{k?��B?�֤<h��}�S����bw= �W?'*i?_�>���{	о3���A�5?�e?��N>�bh� ��.�.�ZU��$?�n?-_?]~��#w}�w��n���n6?��x?��~�#���뻾x���w�>V��>YK�>#C�?`>?,\Z�sD��X뺿3�;�5H�?��	@9K�?�-�=�D�i��	?�b�>'u������x�����5q=uX�>�A�Vss�e�B���j��Ib?a��??*K����"��q�=�K��I�?��?�����|�<���@l�������<9��=n;"�Î'��h��7�9�ƾ��
�[ݜ��6��]��>�R@o�߽���>��8�(E��bϿܵ��:UϾ#�s��?Ù�>�˽ki����j��t���F�J�G�������>��>����c&���{���<��j�����>����y�>��M��(���t��5<���>�j�>ߨ�>h5��F���"�?Y����hο\���k��-�X?�?�Q�?� ?��;%S}��s���vFG?Ӗs?��Y?�T5���Z�M	Q�%�j?�_��xU`��4�sHE��U>�"3?�B�>T�-��|=�>���>g>�#/�y�Ŀ�ٶ�9���Z��?��?�o���>r��?ts+?�i�8���[����*�J�+��<A?�2>���I�!�D0=�QҒ�ż
?X~0?{�f.��d?�zy���i���1��.���>�@���!������+<a�x��(���P\����?2�@���?`"ֽ��&��6#?�Ɗ>�i��,����=6�>���>�w�>@�=���>�s�6�Z���>��?���?R�?<?���[���d�=X�y?���>!��?M��=�X�>�=)��������!>\6�=`;&��?,jN?���>݉�=��:�^j-���B��bQ����D�\%�>%da?�LN?�8c>a����.1��#���нc>/��-�`j6�i�N�e5>��;>'->�G���ʾ3$?D93��ӿS]��p�ݽG�3?��>�� ?^���̴�f6>��M?�1�>�&���k�����i��*�?�|�?\�?�� �<�9>�?���>��u��A��~�?�o>4�;?r��F\�@�[�CR�>z^�?��@.��?�T�9N?��n_���k��Iܾڷ{>)K6?W�����>�
?���=y@e��6���Q{�}W�>�'�?���?�?g#f?@t�M�/��Z�=��>�e?��
?O�@<R���X>�d�>??�����D� �i?�@ה@F�]?�!���kֿ�����L������j�=���=�~2>%ڽn@�=I�7=��8��s��]��=?�>��d>N q>�8O>\p;>q�)>�����!�.n������� D�u�����Z�}���Hv��x��5��6���x6��2ý)�����P��4&��`����=�GU?RjQ?��q?p<�>�TY�L�$>]�� O=��#��q�=j�>��2?��K?��)?9��=�1���c��N���Ϩ�����q��>�F>0=�>n��>H�>��!;ݗL>k�:>��~>�+�=�Y4=Q;9�=0�K>Bϧ>���>���>HA<>w�>.д��.��נh��w�
̽ �?����ѴJ��/���/��'���r��=T^.?s>���a>пi���w2H?]���@$�q�+���>P�0?�cW?X�>d���fT� >ֺ��j��h>^ ��|l�n�)��Q>9e?��g>�V>:�F��o ��-t�DLȾᥝ>ou=?���M���mL|�Z�%�e����T�>�S�>]�t�@���� y���w�G>��E?��?��ּ߽ܾ�2!�������M>�t>���&�=V�y>�Ɲ��y�2R���D;��=v�>K3?Ę0>�m�=C(�>�4��$�Z��i�>��?>�,>�3@?_0&?�¼&�s�̂���0��Dw>k)�>�{>:�>��U����=�z�>�yq>�X��qW���KO�/�Q>�)s��c�gF�c��=����=r��=+����	@�v�m=�
?�.���|��N���=.�J�]?�0?�~<�6�=y�#�ĳ�Iվ<b�?v@�۬?dϾ��a��1�>��?�K%��_�>Q�?��t>��%���l�?ƀz��57�-7�ʵ;��ܲ?�S�?ɀ&<�]����o���=�~$?ȶ�3��>�^�ч��U+l�Z;��9uh�c�>�>?%d�Z�=Y����	?�>����笿�MǿN�g����>���?I��?�Ǒ��3����F��~$?� �? �B?�U>+㺾�$�V$�>�/?�W?���>"�)���׫?�K�?���?�y=>S��?�?���>�먻�@,�$B���j��ZT'��=��>Ȩ�=V�¾ZIR�g��ʏ��@ib�D"��	}>t��=���>��=��ð=���l���RC�;��>��>]�T>Cw�>���>q@�>�W�>OZ�<lk!�����&%���aY?�y?�n��.���2G>k><\�E�J!L?�o�?�叾�(ɾA�?>�a?�^?l�Q?�?�g5�w\���ȿ�fؾ��e=�a>���>���>0v����;�A\��AA�>��?�!s�2���ң�d�(���>�(E?n��>��[��t?1N!?���>���>F��������?���?�n[>��>�`�?�k)?¤=����n(��+ײ�|�O��f3>�Vx?,M?DT>Ip��$���h�y��`��>j�?�J�?�������>֘?O�q?�
x?��>�A��i����Iq�opH>�!?� �P�A��C&��l��q?#P?���>b��Jս��׼�������?�\?�4&?&���9a�Bþ���<�� �x>H��e<�G�M�>��>�D��Gܴ=�>>�#�=Am�)6�7li<Bʼ= h�>���=�K7�����0=,?��G�}ۃ���=��r�?xD���>�IL>����^?kl=��{�����x��	U� �? ��?Zk�?b��@�h��$=?�?S	?m"�>�J���}޾6�྿Pw�~x��w�\�>���>*�l���K���ڙ���F��Z�ŽH�5����>�^�>Kq?�-?��>[��>����9�F�t��]D޾�}b�h�3�d�.����z��pоAԣ�(�ܽ52׾i}����>�rN���y>�_?Y�T>Q�y>�>�i=I��>n��>ڌ�>C�>&�C>Z�L>��=0�׼P2׽��R?Z��F '�n��深���A?z;e?m#�>Ib9��Å�ޘ���?�ݒ?䡜?3�~>�Tf���,��W?J�>Y{����
?cC.=k�L��<������r��E=�#�>�9ڽ+h9�Z�M��h��?�m?	�R���;�H��`���r=4Y�?�*)?��)���Q���o�A�W��S�A���g�-�����$��p�KƏ��\��Q��ht(�{,=�h*?�?*�1��	���$dk�!?��5g>g��>�W�>ZY�>}H>A�	���1��^�F'�oƂ����>P{?��>�K?�",?�h?A�B?V�>W�><���S!�>��;=ӈ�>��+?	�c?J�?>�>	?��,?7�=���<P��u��U?U-?9��>�-.?@]�>�CվVg<�&޽K���G�|D��=��=i���.�ʊ5=Vy�>�X?�����8�����`k>z�7?��>Y��>���-���<f�>�
?G�>> �~r�c��V�>���?}���=��)>���=F�����Һ�Y�=H���*�=d5��z;�+d<���=s��=QIt�f;��W0�:g��;�n�<���>%f5?:��>�d>�������m0�=d��>Y3 >���=����#`~�{#���@r��RH>���?�d�?�d�=U��=�E�=�
k��Vξ���r���$��,0?�^?�V5?lK�?��V?��#?TI�=>2�츎�xm��
���J&?5\?�֎>���ٜ��̵���K���?ٌ?�U�*��<�94�}̆�����O>ޠ��󀿩��1�Y��o�|y��X����?mΓ?�Z��EC� � �>ɕ��S����&?g��>�>���>��H�
�i��n&�N,>��?��{?v!�>}�O?�={?��[?(qT>c�8�G0���љ��4���!>"@?}��?a�?8y?p�>y�>6�)���L�������߂�)W=|Z>i��>�*�>��>���=t�ǽX����>�gV�=�b>o��>�> �>~~w>�,�<�G?��>>W��0��@褾Ƀ��<=���u?Λ�?��+?�T=ԁ���E�fI���D�>�n�?S��?q4*?��S�m��=`�ּ`߶���q�%�>fӹ>@4�>p��=�VF=.n>��>{��>�$�a��q8��pM���?eF?n��=��ÿ�6n�ep��4U���SO������\�%Si�@lg�!�=`Տ��,
����� FM��^���%�����$���OC����?�|]=0X�=��=xA������x^<�MT=b�<���=~��ݴ<wX�D���b#��ؕ�;�ӧ<w)0=Oܼ0*���7q?��:?Q�@?0E?��>��Q>�x �.�Y>�L���,?�<(>���Rm��=7�����ȟ����Ծ�艾w'����>�<K�!B�=K#0>�9�=e�9=�0�=3eK=�s�=z��<�U=��>��=�.�=u�=/Q>e>0|?���� X��1�E�.� �WmF?�>�>��>fl���W?3&>ۀ�?�Ŀ����?4h�?���?�?Aꎾ��J>��l�v����?�}|b��*>>=>��B���>��`=�!+�pc��RW���{�?�@h�*?�˔�2�ֿ�� >��7>s>��R�܄1���\�8�b��oZ�A�!?�I;�7̾�3�>w2�=B7߾�~ƾ�Y.=8x6>iub=���T`\��,�=��z�(<=�"l=���>n�C>���={'��^�=�{J=[f�=6�O>�����k7�7�+���3=���=�~b>��%>"��>P�?�b0?�Wd?5�>�n� Ͼ+@��J�>�=2C�>�υ=�nB>ዸ>��7?�D?i�K?a��>/��=��>��>��,��m�5k�!Χ�ꁬ<��?oΆ?�Ѹ>$�Q<��A�#��!h>�a2Žxv?yS1?pl?V�>B/�Wտ@K?>��霼�T��[�⽏�پ�t�67��s�U�>�g���<%��>	T�>2��>�y�>�2�>M��>�[�>g�=o�Ƽ�c��#�������>,�ɶ>������N<Q�����SA�<��n����.�y�����9-��'=�4�=��>ds>���>��(>���6�B>ƣ���N�"��=tH����K���f��py��$�:�+�#�>�m(>�Vr����H��>�S>α�>�
�?I�r?I�>���;�쾧���>����W���0=�m@=	���x!7��]���P������>�ߎ>t�>Z�l>(,�.#?���w=b�lb5�S�>|�����)��9q��?������+i�Z�Һ��D?�F�����="~?R�I?C�?Ӎ�>����ؾ�70>eH��g�=��*q�Hk��_�?~'?���>��!�D�&2̾�6��^��>8�H�8(P�T����^0�a���K��\�>L���о�*3��;��e4�B�NBr�y��>�wO?���?!Md�
^���*O�*��s����?3?g?���>�D?eW?N����?��R��T�=�wn?�s�?�1�?b�>��=H����H�>)�
?�!�?]-�?�Ps?ۻW��w�>�
�<��%>�����Y�=�>��='��=;�?.�?�?}u��;�ơ����tq��I=VD�=��>�[�>�ށ>���=��=ƹ�="h>���>ᔔ>��b>�9�>��>)���v �΄?�P>�R�>�R?�i�>���nR�Q�	>��<�Y]���f`b��k���=t���c摽ln�W��>㷿$��?��>tc��?����_��Ԏ>ftd>�<��)]�>�~>���>�i�>�A�>��=�l�>}�%>&Ǿ�?>�L����<�d�%�o�
ȵ���>@z��Q$�����t��^���хľğ	��z�Yt�n�=�ϻ==��?I���[�]^$��H4���?�*&>��?�ݝ�-����>��>]�">"�}��������nϾ�ؘ?�4�?A&%>H�>R,u?�?�W��YͽNQy�+n�����d��S��x��x�y	�yZ���@?�I[?�oH?\����T>�x�?�B�3׾#�>@�S�R.J����=���>rB��/Ͼ�D�dX����ž>�=�G]?�8�?�RN?X����q��U�>�,4?��~?q�S?R�+?^|B?�R���EA?���=Ģ?P�?W�@?�O%?��>��>��9=�n���O=&lb�횾nt@�5fl�P�?���p=��=6}7�	g!<UD{=4�r=�.��=н�0�=M�L<��:�O2�'�9=y �<\��>��u?�l?�P�=d/?R�G�"=d�]=۾�(;?�O�iw��g���͹�=�3����ٓL?��?��?DP>�w*�.W���=RR�=z�>��>X�}>�\���w;�z>_�[>���>m�>d�ؽA��V�ı��@E=�|�>��>�H>6����hc�����������>�2վ�����!�0ꉿo4��o.�]�?�g?�Q?����ѾQi�=�v����F?��?�J?{}�?� �&\��C��p�=�;P�>��0�ڃ?��6��.׬��<#�Ԕ�=��.>R���c���]�~>�+1��B��s�}����Mɾ�Y>������> �V)��򣕾�S(>NZ1>�+�����W�H/��.v^?��X<?���5Q�Y)��%�0>�Y�=l8>l5�	d<i�?��_�+��>B��=ؽ&�����%I�n
��"�>�x>?u?I��?�C��y�p���N��<��(q߾ZUY=,'?��>r�?E�->"���R�վK���j�_�-���>���><��8�M�lK��Ϩ���?���>�?U1>>Vu�>؇<?,u�>�s?�*?fL?�Ƃ>Vl�~�ɾ\�+?C=?��x=�7���s���5���5�ot?��5?�׆��`&>e�?@@%??�3?��V?@�?�="��XN��g�>C��>�m��E��-��>zML?F��>j�M?{��?�{>%z=�%����ӽ��=�9O>w�=?� ?�y?p+�>���>�"��N�|=��>��b?�M�?~p?��=�x?>�4>F�>}�=}�>(�>�f?�|O?as?��I?���>h��< ���ٰ��,x�{f��\�;���;��x=/����{���n�<�'�;导�񉼔��[sB�����<t��>�Ӕ>fi{�g=>'᷾G=���}�>A�:���������\+)��vP>���>	?)��>t<0���>@�>t&�>�G4�
t0?7�?�G,?J0P��iG��̾�H���K�>��L?�s4=�fe��ȑ��+l�Y�=�Rq?}2\?ɞ��kV�>c?]?mA�,�=� �ƾZrg�7>��}R?=?;UQ�'v�>��|?A�r?WF?��[��nl�����P�b���x����=�ݛ>w��?rg���>�8?�g�>�d>��=����z������?�Ë?8�?�}�?��)>B�k�X߿A���샿�YP?�G�>����:?�`��	��k毾M�X��~��Do;�P�L쬾������KN��66!�1�_<"�
?�'a?ֵ�?@�F?�u��[�}�����q�;9M�r���G���5�zeB��B�]����%�>���]�/��=>�|�eW?�S��?TM'?QU*��%�>yp��@r���qо��F>Q������v=G����W=��v=�Ik��4�L���z�?��>���>��9?@f]�{=�P�7���6����X�">7D�>���>���>t ��xyA����d�ɾb���PȽ$l>qX?-�z?r�?:���05��W���*���_D�ټ����>��6>Ck�>�l�����J�D��7��d��)��ǆ����<�=�"?�:>�c�>pG�?,)�>�$A��y3���Óf��8 ����>;4=?T)�>kY�>;ƾa ���>ՙ?��4?J��<n�Խ�=���� �<T�'?q��>DJ?���>ojh>t����`���]����q�m�(>�;h??K.�6_Ǿ��>��r?N=��Ƚ;���]�>M�"�+54����h��>��>��h>mN>�����R4v��f��j1)?�D?���a�*��,�>�)"?�7�>Tʣ>~��?
��>C�¾���8�&?�J^?3J?�JA?���>zC=>��f0ʽؾ&���1=Jj�>A�Y>�n=�}�=�j�5�]�DO!���N=m��=��ʼ�⸽Q��;���"Q<	
=[R6>;�̿e$-��a����1j(�yXA���ٽ�>���drS�۸���X�2<����&^:Y}2�\�V�#�X�w�5�r�?a��?I���XX<w�� ���2�����?,����=dMf�z/�ܨ�o�Ѿ(7I�k���A%�3�>�g	a�7�'?�����ǿ����	;ܾ
! ?zA ?:�y?O�	�"���8��� >bG�<�(�����˚���οB���
�^?���>;�1��1��>��>O�X>$Hq>����螾�/�<��?��-?���>Ǝr��ɿ:���ͤ<���?3�@}A?��(����a�U=`��>ێ	?r�?>UJ1��F����U�>Q<�?���?0�M=�W�Q�	�~e?�<I�F��B߻��=�E�=�r=T��a�J>�Y�>���YA�?ܽ~�4>�څ>�n"�Ū���^��R�<�]>�ս$��G��?"l��VK�ԝ1�Ve��'ϲ>k�V?B�>kv>(?HY���Կ&�v���1?p@���?W6?�þMd�>G��eMl?t/?��c>(�T��~�|>�>/LW���>�U׾V�~��}�=�'�>���<�T�H)����2I&=�Ri>*��dſ1�#�9�"��kC<�G��d��c����;<���k���h����sf�=�o�=�dM>2f�>v�Q>3�]>�W?}k?��>�E>�G�h���Qƾ��<xy� J��W�����j.��]&��ܾ����t��*�W�ɾ�z=�..�=w?U��̍��%�� j���>���2?� )>~ȾN�I�P�P<�/Ǿ����A�@=���dƾ�l-���j����?��D?�����5L�_Q�eu�M�ͽ�2V?N������f��:��=���@��<%�>X��=o^۾Ϥ1���U�ގ6?&?%����P�G&�><�9ܸ=��-?u�?�ž� �>3�B?�gg={ژ=(/>G|�=�Ď>K?��;�D��Q
��F?��_?�it��Ȩ��?��龉W��b6ý=�>)ռE�0>{��>8X��jѾ��2=L��k<�>�'W?
��>��)�,��_�����L==�x?��?�/�>6|k?k�B?7�<�g��R�S�u ��Mw=��W?�)i?'�>.����о����?�5?k�e?P�N>�`h���龁�.�?T�%?��n?^?�~��ov}�$�����o6?䙀?dt��dj��갢���K<W��>!��>���>��B� ?L�8?Dl�����绿 ==�?�?�[
@<��?4���=b9L�1T?���>~�a�XǸ���=�#���&E>��>�ξ~Og��0����Ќe?y�?i?�,��(����=�֒� ��?
=�?����"�<[��mm�y���Y�<���=$�E�U��X�� �7� Tž�j�{���������>'O@�d��c��>��J��kῥ�Ͽ���`�ʾ�w}��d?Y��>�]������Ln���u�.XC��-A�������>��?>��=�Ns�ڛ��N�7!���"? �ýSEp>�,������o��fI>��[>��}>A<>������?�ѾZ��-���a`����A?ç?�Z�?��l?FX���-���ٽC�>�)d?l|�?��n?���0q��\V��$�j?�_��vU`��4�lHE��U>�"3?�B�>T�-��|=�>���>,g>�#/�v�Ŀ�ٶ�,���X��?��?�o���>q��?ws+?�i�8���[����*�x�+��<A?�2>���H�!�D0=�PҒ�ȼ
?]~0?*{�f.�h�_?B�a�:�p���-�w�ƽ�ۡ>��0��e\��M�����tXe����Ay����?P^�?s�?״�� #�46%?��>����8Ǿ?�<��>�(�>c*N>hH_���u>����:�jh	>���?�~�?ij?䕏�����U>�}?�G�>J��?��=,��>B��=O���>g�=�V>��=����>�5X?$h ?�y>n 6��,��i1��BG�IN��pO�U��>�Nb?`V?-G1>�������45�� Ľj!ɽ�v��i?��v�����->o)R>IE>�M����þ�&'?>q6���ۿl4�� 3��R�C?�Z >�H	?�Z(����ǁ�=UOB?Wd�>�Y��4(���ד����?�c�?az?�Y�� �=���=���>�`Z>�ˡ��F	�)�2���>
\V?��@���Ds���}>��?Ǻ@pY�?f�x���?�d�b#����s��C�i4	��B�=�t7?EB�$��>��?�@�=�m�����vz����>��?b��?і�>Aj?��t�t-����=f=�>"�Z?;?�v�h��%�i>�?	U��f������_?G�@�@0yZ?ꦿ�hֿ����\N��v�����=���=��2>Aڽ\�=��7=s�8��I��U��=��>�d>�q>�'O>�_;>t�)>����!��q�������C���"���Z�9���Vv� z�l2�����I@���0ý�v���Q�Q1&�GF`�?B�=�T?��N?a�p?8?]J�c�.>^ �r�
=����o=��>��-?}H?�+?�=�띾��d�7r���ר�<Ն�K��>2�D>�v�>���>y$�>�%�;5PG>�X@>
��>ql�=L�1=�i8;�=��T>��>�,�>ٺ>L<>��>Ĵ����ԥh��}x�g̽��?�;���J��1��y��|���Sߠ=ob.?">����1п����<H?�0���6���+��J>1�0?pW?�>�����V�<:>���;�j�/>Ѐ �E�l�*�)���P>_?� f>��t>�3�p�7���O�+����s~>�Q5?m궾w^6�:Su��H��޾�LK>͝�>�_ ��1��ؖ��	��*i��`x=ú:?��?+�����ņy����O>!Z>*�!=s�=WQL>0�`�3�ȽդG�`2/=���=Qx_>�?��+>C��=�>[>��S�I�8�>��=>�*>�f@?Tg$?ϸ�2��:Z����(�f5z>C�>9�~>>c>&)J��=�=�	�>��^>\v��~�#���k?�('S>�����Z��큽.�r=✕�J5�=��=�,��P�:�z+/=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ��>Ygf�� ���\���i�:��=�ތ>X�P?�D-�����cq��� ?X ?+��k���5ͿZ.���?@��?�6�?h���OW��w�M���'?c>�?\0:?�f%>���wL>�1'�>1?(e?��>�I'�=h��h?^=�?x�?r�/>���?�;w?��n>�"���c��W��gJ|���>�_�>�C�>��2�:�J�ԫW�f��?�����a�ج��<�>�>=<��>��齨�
>��N�����<�3�>w��>`x>�&�>#�
?�b�>m��>r���xC�������&��V?tǄ?1������)>�]<k�z�5?@wZ?�~\�Z)�Zo�>;M?F�}?T.P?��>2b�C��t�ƿ�T¾�/�=���==Y�>�?��2=[�<����|��Ä>��?hJ�=���˾&& �+ܞ>#r?j?:��=��?�l%?�6>�t�>�D�2��4	G���>Z �>�?-�?��?�S��7=4��\�������Y�2�W>�zw?��?�+�>�c�����G����y�?�w��G�?Wi?ҳ��ʧ?(I�?X�@?��C?�d>�A��t߾^}��7|>�=?��
�B�@�"��   �*�?k5?P�>p��������<�=
������R?	^?L9'?
����`�;|ʾF�<�s���8'u>��?����$>x >�gv��=��>��=a�s���/�`D�<|8�=�6�>I��=a�+�v�n�3=,?boH��ۃ�И=��r��tD���>�:L>+���[�^?Q�=���{�����u����T���?6��?�g�?����h�l(=?��?�?�0�>�M��σ޾��qtw��mx��w���>&��>F�m�9�ݐ��:����C��+ƽ�7 ����>�>S?&?���>�0?\���E��]���,���Y�A���L�n|��nھG�� ȡ��b�����e�9���r> {�a�x>���>]�>��>x��>�c�=��>Q��>NS>���>��>��V>��>|E�.�νODR?Z���ا'����΀��B?!d?�(�>2oi������B�?���?�q�?�	v>-sh��
+��d?+.�>�i��f
?h�;=����<�?��m!��/��{���Ԏ>��׽v :���L�`[f�T
??������̾^�ֽ?$����=^��?s
*?��3�O�'�dOt�X�_��T�g�K�V��^`��A<��o{�S��� �u�fz{�J���<��?X��?�鬾��վ1ľGjv��QN�Z
o>��>X�<>��>Ӊ=>�{վR�F�Pi�K$&�% ��N?jx?��\>��a?��3?�]y?��P?�b~>I*?]�w#?���}>3�?֬5?�0:?v�?�r?	�(?t��=�Z�<�����@�?�G	?�,?�A
?�ѻ>����pۚ;,N�=(K���b[��/ݽKH�=#z�=�L��P�O�5y�=��>�X?m����8������k>k�7?��>d��>���-����<|�>�
?�F�>; �~r��b��V�>���?����=��)>���=ߎ��i�ҺZ�=������=�6��\y;��d<���=E��=Qt��%��8�:��;�o�<�>��0?��>�cZ>������ݾ(Y ��`P���>��p>ϧ�>��	���n��T��w�m���=�v?r2�?>�>��y=k�=>�(�����8Nھ�"ƾ�5�=�D�>YW)?���?�#�?�?\?�h~>|P�Z��_�A]<�Q,?^!,?��>d��j�ʾ�񨿉�3��?.[?v<a�Q��Q;)�J�¾��Խ"�>�[/�%/~����D�������~��-��?ؿ�?�A�2�6��x�޿��\��?�C?�!�>�X�>1�>:�)�v�g�j%�2;><��>HR?��>��O?!�{?��[?hsS>��8�_?���7����r���">�J@?T�?�?^hx?X��>��>��)��$��=����]���������Q=]�X>�Б>���>S�>���=����kή���@�s�=�?d>O�>I{�>���>��u>���<s�G?���>�]�����褾�Ã�M=�q�u?���?g�+?�X=׀�&�E��E��}J�>o�?���?�3*?��S����=��ּ8඾V�q��$�>�ڹ>�0�>]��=�jF=�]>}�>��>(��`�\q8�[M���?�F?l��=tdƿ�tp��Vw�%���Z�k��[���``��Ɠ��pW��I_=暾0U	��/����A�{����[��lE������Zk�?*��=몳=��=��<����=��=���<�%=$��ܨ;1a*��T����� ���t�;��P=���v�ʾ�x|?A�G?m�+?��C?D�~>0� >W:H��>ϧj� �?7T>��d�/�����4��٥�{��i�پ^%پ��d��ԟ�v>�iR�"!>��4>���=-��<��=��s=���=����wU=/&�=��=��=�)�=�>p>'�?Å��1Y���:��э=��O?�:�>W&>SW���Y?�b.>͇������Z�2ʂ?�c�?��?�x�>�?�'j>����=�O���Y��U�>]d�9�𽃟�>p/�����7��_%����?���?�W'?�}���@Ͽ�/
>!�7>��>�R��~1�K[�k�a���Y��i!?!�:��̾s�>�l�=�!߾�uƾ�%1=�7>
�a=V7��t\���=@L{��==�Kl=Ǒ�>D>�ѹ=<���~�= �F=��=��O>䍻�S7�b�,�v�2=tT�=?�c>W�&>���>��?qb0?�Wd??1�>�n��Ͼ�B���E�>��=�E�>aυ=�eB>=��>~�7?��D?��K?Ӈ�>ξ�=��>��>�,�P�m�^h��Χ�?n�<ߖ�?�͆?�и>�Q<��A���zg>�G0Ž�t?5S1?�m?e�>%������T�i'<�ݚ��U�=v�������w�����q��n���kӅ= ��>Ͽ�>"}�>�?5>�[6=?��>a^�>�7>kJr��V��-�ɽ:�l�P^�=��j>-,�<����C��[�=�ǽ)����������(2��@=��'����=��>y��=9��>�>薆���E>e,˾��Q�7�>ިྙO���m�^����#�����j
>��'>xB������?�B>ll>�?b }?��0>p�R�(�C���dY�Q9���=]�4=
a�P\>���k��M��Gؾ���>��>��>��l>�
,��"?��w=⾾a5�	�>�u�������6q��>��5����i��g׺�D?nF��4��=� ~?d�I?�ߏ?��>9���ؾ*30>�@����={�z/q��g����?d'?d��>�쾜�D��;̾�׾�	 �>YI���O�ʽ����0�����䷾:��>�֪�D�о�3��f��������B�G@r��Ӻ>n�O?��?ab��T���UO����逆�Ds?"yg?�!�>�G?�7?�K��dg�g\��K��=��n?���?�9�?��
>Q��=ԝ��k�>�/?%�?]x�?��z?Yg����>:wi=8�>I���#�i=֪�=J��=�>�� ?ί�>���>�����M	��@�B.�J�g�L=S=?��<��>�n>Ϗc>�>�R�<9x�=�l>��>J��>�T{>p}�>�q�>Ԏ�������?j>Sj�>ң;?>�>���;e�ʽB]�=H�_�T�gU� 1�A�S���=��,�o,�<�����>�S��F�?rT.>
�-�?���4�=��&>�p>ٌo�E�>5�(>j^|>sē>M��>͖>;6�>I�=>a����>f�#�]���R�|\j�� ־���>�缾�齘j����Fmh�u/�����dp�@|��>�<��眽�?���_^��j$��k���PF?d+�>��"?C�ʾ�r+����=�?�߼>Ps��󘟿o��h�$�?��?�ZX>>S�>�^]?�?�z]�;P�7\a��v��^<��`��RO��B��!:��qM����JR?s�l?-DC?�e�<�D]>gJ�?t�������)�>ʶ4��}5�<�=f8�>�E����S�ݢؾ>P���Q�ʢ3>�|a?�b�?%�$?��'�?Ŷ>m~.?ڢ>?�9�?�'?�/W?X̜��u0?Q��{�>ԽV?��#?��T?��>��>��b="�<���><n�� - �!*�Όн�B/�>�};\���>H=��I�����<k���'��WIW=T��	>I�<!�0=@�=p��>��]?BS�>�u�>U�7?��x8�|ͮ�t/?}�8=-v��� ��Ѣ��R�l�>��j?�?�gZ?$d>�B�ׁB�+><�>��&>b�[>@Z�> Cｈ�E�#C�=�>k�>�k�=,M��ā�A�	��k��30�<�>���>�>`p�*f>*ܾB�G�1s�>iٟ�����⽟M}�زG�3�־�V�>y!T?�.?7��=9/оD��ㇿ�U<?+?f�X?��?l6�=���Cv�2^x��ˍ����>�J=G���f��<��,�X��P%��0>�c޾Vݠ��Yb>����p޾��n��J����{5M=P��SV=h�O�վ?2�פ�=''
>����� �	��X֪��0J?Фj=�w���bU�<p���>Ⱦ�>�ޮ>Ѷ:���v�o�@�����7�=I��>�;>vW��E��p~G�H8�x��>WC?��k?�Z�?�g��a�j�����A0���L���i<���>���>Ba?��f>->�ꑾ�]���j�~3>���>� �>�]+���M�0Ã���پ���g>v�?���=C��>b1?ys?�Ň? /?���>��_>�����s���%4?���?Zq�=>�&�'G�~u5�k&B��6X>�F?xx���=V��><�<?�b?O�q?��?eoj<��"�.�L�:�>*gk>ܰh�-�����>uA?�>��v?ɒ�?���>�z?��/���F�b>�>�3?�(?�?�G�>���>�����=ޞ�>�c?�0�?
�o?ۂ�=<�?b:2>4��>���=뛟>k��>�?GXO?$�s?��J?���>n��<�7���8��KBs��O�tĂ;�|H<z�y=ؚ�b3t�"J����<!�;�g��eJ��Y����D�'������;d^�>w�s>�����0>��ľ�P��<�@>���]P���ۊ�4�:��ط=�>R�?���>�W#���=��>bH�>���7(?P�??�!;6�b�C�ھڬK�?�>�B?��=r�l������u�th=��m?ڋ^?ϔW�$����b?��]?�G��<�l�þ��b����O?.�
?N�G��۳>��~?��q?���>��e��,n����TJb�1k���=�p�>�h���d�I�>֔7?�"�>c>���=�d۾�w�-����?~��?&�?2��?�1*>��n�H+࿓��^��{:`?�i�>F��W�*?��;��̾����叾LGϾ�֠��(���	�������p�*���ҽ�ة=��?�Yv?K7j?U	g?c���GHi��@^�������P�y^�>���E���@�^mB��;o�9��j����ٝ�!Fb= �k���Y�Xo�?Ȥ?�Ȃ�ͤ?��k��)۾�ھT�$>V�K�V���A�=���|�;v��=&�L��h������?"��>~��>^'N?9�H���>��%*���D��뾧o7>���>���>#�>�{���_�ν�ξCԓ�S����7�>��c?Bn@?��w?#냽͋)���b��i����
��}V>P&�=ެ�>9���F��*-�*T?���j����5s�����">s�8?�^(>z��>��?	�?3�������۾5��<L��>��s?��>�:>U#��I#�q��>�e{?+��>L�>a��a$�(��u�����>|'$?�.?O�Ƚ"���%9�zց��ы�z�(����=]�`?�/P�b�7�#N3>��G?
�=xx=$3�>N���
4�Q�
��J$�C#>�(�>n���D>g����N���}�9���y�,?�?k��T;!�{<�>�#?Ӛ�>�"�>5o�?V%�>p�žM�μ?}?h>b?0P?d@?i��>�e�:���0̽�"'�	H=S�>|�p>�=�>�G(��v��/��j�=�u�=�<�������L��Rμ,��<��5=�:>��࿴L���\�F����D~~�9V�SAA�>:��ʾՊ���j�F����(ͼ.��Nku����}N�(��??l�?B����������py�O&�۰�>5%����!r�(/h�;��"�پ�b�d�7� `Z�e�Z��mE���&?�q��>�ǿ-����Qܾp ?��?��y?��e.#���7�-$>���<����$��a̚���ο�#��4e_?���>լ��쥽ȵ�>�P�>4Z>�%r>+/��Nc��	J�<�?�-?!3�>�Xq�0gɿ88���>�<&��?��@hA?�)�HO쾖�T=EJ�>��	?�5@>1��Q�������>�7�?��?!�K=#�W�^��9le?�<��F���ػ���=G0�=��=��~J>e9�>T9�q>A���۽�b4>�ׅ>F� �����^�?�<6$]>�pֽ}���Մ?"{\�^f���/��T���R>��T?A+�>;7�=ò,?b7H�2}Ͽ��\�+*a?�0�?	��?��(?;ٿ�ؚ>��ܾN�M?�D6?f��>ce&�*�t�0��=�AἭP�����L&V���=Z��>�>��,������O��X��{��=`7���ǿy�+�5�D=���;Ϙ���[s��<�:*"���\����a�ڽ���=T�!>�w7><*w>�1>�R>�bW?��w?�x�>Z��=��,�����t��m�GՌ��C>�h�*�ͽv��=��_1���#���$��������"=�
�=Y7R�"���
� ��b�x�F���.?}y$>��ʾ��M�#�-<�oʾ����1ք��祽�-̾��1�#!n��͟?��A?������V����.^�����ޮW?�R�!���笾
��=묱�О=� �>�|�=!�� 3��|S�+r0?J_?q��T���*>�&��0=ܽ+?��?��_<kH�>�;%?4�*��N��0[>��3>�ȣ>���>�g	>5���۽��?�qT?����뜾��>@w��ƴz�طb=>�c5�Ϥ�+�[>}D�<M����V����,�<?W?b��>��)�$���[����9�:=`�x?�?�e�>݉k?I�B?��<�a����S����w=o�W?"+i?Ϲ>.����ϾP���%�5?F�e?�O>M�h�	�龈�.�&U��?�n?%k?g8���}}����g��)k6?�g?��]�HC����(�Hw]����>��?��?+eT����>)�>MJ'���a��h��I�?��	@��?u������V�S=�1?,�>zH;RC�Z[<Hɾ��i>��>�����Q��.�!�������S?2��?�?9J����
����=O����?U?�?Ž���Q�=L����ga����
%��7e>v�����<y����O�z��辀듾W�E��pk>��@dg�QW?PM��k�ￅ�ؿ��v��A���{��-�>�9>hqk����qG_�`�b��4�D6��a��M�>�>.������,�{��q;�V)��k�>(��	�>L�S��&��횟�K�5<|�>��>E��>�*���罾!ř?]c���?οS���ӝ�<�X?h�?�n�?"q?כ9<��v�T�{���V.G?��s?4Z?�o%�,=]���7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�ط>���?b��=f1�>�)�=Ѱ�QX���y>F�=4�s�s��>��I?�G�>x��=�}*�z�/���F�T�R�)�rMA��>�]b?|�K?��]>Ԥ�������!���ԽY~*�L�L�m@�V]7�р˽�M<>`�>>�M>�2M��׾Y�?���u�ۿxZ����=�LH?^ט>f.?�� �2|t��]C��?��>5� �OQ��"=��fO��_�?�_�?op?��ܾS����<��>�X>$?��/��+þo�>�O�>&X^�{ĥ�Nt��H �>�H�?��@�Բ?�����?�*	�$���ք�yվ�v ��T>�=?B��:o�>b�>!�+>��}�ʔ���Yq��I�>� �?�}�?*��>�a?��h�LA'���=̚�>H�R?��?�1�ɝ쾏mS>��?�p"�����u��Vm?�.
@|@��_?�E��o��u����׾�s��9�(>"M@>�ɐ>b�i=�ƃ>������ؗμh >���>Bc�>��>�No>X0 >h�>*�gf�����%���;��U�DF�B ��~������SH8�v=��~:߾H[���+��̼)�oEx�2B��ּF�]>�XQ?�bV?��?d?�E��>�"����=D����˽<�>��-?��,?,�-?�=Fܵ�r�ջw��Έ�զ��;��>*ʂ>��~>.��>3R�>�Yr���>�	h>���>��]>1��=F"��j�X�r>H��>�B�>�q�>�C<>��>Fϴ��1��k�h��
w�q̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��v�T�4:>9����j�5`>�+ �~l���)��%Q>wl?Nif>�u>��3��V8��P��y����|>�36?���R�9�Z�u�n�H�Nrݾb�L>�>�SD�fU�\���bi�+�z=�~:?�x?m~���밾^�u�	���R>�A\>�v=\�=NHM>��b�	8ƽH�G�=T/=�d�=��^>�@?��->�̐=�o�>�%��bXS�`�>�A>��->�@?��%?`��ܪ�����Ԏ/��lu>EQ�> {�>c�>NiI�xe�=q �>��^>�`�G ������B���V>Xg��`�򏀽���=@���e��=��=�� �
�:�ޕ*=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾHb�>�j�1ȉ��fY�X��=���>?�i?rOؾm �����)�@?3$?Dg�$��� п|~�����>WA�?��?*"Y��f��\�B��?'�?��V?�U�>'� �X����!8>�#N?W�P?F܁>�t��O�v2?Ri�?�Z�?��g>F��?�_?� �>e~��PF�ض��=�n���3>�I@>�J�>C����Ǿ9=2�m���i�҂I�VkѾ��>�S_=�8�>4S�ύ���!>	,����q������>Y��>Ʒ(>��&>ߧ�>���>���>�	۽�E����(���T?_��?�l��i�K��h>yx�=�_��T�>�WV?%�=R��(�:>6�i?��?6}?I�>X6�RY���G���ޢ��3;�C>�n�>X�?��p=$�q>�´��1f�<�[>Q��>��;�Ⱦ��ʾFؽ���>}I?;t�>�1�=��?�#?M_m>F1�>�fD��]��r�H�(S�>M:�>0�?�U?~�?����S3�)�4A��UZ��ZN>�Ex?�h?�5�>&���(r��k�ٻ"S�/����?��g?�ǽ�?�և?�O=?��A?Dj>��׾O(���<�>��!?���A�gJ&�>��+|?4I?{��>���ս�-׼����n��<?/\?B&?X��8-a��þ�1�<� #���U��p�;(C���>�>�k��
��=c>D�=HNm��I6��4e<�\�=�~�>>�=[7�z���� ?��׽����� ��~�O[�Ͼ�>��m>�_׾��f?�����r� "��v���ɻ���?b��?[��?�a$��Ga��-?yZ�?�w?!�>�ߋ������>�:V���������k>���>+G������,��喿[��OJ�Ue�>6�>E�?��
?EX>wt�>j���6k3�5a�В�l�T�Y����<��C*�N���~����,�����3��Qfa����>��A��e�>�;�>?c>��>���>��<�Sl�>W>G{}>���>�7n>g�'>�Z>"�=Պ��3KR?�����'�5������3B?�qd?�3�> i�7���[���?���?<s�?�7v>�h�l-+��n?�B�>���p
?�P:=�l��b�<�T�����5���)����>pS׽�:�JM��tf�j
?�/?����̾17׽>ȕ��B�=広?/?�o/���S��4s��Q�ѠH�o#���9������/ �rGp�2J����w��T{�y�!�<�Y=^�#?$C�?��M�쾥����q��/X��>��?W�>�U�>2/>���# �xCN��#��9���5�>��{?0�>�sJ?}#9?�LP?�KS?�<�>j��>����*��>ՙ@<I�>/��>��>?0?i"1?y�?�\'?��E>���'��5�پ��?�?��?���>��?�Z�����.���`���V��	a=���:�ݽ"�N�\3x=��^>�X?&����8�h����k>F�7?��>F��>����,����<'�>��
?�F�>E �~r��b��V�>���?�����=��)>���=������ҺnZ�=������=�5��'{;�B]<ق�=���=�<t�^べM2�:蝇;�m�< ��>�;?1��>�~�>Q����(����к�=Nc>�1X>(36>$�ؾ�q��骖�� h��Ay>/2�?���?H��=u��=�=<%���Ⱦ�%�����Y�<7�?#?�5[?�r�?�58?T3!? ]>���^��!���Q���k?w!,?��>�����ʾ��։3�۝?i[?�<a����;)�ߐ¾��Խұ>�[/�i/~����>D��텻���V��6��?�?MA�W�6��x�ۿ���[��{�C?"�>Y�>��>U�)�~�g�s%��1;>���>lR?�L�>��O?�E{?��[?.S>�8����ؙ�/�$��">j�??Xy�?�Ў?h�x?c�>�>�*��p� ���^����D#��O�P=j9Y>;�>+��>q1�>�}�=Bƽŀ���>�R��=F�d>���>�4�>�s�>�Bw>�<��G?��>�[��&���뤾GɃ�I3=���u?E��?7�+?Xq=��Y�E��G���G�>�n�?���?4*?޷S�%��=�ּ�඾y�q��#�>4ٹ>.2�>N��=ņF=�n>�>T��>%��^��o8��dM���?F?	��=��ſ�[q��p������Ey<.�����b�'ߓ�q}\�p �=z4��������D�\��������p���E����|�7`�>�=��=[W�=b��<��ͼ��<ZVP=�ǔ<J�= zn�2g]<��7� (λ���������e<;NL=��оXm?�9?i�$?�I?�y>�q>QA�H�/>l\���?��4>�8����;�<<�|�������߾�`羃�k�q|��?�>�z�x��=F>Ɲ >]^X=��>�}<F�=I8� �Z=H�=�}�=��=c��=�>y��=� w?Q���6���JQ��+罊P:?���>,�=��ƾ�$@?|�=>�"������v�&?���?�y�?06?v�i�X�>1â�?v��!9�=����G�0>W��=��3��>3K>>�tD��������?�k@N�??�ǋ���Ͽ76/>�3>i�>�>R���0��X�la�q�S��Z!?��;�E�;T��>=��߾I�ǾG�(=��4>�e=����Q\�8��=�ky�B�@=w�m=�k�><wA>�l�=*צ��ͻ=wYB=���=GL>���B6� �!��F5=h�=�id>_&>y/�>B�?td0?dd?>
�p�� Ѿ�����W�>1��=�>�`�=�{@>e��>^�6?7hD?FDK?7�>a��=<��>3��>��,��m��i�5���2x<��?�?�^�>��f<�*A����:d=�����L�?b�0?D�?x��>�U����:Y&���.����P4��+=�mr��QU�l���Pm�3�㽱�=�p�>���>��>9Ty>�9>��N>|�>��>f6�<pp�=�ጻ���<� �����=#���|�<�vż񖉺�v&�A�+�e���X�;���;�]<���;��i=��>�8>ҕ�>��[=������>$T|�[[��9�=�;���:/�3Fm�Vy��U%��r��' g>��F>꽱䎿�S?�� >[nd>���?�ʀ?��]>�L
�S��J����Ƚ{j��5E>��=����>�]�8�y�*�p��g;d��>�ߎ>;�>��l>�,�Q#?�6�w=��1b5���>�|��r��)��9q�@������^i��JҺ�D?�F����=W"~?�I?S�?э�>V���ؾ ;0>�H���=r�P*q�fh����?�'?җ�>�쾐�D�#@̾Q뾽��>UI���O�����Q�0�P���÷��v�>!⪾u�о#3��f�������B��Ar�o�>y�O?M�?zb�U��pUO����i���X?*�g?K5�>�L?�??+��+��_����=0�n?��?�9�?#>���=n�e�>) 	?���?۫�?�s?�=?�p1�>y;R� >7����=�_>�Z�=M��=ep?O�
?+�
?^m����	�j����D�^���<r��=���>7��>�r>~ �=OFf=�l�=�,\>�>��>�e>L%�>U�>�?þإ!�Y%#?Q��~ӿ�9n6?���>�Z>
��~�#�bb>v:{�pTx��뀾SϽߠ�==1#>�U>C����>J]ʿ��?���<�6��`G?G�ZV�[O`>���> �=D�?1��>*�G>=7>a7�>�=�Г>�O>��G$>B'�T4'��iE���D��eǾ�7�>�J�㕡�
n��	���o*��l�f(�������:a3�_�>"Z�?0�ƻG�l�C0�V=���	?�h�>�L?O����� �)C�>r�?l�>����"���r��F� ��\�?��?�}b>[>�>|�W?��?�8�s:�ɂ[��It�x?�+e���]�ub��w����.�b�Խ�^?�w?��??���<sgy>)ۀ?m?&��E����>\90�]�>��'k=��>���u]�Z�ҾE�Ǿ���;�H>N>m?��?��?K#M�AQ(��t3>I�8?��2?"x?:"3?^�7?�A&�b&?��1>m�?��?�t9?l?0?��?.�9>���=1��W��<
떽����Ľjg����|�)=S��=���<��k�
=Z6�<� l����R�:�y�i�x<$LI=��=���=Dצ>V�]?P6�>I��>�q7?4��D�8�����A8/?r�C=����(R���٢����6�>��j?���?J)Z?+ce>�LA�a�A���>R?�>�m&>�!\>(ұ>'��E���=��>��>P�=%fE�-���
��j��AF�<T�>��>j5|>}��E�'>uv��$*z��d>��Q�;ź� �S�1�G���1��zv��\�>��K?��?��=:a�X@���Gf��.)?�\<?�NM?��?��=��۾U�9��J�C���>�x�<k�������#����:�V��:i�s>$0��>砾�kb>���2c޾�n�eJ���羦�M=Ih�nU=�2�B�վ+��\�=�A
>Z���N� �q��{Ӫ��9J?��k==w���oU�MZ��r�>���>��>�:�4�v�qs@�����=��>��:>�L��P���{G�2.�'�>1�W?߄R?ߍx?�E���p�5B�G�5�(�4�V`>'L�>ݯR=�(%?<�>���=��
���&��d\�Y�O����>Q��>���+o�F��ܙ��%�T�;}9��,?�5�>l�!?��>L�*?j�?�G?l�>ߧ>���s��ql&??N�=�ӽ�Q��g8���F����>�H*?'�>��u�>7�?I�?�M(?�R?�?�c>N��;@�J�>p�>ҮW��'��U�]>��J?�	�>k�X?|W�?a�>>�z5����������=�V$>/�3?[�#?��?mŸ>�@�>Z窾�R�=`M�>4�]?�}�?ũs?g�=	�?+�7>���>�[�= ѫ>���>?A?~�O?v�n?�E?���>�n]<�έ������<��,ּ�:h��GA<m�j=9���H�Ȗƻ�%�<�l\<|4��mሼ_�ż������/��<)^�>|�s>o����0>C�ľ-P���@>����N��ي���:�xݷ=���>��? ��>�S#�ᾒ=���>�J�>����7(?��??��";��b���ھr�K��>�
B?k��=y�l�3�����u��h=��m?Ή^?��W�$����b?K^?#F�i=�E�þ��b�R����O?z�
?w�G���>�~?V�q?��>(�e�N;n�/���Eb�k��ζ=Xl�>4V�*�d��2�>�7?w)�>h�b>{��=jj۾2�w�4q���?���?x	�?q��?�*>D�n��"��e��Ϛ�pd?�&�>�ؾ�7?��:�Ѿ���)��3���Ե���c�������t���dO���D������� >�?�Yu?��_?L�^?��㾧�m�Te�U����F��0�s���C�ܻN��
H�s/w���)z�#"���@�<
ln�n�Q�R�?A@&?W�v�!�?H�����ؾt>�r�P�����=Slp���<���=��=�Jb�!.����?�¬>���>��A?��R�ey=��D8�N�A�����3H>tӏ>���>o=�>�ɔ��H@�<;��ү��?��I�ƽ��w>�v\?��G?2gu?eo�GS��c�=���<RO��`�|=��]�3R�>��������/���H���g�Z�̾d�������v=֊&?/k�><"&>c��?�@?��쾦|��A�ľ2	�&��<���>��g?�t�>��=����^:�uǮ>�>f?r� ?��>Ҙ־������;�k�>��$?#��>�ڂ�ə���+S��wx�Nq����_�=��g?�{��6̽@�>�_T?�?���|����>3�M�����s�Ww@�А��BO.?Y�=?�`>�������qY�j�h�0U)?��?<�k�.��a{>��?���>�&>d�?>�>o4���
�P?bn?ԝZ?�lG?K�>&���k;	���A�u9�=V��>v;H>(g=2��=,D3���;�.t&��A=�=�����7�rCx��c<���<�s=6��=6�鿹�d��F�&I�G���G���j�7p����ĩ��3�"�� ��M��>v��ϽN=!����줾�@�� m��1�?q��?�ξ5-���͡�+i	��	^�>g��;4!�s�Ǿ՟��]���`���{���$��SZ�B�a��Ow��M'?�O����ǿb����[ܾ��?��?��y?���U�"�W�8���!>eF�<n����뾙�����οԚ�I�^?�%�>r�đ�����>�@�>�qZ>i�q>p�����:#�<Gs?�-?>��>��q���ɿ���S��<N��?@tUA?�T)������W=0��>
?��?>�21��d��1�����>*�?��?�N=��W�ȥ��}e?�<%uF�l�ݻP1�=�Ϧ=�n=���4�I>]s�>h0�)A�8�ڽ1�3>�u�>�M%��l�^�v
�<O]>x�׽9���5Մ?+{\��f���/��T��U>��T?�*�>U:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=l6�򉤻{���&V�|��=Z��>b�>,������O��I��T��=�:��Eӿ4p+��!���x=���<�%��QIֽ!��C���;�ǳY��r���P>��%>F:;>	<>>]�!>���>�Ll?=d?�y>���=#�I����������J
>�駽
͛��ؾ�N�_G��)�Ҿ��D�%�L�������O��ƃ=v�g��*����F���x�y5?��L%?\�>���������=�[ľLq��#u�=�b1�dl���;��~�ϒ�?��g?.���ۚR�������@�C��N?oS �&�־M�^�O�=��#�=ϯ;?�j>�=&׾{WI��YF��/?g�?a���+_����">`h�.�<C�)?��?�t�<dЫ>$�"?�5������Q>��2>��>��>�>�Z��b8ӽ�c?�P?����u���Ս>�jžL�p����=� >�CL�����.^>�i�<����#s��������<�"W?.��>��)�?�"h��GN�օ<=4�x?�?P3�>�wk?��B?T��<�n����S�z���w=��W?+i?ߩ>br���о���&�5?ϛe?�N>��h���g�.��T�?�n?^?<I��%{}�N�����*j6?,�s?Y�N��<��fF���= ?�>K��>:?�{[���;>I�7?���=\��e���L�7����?�W@@��ٽ�`�ݩ�=��H?��>e��9H�����3��`����?Zzƾ�h���3���̽�?�]z?�'?�þgH�����=���G�?�?	�羒б=)u�%o��t�1<6��%!>�0ʺ�r��A��o]I�����y�оʐ�?=SM;>�@n�p��ˣ>Ә�n�濳�ϿW{z�a���Fz����>�ą>3;����ؾ"�q��fs�Mf6���>��ە��H�>��>����s�����{�yo;�H'��>
�>?�����>ЛS����󯟾
�2<(ǒ>?��>|��>����Ƚ�U��?lP��0=ο��������X?\�?�i�?S�?^@<��v���{��S�)G?:�s?�Z?��%�h$]��n7� �j?�_��qU`��4�tHE��U>�"3?�B�>I�-�Ѳ|=�>��>�f>�#/�v�Ŀ�ٶ�3���W��?��?�o���>o��?ls+?�i�8���[����*�C�+��<A?�2>+���D�!�;0=�FҒ���
?M~0?{�a.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?B�>	�?C��=M��>7T�=�᱾[�3��#>�%�=�?�s?E�L?��>-��=I�8�c/���F��:R����O�C�>Ӈ>�a?�@L?�c>�
����2�!�L
Ͻ	�1�ab켴�?�Y,�T�ݽ�5>�=>N�>~�D�ZHӾ�[?�z����������� tY?��@>�z?x6�(r��<�;ڼ�?��5>�E�簿x���N�ڲ?��@�?چ�����ͼ���>���>1�|��핽a��(ZN>��.?`��P��𷅿�ȩ>RS�?;�@V��?�W��Ӹ?�"��'�����8ͧ���/�V��=��L?�`���.>�� ?e1�>������?1q�=��>=ܲ?�e�?�0�>p�Z?�rg�2���X��<�>{�1?�?���=?��v�>�
?�9�xo��xLܾHi\?P�	@G�@F�_?<����hֿ����dN��N���.��=���=Ć2>�ٽ3_�=��7=��8�w=����={�>��d>&q>0(O>sa;>��)>���M�!�
r��X���Q�C�������Z�7��0Xv�_z��3�������?���3ýy���Q�2&��>`��8[>��S?��<?�Q?.�?�[=S=�?��~g>�%=ʎH=�C�=%�<?�^]?
�A?xW>����3=c�gRy�낻�0}����>t�>�M�>��>Oϓ>�G='>{�o<��n>���>g�8=������H>qh�>֯�>/>r>m�0>&�>3���᯿mhk�񊅾L�޽C�?3Ɠ���M�;՗�32��;5����=�d.?���=Bd����Ͽl�����J?����M]�z�6���>{�/?;�T?[,>�V��(�U;6>�'�<�j�ߪ	>z3��&y��%���W>��?��f>P'u>I�3��Y8���P�V���U^|>�16?�඾�;9�+�u�X�H��[ݾS1M>���>~�E�fo�����M��yi���{=v:?��?���~ް�d�u�a;��0>R>+\>P�=|g�=�KM>�Ac���ƽ�H��1.=���=p�^>�8?��/>n�=K�>�6���&\��>d�;>��<>��@?�v#?Fy+��-ý����R$9�M�r>Tc�>��>٣>�IN�j|�=k��>�AO>K��Ԃ�ߌ�_�X�Ib>�,����f���Խu=뿁�P>Y�#=�M�&t4�G�&=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ˧�>���ƙ��J@��+aa�ڈ�<�O�>O�[?�PǾ���Z����+?Cu�># Ⱦg���Կ>x��r�>;<�?]*�?��c�����L�^��}?t�?�U?�q>���_sٽ�A�>��M?�}H?�1d>�.O��'��K?k��?͔�?ѠP>��?8%q?�`�>]�t�3�=��꧿M���gj=��ٻ�.>��*="e��ۆ?�<����Y��P�m�%N�Bm0>T�<qI�>\������U��=R���=J���%A��ٛ>a<|>��K>xp�>W�?��>�:�>p-	=�`ݼj[k�SΩ�ބJ?�<�?���p8V��Σ=I��="�zΓ>��@?�u>�3Ǿ�L1>,g?�G�?R<o?1D�>�4��z��}#���Wž�rj����=v��>3��>|����>���ҷf��Ś>>�]>�>�;�Z꾷O����>;�|�>� ,?���>�2�=ˎ ?a�#?1�j>q�>�`E��3��O�E����>I��>�1?��~?��?O���^`3�K���ϡ��t[�7N>��x?BC?&ҕ>W���Y���&�C�K�I�툓����?g?m��t�?��?No??P�A?&�f>D���ؾ�d��d�>.�!?��ĂA�}'&�Ƿ��{?b?&�>�,����ҽ*�׼������4?G\?�S&?���B8a�f�¾B��<
�(��I�	�<BD�D�>�>�򆽐j�=�>���=� m�g�6�g�Y<v�=.��>��=��6��ڎ�aq&?�W��Bʔ�M�T���\��L��u>��>.���Y?i����=�2���pꜿd����?^�?四?e,��)��{�0?o�?��*?�a>g]ξ~8������p�����cӾSb����>,�����֛�,��9ё����}�M��� ?��>��>�4?.��=���>p�*�AkD�N��[�߾Օ`�D%��"R��>��o��"�b�M"��Ⱦ��z�Z��>J)m����=k�?̙�>�r#>��>�R�=d�u>hY�>i��>���>�>��>U�&>:�����;�KR?����!�'���达���g3B?�qd?P1�>Pi�:��������?���?Ts�?'=v>h��,+�~n?�>�>H��Uq
?bT:=9��:�<V��p��3���3��>�D׽� :��M�=nf�vj
?�/?�����̾�;׽N����k=�5�?G�(?�G*�{)Q��o�x�W��S���"��f�&\���%�d�p�E!������a��^#(��-=��)?��?;��]�(��F�k��@�?�h>���> �>��>��H>��
�Y�1�Vr]�}�&� ���G��>9~z?I�>P7;?��9?agQ?u�M?GU�>|�y>�ʾ{?}@�<"��>
}�>3	H?��'?��8?"�!?�,?�9>р��7�X��G� ?�� ?��?4��>z�?���Gٯ��C�����~8���5z�̈́W���>�Xƃ�^l=�"Q>�X?	����8������k>�7?��>~��>���-�����<��>
�
?�F�>% �.~r�c�JV�>���?T���=��)>���=뉅���Һ�Y�=������=S8��{;��f<��=���=HAt��ہ��!�:$��;!k�<�d�>!U?��>Ypg>�g�����2
$�`Z�=��u>��">b�?>0L���ҋ�E��Pvk�/��>DD�?:�?w(>	�=��>v�ɾ��!"�_輾�GX����>Q�C?Bnz?�}�?`�?��?v�>#;ƾ����H�� ����^?n!,?��>����ʾ���3�ĝ?`[?z<a�׸��;)���¾�Խ��>�[/�i/~����6D��腻���2��-��?⿝?�A�I�6��x�տ���[��u�C?�!�>�X�>|�>C�)�c�g�y%��1;>��>WR?�e�>�d?�l?�KE?Q��>D]-�����X��H�>ʹb>g)3?��>?�x�?�a�?�-�>ۣ�=�ŗ���ɡ�.yw�I
�������w���$>��>���>٘�>�|�=î�������	�܎S=��>��?}�>���>s4>yev=��G?���>�O���������΃�uF>�!�u?���?��+?��=
w��E��S���$�>�j�?:��?�-*?�xS���=�Gּ�ﶾ�r� �>�ʹ>��>���=��G=��>���>\d�>_+�5S��U8�{DN��?�F?4��=n ƿ͢q���p�����gd<P��3e�����{�Z����=*Ř�m��-Ʃ���[��������k ������.�{�>��>(x�=
��=��=��<iKɼ�½<$�J=���<"�=�Rp��Ym<��8��]λ򛈽�j�=\<D�I=.����)����{? J?E0?V�<?vh?>��	>i�� ْ>`P��5�?;t/>M�;�9R¾Hd1�8�������<ݾ�BϾ��c�癜�g4>��8�؇!>��:>��=^�ʼ���=�7=�~�=n��;�Y*=�r�=)Q�=�y�=]P�=��><��=�6w?W�������4Q�Z罣�:?�8�>{�=��ƾo@?��>>�2������zb��-?���?�T�?A�?Cti��d�>J��i㎽�q�=i����=2>f��=~�2�T��>��J>���K��<����4�?��@��??�ዿТϿ5a/>�4>\�>�FR��X1�<aX���a�RsW�͇!?v*<�jB;�
�>q�=V��B�ȾJ�=�3>��o=F���\��G�=vc|�� ?=��j=���>��F>g~�=M�����=a$R=���=P>���93�3�+�/�n�>=���=Z�`>�-(>���>�N?�'/?X�_?a'�>yPu��پb��	8�>vأ=��>�ޙ=_#>� �>Ʀ,?y�E?8K?z�>8d�=�Y�>��>z�2��mr��d۾�ɬ���߻�M�?�"�?,w�>"/<*I��Z�=:�#F��dM?+�)?�?��>5���	�'�,�%�.;�J�&��ڽ�������0�Մ���O�&����,>^�>bW�>c	�>ثU>��>=�V>��>�{�=|���sͬ=����2X=�#���=)�=�^�C��ٷ<�x$�H+`��(��kK[���Z����2}=qoH=&9�>��=x�V>HW
>�X龂iP>�w:�܏z���^�.3/�d,�������k?��{)�V��>�;�>YKS�]����I ?��$>�8�>%��?
k?�>�3*�ƙ׾�{��e�e���:t�=;��=LVI��_��j���P��վ���>��>��>�l>�,��2?�/v=���U75��,�>Ӆ�����M�L4q�>0����i�IP�3�D?�;��а�=}~?Y�I?�׏?qr�>�����ؾ&�/>����I=���q�����?z�&?�U�>D��K�D��A̾� ��f�>�6I���O�߿����0�!�t˷��}�>>쪾��о(3��g������J�B��0r�R�>J�O?��?Xb�Z��w\O�����\���c?�g?�6�>-M?;?�0������p����=��n?���?�8�?q>|@�=�fǽI��>1Z
?���?�t�?�t?� 8����>��;{,>������=�5>`��=g��=QC?A�?��	?����w	�II�)n���m���<��=\ߎ>� �>v�w>O��=�k=IM�=f�d>K-�>�<�>�g>9�>Ɗ>$ʥ���d]?a;:=p���T�K?ru�>�u�=`���!'�S�h>�j�������)�����,m>C�>>�]>W�y=�	�>�%ٿ��?��>�B1� �:?���C�꽘vr>rX�=Rq�=vl?���>ZZ?���>U ?��(="H�>��>��ݾV�D>�'��@"���P���g�ZQ����>�'�o�����!�C��R�h���z�ϻq�:ބ�O�G�X�Q�"��?Gݽ,�_�k\9�s�	=eZ?���>��B?:����g�<�k�>	�?Q�>����� ڒ�F⭾ߕ�?P' @�U>8̔>a6U?�e?,�h�i�;���\��Mr���=���e�bMH��<��������^J�a�Z?�s?f�3?�DA=�\>���?Z:��ZǾP��>��;��L���>�'�>#����o��ľb��D�6��_U>��^?�]n?��?w1���>s�!��.E? �e?�uc?38?9 �?"e�=WM�>+�>Ù?���>�pJ?	kM?�>N?)�o>��!=�X?��T���*՛������+=[p�=�Dl='�ؼ��#=�Z�=7�<8
y=.�=IƼ��ͽ�fG��#m��[}=3�>��>�Q�>G"]?\��>�v�>m^6?6��9R9�C����j/?�H=�G��d3������9��c�=�-j?)t�?��Y?�g>ԃB��@���>�U�>>�%>E[>�>S��B�A�j��=#>�~>�h�=E�Ԛ~���
�*�����<�>���>T:|>�č���'>'`��Yz��}d>R������S���G�>�1��;v��]�>r�K?��?���=�`龓����Jf��)?r`<?�PM?��?
�=̹۾��9��J�XG���>��<���¾�������:�)�:x�s>�&������¤b>E~���ݾ�\n�aJ�u��I�L=|��"T=�/���վ��~�I�=�|
>����� �����Ī�J?��j=JG��B-U��3����>45�>}خ>n77�]x���@���$�=���>\Q;>�И�6����G�� ��#�>%2L?ƴX?� �?PI�Yz�O����Ľ]ym�M�=���>j?�>��G>��꾌�*�g�v��)�}��>8��>��6�/pS����_��BT�?;h�@�3?���>���>�D?�~(?��X?5D?��?N=>��L�����3(?���?e��=�н�)O��#;�3uO�n��>�N/?��$�?J�>Q7?�O&?&�+?SU?i�?���=Ze��>C����>�p�>p?V�!诿�to>G�H?��>HjM??8�?m�r>��0�a˼�a����7>�iY>�0?%N?1F?MM�>:��>����Zt�=_��>�3^?o�?aw?��>�j?��G>�%�>���=���>�(�>-Y?�O?�Vo?��E?e��>���<�w����½�����뼁���3<L�=���"�3��}�|6=��<�hX���_Wm�[�q���@�<AZ�>
�s>l�K1>O�ľwR��!�@>a���^��V銾t:�V�=z�>��?���>C#��Œ=2��>Y9�>����;(?��? 	?|2;�b��۾�K�h�>��A?ey�=��l�΅��6�u�7�h=o�m?c�^?Y�W��!��y�b?��d?��澣84�.����߄�����9?��?*�.��̩>�6q?Vjz?H?{�/���e�����5g��G���6�=:��>(�5)k�2��>L�3?Ù�>e�G>}Y�=�ܩ��Bm�t����z?V?<��?FO�?.l>%�c�"dۿyZ��ᒿl-`?���>dȲ�:�&?�w�S�;f���f͎�uھ�Z���~��E7��E�����a���tGؽ�	�=�F?�Gr?Ro?�_?����J�a��N[�^����Y�?:�h"���B�$�B���B���q�;�����Bߞ��_=��f��O�Q�?:+?�<���?��Jݾ���d?(>YLo�˯�+�="�/�9?�����=�?�-�'�����.I?��>���>Y�@?0�I��)��Y"�V{L����d!>�G�>4i�>���>���;�����ὭվDέ������y>��\?z�J?���?L��N9?�N�Z6�Ŋ,�q�ľp�^>�K>���>ssP�^_��t@��QM���`���Ҿ��������=�?+�w> u?>�!�?��>!J�������O����=o�>�:s?� �>�I>����4�;1�>�Yb?Ӗ?�>�V�1��Ƃ�@�z�� Y>z�>�7�>� s>_�/[������q�Q'��Ի�p?�QY��]9�+�>N�?���=�ѵ<�n�>�Z�=�����;�m�C��9K=+Z#?�
�>/r>���+�6��Xa��ٽ4'$?�B?߳C�GF����=�?�<�>�!F=�ޑ?'?Z�ž���e%?qȅ?�Tx?��?p��>h����g-�{�R�n�*�R>7��>�nx>,�&;��T>�q=�#�gs�����K5 >qy�������ӽO����=�����e>��ӿ.<N�3u�����h�Y����p�ۂ1�o}��o��c[��0���߽�2�Q���w��ƌ�А	�Hs�?"7�?��Ҿ[����ő�%y��$n'��Ǉ>(�P���VdI����=^t��U��U߾؇J�1#i�eZ���`�׎'?������ǿ㭡�>@ܾ ?�2 ?רy?�	���"��8��� >'��<������ў��_�οۢ��k�^?)��>���E�����>O��>��X>�:q>�釾H잾�<�?ʋ-?���>ׇr���ɿ����U�<��?�@|A?��(����V=3��>ђ	?"�?>�P1��H�@����V�>h;�?~��?�oM=��W�Ġ	��e?<�<��F�t�ݻ3�=�B�=�L=��a�J>�T�>̌�[A�^8ܽ��4>څ>�z"���c�^����<8�]>��սf/��Մ?\z\��f�@�/��T���T>6�T?�)�>*B�=O�,?V7H�~}Ͽ�\�Z+a?�0�?u��?��(?�ۿ�7ؚ>O�ܾ�M?�D6?���>d&���t����=�%�`o�����<'V����=n��>�>?�,������O��Q�����=~m�1�ɿe�&������<=�=�*�<'���ꌼ�)�\wݾ8��y��� �=u�>*�(>�zz>��J>q��>��\?M�n?��>�[,>{�)�>���O�Ҿ+����V��c���u��7<�Ծ����Y���*�������ʾ�B=��ψ=T�໎�
#��~i�!�E���,?�1>j�о�DQ�o=�<݊ξ�d�����������Ҿ��/�!i�S)�?n�I?g����S��e�sܔ������ZX?������������>e
�h��<E"�>� H=��q�.���P�P10?�y?�@��h���!�)>"� ���=m�+?N� ?��Q<�T�>��$?Lh,�� 轢$Z>��3>A<�>���>��>����4۽I�?�T?�?�c��b)�>7ľ��/y��Pc=��>��5�Bv�O?[>�e�<���� jS����� l�<�'W?>��>S�)����a����D<==��x?��?B1�>~{k?A�B?���<�j����S�F�Igw=b�W?0)i?ѹ>r���о�~��2�5?v�e?��N>8ch����.�.�pU�0"?B�n?`_?�g���w}�/��>���n6?P)u?:�-������)m���>�?�ۊ>.�@?��q�Z�=~w:?��>�7��<�����!���?6V@�g@�����
��w�=ro$?�$W>Nu��	�/M��_��54���>����,p����ɾǁ��9��>�Y?5��> �Ⱦ�{�}E>xذ�؂�?`�?�n�HV>�۾��j�:��u�G�~��>�Cռ�-d�m 侲�e��>U�]I̾+ ����C=>�j>�&@	��Fc�>�b�=k�⿂����P���Ƽ��(8�>��>�R�����<�e���W��j#���.������M�>��>���'����{��q;�a0����>���	�>��S��&��m���B�5<��>��>鷆>�,���罾ř?&c���?ο\������>�X?h�?�n�?q?�9<l�v���{���j.G?��s?FZ?�p%��=]���7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�[�_?#�a�G�p���-���ƽ�ۡ> �0�f\��L�����Xe����@y����?M^�?e�?ܵ�� #�b6%?�>e����8Ǿ��<���>�(�>*N>"H_���u>����:�i	>���?�~�?Ij?���������U>�}?���>N?�?!�>��?R��=X:����<�n>b�=@Յ����>��G?M��>o��=�&��l5���I�8>N�L��<����>@"_?��C?�Wd>�)��&[��������Ō8�ʨ����8�K�.�|߽�`>?�4>@�>@�Q�n�ھ��?�f �e�׿$���$l���'?j>�|3?_���r<�0���AЈ?=�*>����b����u�+D7�(��?	�@��?��о���vA=�Q�>�?�"�=!�dǾ�MC>��.?����W��|��E��>�)�?K�@v��?q����M?�����	��^&��a����Y"=��=?^U?����.L\>�?�`�>{�~�a���b����>et�?kp�?x��>�T^?�b��8��@;4��>��d?��
?0V������=l\'?�+�b癿����Wp?N�@��@H��?cZ��{㿵���(��+���6F>���=d��>�
� �߽�=2��������>؇�>�
I>,+I>z6�=t�=��>�������~��u,����7�^?�W� ��T�PN�����"�+���澲c־�\��B�J�H/����}��7�ۦ���>Y�5?ƛQ?��t?���>�o����D>���=�3.<:,Y��s>YE?hP?�~3?�0v��a¾1�j��5h�܇��Yw�����>=*�>�>ѽ�>I,�>ٻ��� ���5+>���>U>ֆS<V���ؽ���<�P�>�t�>�G�>�C<>��>Fϴ��1��l�h�*w��̽/�?q���U�J��1���9��ڦ���h�=Cb.?�{>���?пa����2H?���})���+���>x�0?�cW?L�>��M�T�d:>����j�7`>�+ ��l���)��%Q>zl?��f>�ju>�o3�N8��P��a��v|>}�5?�g���]8�3�u�I�H��!ݾ&�M>�>ػD�(T�o햿��~��|i�1Ez=l�:?��?ɕ��Tాe7u����%�R>(l[>t2=�d�=O<M>��e�d�ǽ��G���-=�=��^>�M?��?>q,�=}4�>q���"_����>�c'>��>��A?Ύ&?뢩�뾿�����'?�u|>�5�>�w>Z>�_B���=��>��U>�x,�Ԯ<�|'�-pI�$�Q>��ˏf�D���`�=$_�ai>d$>=d ��m:�I�E=�~?���!䈿��e���lD?N+?$ �=�F<��"�E ���H��C�?p�@m�?��	�ޢV�3�?�@�?(��#��=}�>׫>�ξ�L��?��Ž:Ǣ�є	�G)#�lS�?��?N�/�Zʋ�7l�j6>�^%?��Ӿ�ګ>�q��(����Ł�	e��ؽ�7>6d]?����^���T�ݽ�J1?���>q�Ѿ�Ҥ�{�Ͽ#2z��u�>h�?���?�[� ����dC��c?OR�?��P?��>9��L޸���M>n'E?�N?�>r>�D��@�=��?G�?�n�?��U>;.�?ko?���>)6�e:?��[��엃���;~�=�Ȫ>mSo>�־s[�
�����U���B�}�=�`>��c=l�>`������W`=HG��iͬ��ڽ���>���>��=P�U>�O�>k8�>9}�>����ɽ{��>���G?0�?z����S���E<���;���ޑ�=|\b?�ϟ>),پ���gfz?o�?cd�?i~>*$%��t��-&���y��V쵽-��=�L�>�O�>�)�=���>�Ц���&�>��>8͓>�_�)	�gR�×�=���>�)?^��>��>�� ?P�#?�]j>�>�_E��=��[�E����>I��>z<?��~?.?�۹�vT3�o��d顿��[�a.N>��x?�W?�Ǖ>싏�w���?jC�H�H�(��⠂?+hg?��-?�2�?�??�A?,�e>d{�)�׾�[����>7�!?N �g[A�g<&����PX?��?6�>3����˽��ּ�v�����f�?0�\?�&?I���a�\þ�@�<29�<��Bw<��N���>��>}ރ�A�=gJ>ɀ�=��m��~7���U<2O�=��>[��=L�6����92,?Н�<�ߣ��J����q�']9��\H>��>�v���AL?�M>=z j��W������қ�L"�?~��?Hٗ?��f�Hw<?v>�?�}@?\ѝ>�3׾�u��Y��^��Db��������=;�>8o���پ�����"��%��(�V�a[�l{
? !�>_K�>@�>� 7>A�>��u�Q�8�S����վ�P�Θ)�h�K��#(�h�
���7���Խ"��z>ľy�q���>����V|>��?p�>e�
>��>H�?=�E>��">{`�>��>z T>E�y>�>�bƺ�䣽�KR?�����'�k�辴���X3B?�qd?D1�>�i�:��������?���?Ns�?+=v>h��,+�xn?�>�>C��Rq
?�T:=�8��;�<V������2��}�"��>�E׽� :��M�@nf�{j
?�/?���ŋ̾�;׽桠���n="�?��(?��)��R�|�o��W���R�t��h�h�d
����$��}p��ݏ�e�����4�(��1*=�*?j3�?������鬾�Wk��E?�t�f>���>��>I�>ʓJ>_�	���1���]�eY'����:9�>�{?��>"�H?H�;?@P?�K?�n�>4N�>nv��)�>�as<��><!�>�(:?d�.?JD1?l�?��(?X.Y>?����7���Pپ)M?��?�?�?Խ?���7�ٽ�Ӽs�W���j���u��b={�w<"�޽��}�BK=̆R>�X?���ҫ8�q����k>Z�7?���>M��>���N-��.�<�>��
?aF�>�  �I~r�>c��U�>:��?����=��)>!��=?���>�Һy[�=���6�=�7��O�;�c<t��=t��=|�s������(�:���;MZ�<��>�l ?�:�>$Æ>;�w� ��l���}=��>>�(S>	�>>�*��R#��f"����i�C��>��?���?�y=(�=i�><c���۾�J��m��'ߊ<�� ?͕$?e�_?�&�?��;?�,?��=����񏿹(��U���
?o!,?��>p��l�ʾ��ǉ3�ŝ?8[?2<a�H���;)�+�¾��Խs�>�[/�I/~����ED�E󅻵�����(��?�?�A�F�6��x�ǿ��\��-�C?�!�>�Y�>�>i�)���g�i%�X1;>���>NR?U7�>פS?rv?��V?,Q>�g9�͖���1��\��<j1>�9?�y?S�?ȶz?��>m�>�QB�{��?- �s$��\����'��<��a>2�>��>�/�>s�=s9}�_s���~`�tâ=�#�>�>��>&��>� z>X<��G?���>j[�����:뤾�ƃ�	=�a�u?���?�+?�e=���z�E�'J���F�>3o�?L��?B3*?]�S����=��ּ�඾��q��$�>Gٹ>�0�>�Ɠ=ˉF=�i>��>���>A(��`��o8�QM�r�?�F?���=ƿE�q��p�4ʗ�M3e<v咾��d�ϊ����Z���=Bߘ������?�[�y���b���|W���Ց{���>���=��=8�=���<{vɼ��<x�J=��<U�=�sp��n<x<9��@л������!���\<0�I=E2���¾��z?��I?p�0?�@?aqR>��1> o� r�>ߙ��J?<�S>S��H���>0���������X׾&#Ծ� ^�����>��a��*>�<->���=Bb�<%��=�Q=-?�<�����=��=�p>�{�=�=O>+ �=�6w?���������8Q�C�Ҷ:?4�>#��=�ƾ�@?��>>1������ac�~)?B��?�U�?��?׀i�a�>0���Ŏ�셐=�󜽘/2>���=	�2����>��J>��}K���c��Z2�?��@�??~ዿ��Ͽ:_/>�!/>�e>�pO�� 1��N���Z�6y0��U?OA��(־b+�>�U�=����*׾@�<�+>-��=����]��:`=�\���=�	)=]V�>��O>a� >q��f��=�J=)o�=�C>��{;��t����x�i=���=&RT>�U%>C��>t�?� 2?>c?斯>അ��ھn6ɾ�b>���=�к>�<�=ܽ
>.Ɏ>Q�?@�I?I?V��>�lV=�X�>Rd�>�i)���t�ծ��m�������b�?L��?���>fv�<c�ٽVD(�4*D�	����?�&?j�?t��>�����z�$�?!��<w�>�h>�q���G=�Gr��qվ|d��S5>h�>4��>�Qw>��,>&^�=�R�>���>�>q�1�;��<̐��d�=��ؽ��7>�8>�F��5��[����S�{��{�=�h�\��=#x�=a��n�=F��>_ߑ=�b�>� =�ٺ���P>6--�#
b�'�<C-�Sr7���o�����`�0��B#����>�;�>O�+��0�	?;s>e�I>P��?��k?eY�>[4��W�о�렿�茶��.���=�\�<xrܽ�Q�޾R���W������>Z�>5�>��l>,��$?�x=�⾷b5��>(��ر���}6q��;��D���Ni��׺�D?�C�� ��=	 ~?��I?���?���>C���|ؾ�M0>�K���;=�
�%(q�kf��� ?Y'?ɕ�>����D�MG̾���޷>�=I���O�d�n�0�t���ͷ�č�>;���B�оl$3��g�������B�Kr���>��O?�?q5b��W���UO����.��,p?}g?��>,K?&@?~���{��t���|�=�n?���?�<�?.>��=^�����>y4
?VՕ?���?�v?��8�ʡ�>�45<�t$>�ך�S��=,�>�y�=���=�?�a	?q?���:	�j��9���!h���<�N�=漗>�Ջ>��z> V�=o2�=s��=��\>��>G�>hUh>��>�u�>䍕����Y�+?Fń=���s�-?(n�>4�=�̼�6���y�=8o��BU�#3Y��B\���4>��G>�>�Q�Q�>��ֿ�Ʊ?+��>�~:��7?'A�(K�t��>~9>�Q;�"�>b�?ڋ?F7>�z�>q���u�=��>�[ξ_/7>��&�(����I��n~�c����t�>�H/��T��IM��\&=y��T�����qP��&���j\-�}D=/��?�tɼ�^k�f. ��=�|�?77E>E�[?w���>��R�>g1?��>�9Ӿj���$��2Rݾ�?���?[a>�e�>Y'X?n�?9VX��<�[�T��-v��F��g��PE��h#|��2�xM�۔_?يr?]h2?��y�)un>iE�?�:(�����L��>�B���H�9��=�M�>�_����j�r\��L�����{�u8�>�l?Uy?��?��X���j=g$��V�D?6P?+??��3?�!�?���k?�|�>I�?���>�Z?�C?%-?`>��2=����3[�<�x?��o�d'��Q�Ԁ������=�=(�l>���=M"	>�y�=�p�=��=��=A�r<��&>��>�H�=/v2>4T�>$�]?�>��>o�3?t�+�y�9�"���3�*?� �=̦m��W���o�������T�=l*j?m��?�U?{�f>�;�*�=��?>��>>�`>F�>�t ��[A��ĸ=�R>�>0�=u*�T�t��%��������<��#>8 �>43�>b^9�)�E>Q@��E�����P>H���=3P� �޽֠U�H�;�Dk�{��>��U?S�?fg�<҂ �Y&��]Z��?�q=?nZ?��u?tk=����4�Tl[��q��^�>5 ?>�L�
��� q���V5������u5>]�������¤b>E~���ݾ�\n�aJ�u��I�L=|��"T=�/���վ��~�I�=�|
>����� �����Ī�J?��j=JG��B-U��3����>45�>}خ>n77�]x���@���$�=���>\Q;>�И�6����G�� ��#�>%2L?ƴX?� �?PI�Yz�O����Ľ]ym�M�=���>j?�>��G>��꾌�*�g�v��)�}��>8��>��6�/pS����_��BT�?;h�@�3?���>���>�D?�~(?��X?5D?��?N=>��L�����3(?���?e��=�н�)O��#;�3uO�n��>�N/?��$�?J�>Q7?�O&?&�+?SU?i�?���=Ze��>C����>�p�>p?V�!诿�to>G�H?��>HjM??8�?m�r>��0�a˼�a����7>�iY>�0?%N?1F?MM�>:��>����Zt�=_��>�3^?o�?aw?��>�j?��G>�%�>���=���>�(�>-Y?�O?�Vo?��E?e��>���<�w����½�����뼁���3<L�=���"�3��}�|6=��<�hX���_Wm�[�q���@�<AZ�>
�s>l�K1>O�ľwR��!�@>a���^��V銾t:�V�=z�>��?���>C#��Œ=2��>Y9�>����;(?��? 	?|2;�b��۾�K�h�>��A?ey�=��l�΅��6�u�7�h=o�m?c�^?Y�W��!��y�b?��d?��澣84�.����߄�����9?��?*�.��̩>�6q?Vjz?H?{�/���e�����5g��G���6�=:��>(�5)k�2��>L�3?Ù�>e�G>}Y�=�ܩ��Bm�t����z?V?<��?FO�?.l>%�c�"dۿyZ��ᒿl-`?���>dȲ�:�&?�w�S�;f���f͎�uھ�Z���~��E7��E�����a���tGؽ�	�=�F?�Gr?Ro?�_?����J�a��N[�^����Y�?:�h"���B�$�B���B���q�;�����Bߞ��_=��f��O�Q�?:+?�<���?��Jݾ���d?(>YLo�˯�+�="�/�9?�����=�?�-�'�����.I?��>���>Y�@?0�I��)��Y"�V{L����d!>�G�>4i�>���>���;�����ὭվDέ������y>��\?z�J?���?L��N9?�N�Z6�Ŋ,�q�ľp�^>�K>���>ssP�^_��t@��QM���`���Ҿ��������=�?+�w> u?>�!�?��>!J�������O����=o�>�:s?� �>�I>����4�;1�>�Yb?Ӗ?�>�V�1��Ƃ�@�z�� Y>z�>�7�>� s>_�/[������q�Q'��Ի�p?�QY��]9�+�>N�?���=�ѵ<�n�>�Z�=�����;�m�C��9K=+Z#?�
�>/r>���+�6��Xa��ٽ4'$?�B?߳C�GF����=�?�<�>�!F=�ޑ?'?Z�ž���e%?qȅ?�Tx?��?p��>h����g-�{�R�n�*�R>7��>�nx>,�&;��T>�q=�#�gs�����K5 >qy�������ӽO����=�����e>��ӿ.<N�3u�����h�Y����p�ۂ1�o}��o��c[��0���߽�2�Q���w��ƌ�А	�Hs�?"7�?��Ҿ[����ő�%y��$n'��Ǉ>(�P���VdI����=^t��U��U߾؇J�1#i�eZ���`�׎'?������ǿ㭡�>@ܾ ?�2 ?רy?�	���"��8��� >'��<������ў��_�οۢ��k�^?)��>���E�����>O��>��X>�:q>�釾H잾�<�?ʋ-?���>ׇr���ɿ����U�<��?�@|A?��(����V=3��>ђ	?"�?>�P1��H�@����V�>h;�?~��?�oM=��W�Ġ	��e?<�<��F�t�ݻ3�=�B�=�L=��a�J>�T�>̌�[A�^8ܽ��4>څ>�z"���c�^����<8�]>��սf/��Մ?\z\��f�@�/��T���T>6�T?�)�>*B�=O�,?V7H�~}Ͽ�\�Z+a?�0�?u��?��(?�ۿ�7ؚ>O�ܾ�M?�D6?���>d&���t����=�%�`o�����<'V����=n��>�>?�,������O��Q�����=~m�1�ɿe�&������<=�=�*�<'���ꌼ�)�\wݾ8��y��� �=u�>*�(>�zz>��J>q��>��\?M�n?��>�[,>{�)�>���O�Ҿ+����V��c���u��7<�Ծ����Y���*�������ʾ�B=��ψ=T�໎�
#��~i�!�E���,?�1>j�о�DQ�o=�<݊ξ�d�����������Ҿ��/�!i�S)�?n�I?g����S��e�sܔ������ZX?������������>e
�h��<E"�>� H=��q�.���P�P10?�y?�@��h���!�)>"� ���=m�+?N� ?��Q<�T�>��$?Lh,�� 轢$Z>��3>A<�>���>��>����4۽I�?�T?�?�c��b)�>7ľ��/y��Pc=��>��5�Bv�O?[>�e�<���� jS����� l�<�'W?>��>S�)����a����D<==��x?��?B1�>~{k?A�B?���<�j����S�F�Igw=b�W?0)i?ѹ>r���о�~��2�5?v�e?��N>8ch����.�.�pU�0"?B�n?`_?�g���w}�/��>���n6?P)u?:�-������)m���>�?�ۊ>.�@?��q�Z�=~w:?��>�7��<�����!���?6V@�g@�����
��w�=ro$?�$W>Nu��	�/M��_��54���>����,p����ɾǁ��9��>�Y?5��> �Ⱦ�{�}E>xذ�؂�?`�?�n�HV>�۾��j�:��u�G�~��>�Cռ�-d�m 侲�e��>U�]I̾+ ����C=>�j>�&@	��Fc�>�b�=k�⿂����P���Ƽ��(8�>��>�R�����<�e���W��j#���.������M�>��>���'����{��q;�a0����>���	�>��S��&��m���B�5<��>��>鷆>�,���罾ř?&c���?ο\������>�X?h�?�n�?q?�9<l�v���{���j.G?��s?FZ?�p%��=]���7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�[�_?#�a�G�p���-���ƽ�ۡ> �0�f\��L�����Xe����@y����?M^�?e�?ܵ�� #�b6%?�>e����8Ǿ��<���>�(�>*N>"H_���u>����:�i	>���?�~�?Ij?���������U>�}?���>N?�?!�>��?R��=X:����<�n>b�=@Յ����>��G?M��>o��=�&��l5���I�8>N�L��<����>@"_?��C?�Wd>�)��&[��������Ō8�ʨ����8�K�.�|߽�`>?�4>@�>@�Q�n�ھ��?�f �e�׿$���$l���'?j>�|3?_���r<�0���AЈ?=�*>����b����u�+D7�(��?	�@��?��о���vA=�Q�>�?�"�=!�dǾ�MC>��.?����W��|��E��>�)�?K�@v��?q����M?�����	��^&��a����Y"=��=?^U?����.L\>�?�`�>{�~�a���b����>et�?kp�?x��>�T^?�b��8��@;4��>��d?��
?0V������=l\'?�+�b癿����Wp?N�@��@H��?cZ��{㿵���(��+���6F>���=d��>�
� �߽�=2��������>؇�>�
I>,+I>z6�=t�=��>�������~��u,����7�^?�W� ��T�PN�����"�+���澲c־�\��B�J�H/����}��7�ۦ���>Y�5?ƛQ?��t?���>�o����D>���=�3.<:,Y��s>YE?hP?�~3?�0v��a¾1�j��5h�܇��Yw�����>=*�>�>ѽ�>I,�>ٻ��� ���5+>���>U>ֆS<V���ؽ���<�P�>�t�>�G�>�C<>��>Fϴ��1��l�h�*w��̽/�?q���U�J��1���9��ڦ���h�=Cb.?�{>���?пa����2H?���})���+���>x�0?�cW?L�>��M�T�d:>����j�7`>�+ ��l���)��%Q>zl?��f>�ju>�o3�N8��P��a��v|>}�5?�g���]8�3�u�I�H��!ݾ&�M>�>ػD�(T�o햿��~��|i�1Ez=l�:?��?ɕ��Tాe7u����%�R>(l[>t2=�d�=O<M>��e�d�ǽ��G���-=�=��^>�M?��?>q,�=}4�>q���"_����>�c'>��>��A?Ύ&?뢩�뾿�����'?�u|>�5�>�w>Z>�_B���=��>��U>�x,�Ԯ<�|'�-pI�$�Q>��ˏf�D���`�=$_�ai>d$>=d ��m:�I�E=�~?���!䈿��e���lD?N+?$ �=�F<��"�E ���H��C�?p�@m�?��	�ޢV�3�?�@�?(��#��=}�>׫>�ξ�L��?��Ž:Ǣ�є	�G)#�lS�?��?N�/�Zʋ�7l�j6>�^%?��Ӿ�ګ>�q��(����Ł�	e��ؽ�7>6d]?����^���T�ݽ�J1?���>q�Ѿ�Ҥ�{�Ͽ#2z��u�>h�?���?�[� ����dC��c?OR�?��P?��>9��L޸���M>n'E?�N?�>r>�D��@�=��?G�?�n�?��U>;.�?ko?���>)6�e:?��[��엃���;~�=�Ȫ>mSo>�־s[�
�����U���B�}�=�`>��c=l�>`������W`=HG��iͬ��ڽ���>���>��=P�U>�O�>k8�>9}�>����ɽ{��>���G?0�?z����S���E<���;���ޑ�=|\b?�ϟ>),پ���gfz?o�?cd�?i~>*$%��t��-&���y��V쵽-��=�L�>�O�>�)�=���>�Ц���&�>��>8͓>�_�)	�gR�×�=���>�)?^��>��>�� ?P�#?�]j>�>�_E��=��[�E����>I��>z<?��~?.?�۹�vT3�o��d顿��[�a.N>��x?�W?�Ǖ>싏�w���?jC�H�H�(��⠂?+hg?��-?�2�?�??�A?,�e>d{�)�׾�[����>7�!?N �g[A�g<&����PX?��?6�>3����˽��ּ�v�����f�?0�\?�&?I���a�\þ�@�<29�<��Bw<��N���>��>}ރ�A�=gJ>ɀ�=��m��~7���U<2O�=��>[��=L�6����92,?Н�<�ߣ��J����q�']9��\H>��>�v���AL?�M>=z j��W������қ�L"�?~��?Hٗ?��f�Hw<?v>�?�}@?\ѝ>�3׾�u��Y��^��Db��������=;�>8o���پ�����"��%��(�V�a[�l{
? !�>_K�>@�>� 7>A�>��u�Q�8�S����վ�P�Θ)�h�K��#(�h�
���7���Խ"��z>ľy�q���>����V|>��?p�>e�
>��>H�?=�E>��">{`�>��>z T>E�y>�>�bƺ�䣽�KR?�����'�k�辴���X3B?�qd?D1�>�i�:��������?���?Ns�?+=v>h��,+�xn?�>�>C��Rq
?�T:=�8��;�<V������2��}�"��>�E׽� :��M�@nf�{j
?�/?���ŋ̾�;׽桠���n="�?��(?��)��R�|�o��W���R�t��h�h�d
����$��}p��ݏ�e�����4�(��1*=�*?j3�?������鬾�Wk��E?�t�f>���>��>I�>ʓJ>_�	���1���]�eY'����:9�>�{?��>"�H?H�;?@P?�K?�n�>4N�>nv��)�>�as<��><!�>�(:?d�.?JD1?l�?��(?X.Y>?����7���Pپ)M?��?�?�?Խ?���7�ٽ�Ӽs�W���j���u��b={�w<"�޽��}�BK=̆R>�X?���ҫ8�q����k>Z�7?���>M��>���N-��.�<�>��
?aF�>�  �I~r�>c��U�>:��?����=��)>!��=?���>�Һy[�=���6�=�7��O�;�c<t��=t��=|�s������(�:���;MZ�<��>�l ?�:�>$Æ>;�w� ��l���}=��>>�(S>	�>>�*��R#��f"����i�C��>��?���?�y=(�=i�><c���۾�J��m��'ߊ<�� ?͕$?e�_?�&�?��;?�,?��=����񏿹(��U���
?o!,?��>p��l�ʾ��ǉ3�ŝ?8[?2<a�H���;)�+�¾��Խs�>�[/�I/~����ED�E󅻵�����(��?�?�A�F�6��x�ǿ��\��-�C?�!�>�Y�>�>i�)���g�i%�X1;>���>NR?U7�>פS?rv?��V?,Q>�g9�͖���1��\��<j1>�9?�y?S�?ȶz?��>m�>�QB�{��?- �s$��\����'��<��a>2�>��>�/�>s�=s9}�_s���~`�tâ=�#�>�>��>&��>� z>X<��G?���>j[�����:뤾�ƃ�	=�a�u?���?�+?�e=���z�E�'J���F�>3o�?L��?B3*?]�S����=��ּ�඾��q��$�>Gٹ>�0�>�Ɠ=ˉF=�i>��>���>A(��`��o8�QM�r�?�F?���=ƿE�q��p�4ʗ�M3e<v咾��d�ϊ����Z���=Bߘ������?�[�y���b���|W���Ց{���>���=��=8�=���<{vɼ��<x�J=��<U�=�sp��n<x<9��@л������!���\<0�I=E2���¾��z?��I?p�0?�@?aqR>��1> o� r�>ߙ��J?<�S>S��H���>0���������X׾&#Ծ� ^�����>��a��*>�<->���=Bb�<%��=�Q=-?�<�����=��=�p>�{�=�=O>+ �=�6w?���������8Q�C�Ҷ:?4�>#��=�ƾ�@?��>>1������ac�~)?B��?�U�?��?׀i�a�>0���Ŏ�셐=�󜽘/2>���=	�2����>��J>��}K���c��Z2�?��@�??~ዿ��Ͽ:_/>�!/>�e>�pO�� 1��N���Z�6y0��U?OA��(־b+�>�U�=����*׾@�<�+>-��=����]��:`=�\���=�	)=]V�>��O>a� >q��f��=�J=)o�=�C>��{;��t����x�i=���=&RT>�U%>C��>t�?� 2?>c?斯>അ��ھn6ɾ�b>���=�к>�<�=ܽ
>.Ɏ>Q�?@�I?I?V��>�lV=�X�>Rd�>�i)���t�ծ��m�������b�?L��?���>fv�<c�ٽVD(�4*D�	����?�&?j�?t��>�����z�$�?!��<w�>�h>�q���G=�Gr��qվ|d��S5>h�>4��>�Qw>��,>&^�=�R�>���>�>q�1�;��<̐��d�=��ؽ��7>�8>�F��5��[����S�{��{�=�h�\��=#x�=a��n�=F��>_ߑ=�b�>� =�ٺ���P>6--�#
b�'�<C-�Sr7���o�����`�0��B#����>�;�>O�+��0�	?;s>e�I>P��?��k?eY�>[4��W�о�렿�茶��.���=�\�<xrܽ�Q�޾R���W������>Z�>5�>��l>,��$?�x=�⾷b5��>(��ر���}6q��;��D���Ni��׺�D?�C�� ��=	 ~?��I?���?���>C���|ؾ�M0>�K���;=�
�%(q�kf��� ?Y'?ɕ�>����D�MG̾���޷>�=I���O�d�n�0�t���ͷ�č�>;���B�оl$3��g�������B�Kr���>��O?�?q5b��W���UO����.��,p?}g?��>,K?&@?~���{��t���|�=�n?���?�<�?.>��=^�����>y4
?VՕ?���?�v?��8�ʡ�>�45<�t$>�ך�S��=,�>�y�=���=�?�a	?q?���:	�j��9���!h���<�N�=漗>�Ջ>��z> V�=o2�=s��=��\>��>G�>hUh>��>�u�>䍕����Y�+?Fń=���s�-?(n�>4�=�̼�6���y�=8o��BU�#3Y��B\���4>��G>�>�Q�Q�>��ֿ�Ʊ?+��>�~:��7?'A�(K�t��>~9>�Q;�"�>b�?ڋ?F7>�z�>q���u�=��>�[ξ_/7>��&�(����I��n~�c����t�>�H/��T��IM��\&=y��T�����qP��&���j\-�}D=/��?�tɼ�^k�f. ��=�|�?77E>E�[?w���>��R�>g1?��>�9Ӿj���$��2Rݾ�?���?[a>�e�>Y'X?n�?9VX��<�[�T��-v��F��g��PE��h#|��2�xM�۔_?يr?]h2?��y�)un>iE�?�:(�����L��>�B���H�9��=�M�>�_����j�r\��L�����{�u8�>�l?Uy?��?��X���j=g$��V�D?6P?+??��3?�!�?���k?�|�>I�?���>�Z?�C?%-?`>��2=����3[�<�x?��o�d'��Q�Ԁ������=�=(�l>���=M"	>�y�=�p�=��=��=A�r<��&>��>�H�=/v2>4T�>$�]?�>��>o�3?t�+�y�9�"���3�*?� �=̦m��W���o�������T�=l*j?m��?�U?{�f>�;�*�=��?>��>>�`>F�>�t ��[A��ĸ=�R>�>0�=u*�T�t��%��������<��#>8 �>43�>b^9�)�E>Q@��E�����P>H���=3P� �޽֠U�H�;�Dk�{��>��U?S�?fg�<҂ �Y&��]Z��?�q=?nZ?��u?tk=����4�Tl[��q��^�>5 ?>�L�
��� q���V5������u5>]���>砾�kb>���2c޾�n�eJ���羦�M=Ih�nU=�2�B�վ+��\�=�A
>Z���N� �q��{Ӫ��9J?��k==w���oU�MZ��r�>���>��>�:�4�v�qs@�����=��>��:>�L��P���{G�2.�'�>1�W?߄R?ߍx?�E���p�5B�G�5�(�4�V`>'L�>ݯR=�(%?<�>���=��
���&��d\�Y�O����>Q��>���+o�F��ܙ��%�T�;}9��,?�5�>l�!?��>L�*?j�?�G?l�>ߧ>���s��ql&??N�=�ӽ�Q��g8���F����>�H*?'�>��u�>7�?I�?�M(?�R?�?�c>N��;@�J�>p�>ҮW��'��U�]>��J?�	�>k�X?|W�?a�>>�z5����������=�V$>/�3?[�#?��?mŸ>�@�>Z窾�R�=`M�>4�]?�}�?ũs?g�=	�?+�7>���>�[�= ѫ>���>?A?~�O?v�n?�E?���>�n]<�έ������<��,ּ�:h��GA<m�j=9���H�Ȗƻ�%�<�l\<|4��mሼ_�ż������/��<)^�>|�s>o����0>C�ľ-P���@>����N��ي���:�xݷ=���>��? ��>�S#�ᾒ=���>�J�>����7(?��??��";��b���ھr�K��>�
B?k��=y�l�3�����u��h=��m?Ή^?��W�$����b?K^?#F�i=�E�þ��b�R����O?z�
?w�G���>�~?V�q?��>(�e�N;n�/���Eb�k��ζ=Xl�>4V�*�d��2�>�7?w)�>h�b>{��=jj۾2�w�4q���?���?x	�?q��?�*>D�n��"��e��Ϛ�pd?�&�>�ؾ�7?��:�Ѿ���)��3���Ե���c�������t���dO���D������� >�?�Yu?��_?L�^?��㾧�m�Te�U����F��0�s���C�ܻN��
H�s/w���)z�#"���@�<
ln�n�Q�R�?A@&?W�v�!�?H�����ؾt>�r�P�����=Slp���<���=��=�Jb�!.����?�¬>���>��A?��R�ey=��D8�N�A�����3H>tӏ>���>o=�>�ɔ��H@�<;��ү��?��I�ƽ��w>�v\?��G?2gu?eo�GS��c�=���<RO��`�|=��]�3R�>��������/���H���g�Z�̾d�������v=֊&?/k�><"&>c��?�@?��쾦|��A�ľ2	�&��<���>��g?�t�>��=����^:�uǮ>�>f?r� ?��>Ҙ־������;�k�>��$?#��>�ڂ�ə���+S��wx�Nq����_�=��g?�{��6̽@�>�_T?�?���|����>3�M�����s�Ww@�А��BO.?Y�=?�`>�������qY�j�h�0U)?��?<�k�.��a{>��?���>�&>d�?>�>o4���
�P?bn?ԝZ?�lG?K�>&���k;	���A�u9�=V��>v;H>(g=2��=,D3���;�.t&��A=�=�����7�rCx��c<���<�s=6��=6�鿹�d��F�&I�G���G���j�7p����ĩ��3�"�� ��M��>v��ϽN=!����줾�@�� m��1�?q��?�ξ5-���͡�+i	��	^�>g��;4!�s�Ǿ՟��]���`���{���$��SZ�B�a��Ow��M'?�O����ǿb����[ܾ��?��?��y?���U�"�W�8���!>eF�<n����뾙�����οԚ�I�^?�%�>r�đ�����>�@�>�qZ>i�q>p�����:#�<Gs?�-?>��>��q���ɿ���S��<N��?@tUA?�T)������W=0��>
?��?>�21��d��1�����>*�?��?�N=��W�ȥ��}e?�<%uF�l�ݻP1�=�Ϧ=�n=���4�I>]s�>h0�)A�8�ڽ1�3>�u�>�M%��l�^�v
�<O]>x�׽9���5Մ?+{\��f���/��T��U>��T?�*�>U:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=l6�򉤻{���&V�|��=Z��>b�>,������O��I��T��=�:��Eӿ4p+��!���x=���<�%��QIֽ!��C���;�ǳY��r���P>��%>F:;>	<>>]�!>���>�Ll?=d?�y>���=#�I����������J
>�駽
͛��ؾ�N�_G��)�Ҿ��D�%�L�������O��ƃ=v�g��*����F���x�y5?��L%?\�>���������=�[ľLq��#u�=�b1�dl���;��~�ϒ�?��g?.���ۚR�������@�C��N?oS �&�־M�^�O�=��#�=ϯ;?�j>�=&׾{WI��YF��/?g�?a���+_����">`h�.�<C�)?��?�t�<dЫ>$�"?�5������Q>��2>��>��>�>�Z��b8ӽ�c?�P?����u���Ս>�jžL�p����=� >�CL�����.^>�i�<����#s��������<�"W?.��>��)�?�"h��GN�օ<=4�x?�?P3�>�wk?��B?T��<�n����S�z���w=��W?+i?ߩ>br���о���&�5?ϛe?�N>��h���g�.��T�?�n?^?<I��%{}�N�����*j6?,�s?Y�N��<��fF���= ?�>K��>:?�{[���;>I�7?���=\��e���L�7����?�W@@��ٽ�`�ݩ�=��H?��>e��9H�����3��`����?Zzƾ�h���3���̽�?�]z?�'?�þgH�����=���G�?�?	�羒б=)u�%o��t�1<6��%!>�0ʺ�r��A��o]I�����y�оʐ�?=SM;>�@n�p��ˣ>Ә�n�濳�ϿW{z�a���Fz����>�ą>3;����ؾ"�q��fs�Mf6���>��ە��H�>��>����s�����{�yo;�H'��>
�>?�����>ЛS����󯟾
�2<(ǒ>?��>|��>����Ƚ�U��?lP��0=ο��������X?\�?�i�?S�?^@<��v���{��S�)G?:�s?�Z?��%�h$]��n7� �j?�_��qU`��4�tHE��U>�"3?�B�>I�-�Ѳ|=�>��>�f>�#/�v�Ŀ�ٶ�3���W��?��?�o���>o��?ls+?�i�8���[����*�C�+��<A?�2>+���D�!�;0=�FҒ���
?M~0?{�a.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?B�>	�?C��=M��>7T�=�᱾[�3��#>�%�=�?�s?E�L?��>-��=I�8�c/���F��:R����O�C�>Ӈ>�a?�@L?�c>�
����2�!�L
Ͻ	�1�ab켴�?�Y,�T�ݽ�5>�=>N�>~�D�ZHӾ�[?�z����������� tY?��@>�z?x6�(r��<�;ڼ�?��5>�E�簿x���N�ڲ?��@�?چ�����ͼ���>���>1�|��핽a��(ZN>��.?`��P��𷅿�ȩ>RS�?;�@V��?�W��Ӹ?�"��'�����8ͧ���/�V��=��L?�`���.>�� ?e1�>������?1q�=��>=ܲ?�e�?�0�>p�Z?�rg�2���X��<�>{�1?�?���=?��v�>�
?�9�xo��xLܾHi\?P�	@G�@F�_?<����hֿ����dN��N���.��=���=Ć2>�ٽ3_�=��7=��8�w=����={�>��d>&q>0(O>sa;>��)>���M�!�
r��X���Q�C�������Z�7��0Xv�_z��3�������?���3ýy���Q�2&��>`��8[>��S?��<?�Q?.�?�[=S=�?��~g>�%=ʎH=�C�=%�<?�^]?
�A?xW>����3=c�gRy�낻�0}����>t�>�M�>��>Oϓ>�G='>{�o<��n>���>g�8=������H>qh�>֯�>/>r>m�0>&�>3���᯿mhk�񊅾L�޽C�?3Ɠ���M�;՗�32��;5����=�d.?���=Bd����Ͽl�����J?����M]�z�6���>{�/?;�T?[,>�V��(�U;6>�'�<�j�ߪ	>z3��&y��%���W>��?��f>P'u>I�3��Y8���P�V���U^|>�16?�඾�;9�+�u�X�H��[ݾS1M>���>~�E�fo�����M��yi���{=v:?��?���~ް�d�u�a;��0>R>+\>P�=|g�=�KM>�Ac���ƽ�H��1.=���=p�^>�8?��/>n�=K�>�6���&\��>d�;>��<>��@?�v#?Fy+��-ý����R$9�M�r>Tc�>��>٣>�IN�j|�=k��>�AO>K��Ԃ�ߌ�_�X�Ib>�,����f���Խu=뿁�P>Y�#=�M�&t4�G�&=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ˧�>���ƙ��J@��+aa�ڈ�<�O�>O�[?�PǾ���Z����+?Cu�># Ⱦg���Կ>x��r�>;<�?]*�?��c�����L�^��}?t�?�U?�q>���_sٽ�A�>��M?�}H?�1d>�.O��'��K?k��?͔�?ѠP>��?8%q?�`�>]�t�3�=��꧿M���gj=��ٻ�.>��*="e��ۆ?�<����Y��P�m�%N�Bm0>T�<qI�>\������U��=R���=J���%A��ٛ>a<|>��K>xp�>W�?��>�:�>p-	=�`ݼj[k�SΩ�ބJ?�<�?���p8V��Σ=I��="�zΓ>��@?�u>�3Ǿ�L1>,g?�G�?R<o?1D�>�4��z��}#���Wž�rj����=v��>3��>|����>���ҷf��Ś>>�]>�>�;�Z꾷O����>;�|�>� ,?���>�2�=ˎ ?a�#?1�j>q�>�`E��3��O�E����>I��>�1?��~?��?O���^`3�K���ϡ��t[�7N>��x?BC?&ҕ>W���Y���&�C�K�I�툓����?g?m��t�?��?No??P�A?&�f>D���ؾ�d��d�>.�!?��ĂA�}'&�Ƿ��{?b?&�>�,����ҽ*�׼������4?G\?�S&?���B8a�f�¾B��<
�(��I�	�<BD�D�>�>�򆽐j�=�>���=� m�g�6�g�Y<v�=.��>��=��6��ڎ�aq&?�W��Bʔ�M�T���\��L��u>��>.���Y?i����=�2���pꜿd����?^�?四?e,��)��{�0?o�?��*?�a>g]ξ~8������p�����cӾSb����>,�����֛�,��9ё����}�M��� ?��>��>�4?.��=���>p�*�AkD�N��[�߾Օ`�D%��"R��>��o��"�b�M"��Ⱦ��z�Z��>J)m����=k�?̙�>�r#>��>�R�=d�u>hY�>i��>���>�>��>U�&>:�����;�KR?����!�'���达���g3B?�qd?P1�>Pi�:��������?���?Ts�?'=v>h��,+�~n?�>�>H��Uq
?bT:=9��:�<V��p��3���3��>�D׽� :��M�=nf�vj
?�/?�����̾�;׽N����k=�5�?G�(?�G*�{)Q��o�x�W��S���"��f�&\���%�d�p�E!������a��^#(��-=��)?��?;��]�(��F�k��@�?�h>���> �>��>��H>��
�Y�1�Vr]�}�&� ���G��>9~z?I�>P7;?��9?agQ?u�M?GU�>|�y>�ʾ{?}@�<"��>
}�>3	H?��'?��8?"�!?�,?�9>р��7�X��G� ?�� ?��?4��>z�?���Gٯ��C�����~8���5z�̈́W���>�Xƃ�^l=�"Q>�X?	����8������k>�7?��>~��>���-�����<��>
�
?�F�>% �.~r�c�JV�>���?T���=��)>���=뉅���Һ�Y�=������=S8��{;��f<��=���=HAt��ہ��!�:$��;!k�<�d�>!U?��>Ypg>�g�����2
$�`Z�=��u>��">b�?>0L���ҋ�E��Pvk�/��>DD�?:�?w(>	�=��>v�ɾ��!"�_輾�GX����>Q�C?Bnz?�}�?`�?��?v�>#;ƾ����H�� ����^?n!,?��>����ʾ���3�ĝ?`[?z<a�׸��;)���¾�Խ��>�[/�i/~����6D��腻���2��-��?⿝?�A�I�6��x�տ���[��u�C?�!�>�X�>|�>C�)�c�g�y%��1;>��>WR?�e�>�d?�l?�KE?Q��>D]-�����X��H�>ʹb>g)3?��>?�x�?�a�?�-�>ۣ�=�ŗ���ɡ�.yw�I
�������w���$>��>���>٘�>�|�=î�������	�܎S=��>��?}�>���>s4>yev=��G?���>�O���������΃�uF>�!�u?���?��+?��=
w��E��S���$�>�j�?:��?�-*?�xS���=�Gּ�ﶾ�r� �>�ʹ>��>���=��G=��>���>\d�>_+�5S��U8�{DN��?�F?4��=n ƿ͢q���p�����gd<P��3e�����{�Z����=*Ř�m��-Ʃ���[��������k ������.�{�>��>(x�=
��=��=��<iKɼ�½<$�J=���<"�=�Rp��Ym<��8��]λ򛈽�j�=\<D�I=.����)����{? J?E0?V�<?vh?>��	>i�� ْ>`P��5�?;t/>M�;�9R¾Hd1�8�������<ݾ�BϾ��c�癜�g4>��8�؇!>��:>��=^�ʼ���=�7=�~�=n��;�Y*=�r�=)Q�=�y�=]P�=��><��=�6w?W�������4Q�Z罣�:?�8�>{�=��ƾo@?��>>�2������zb��-?���?�T�?A�?Cti��d�>J��i㎽�q�=i����=2>f��=~�2�T��>��J>���K��<����4�?��@��??�ዿТϿ5a/>�4>\�>�FR��X1�<aX���a�RsW�͇!?v*<�jB;�
�>q�=V��B�ȾJ�=�3>��o=F���\��G�=vc|�� ?=��j=���>��F>g~�=M�����=a$R=���=P>���93�3�+�/�n�>=���=Z�`>�-(>���>�N?�'/?X�_?a'�>yPu��پb��	8�>vأ=��>�ޙ=_#>� �>Ʀ,?y�E?8K?z�>8d�=�Y�>��>z�2��mr��d۾�ɬ���߻�M�?�"�?,w�>"/<*I��Z�=:�#F��dM?+�)?�?��>5���	�'�,�%�.;�J�&��ڽ�������0�Մ���O�&����,>^�>bW�>c	�>ثU>��>=�V>��>�{�=|���sͬ=����2X=�#���=)�=�^�C��ٷ<�x$�H+`��(��kK[���Z����2}=qoH=&9�>��=x�V>HW
>�X龂iP>�w:�܏z���^�.3/�d,�������k?��{)�V��>�;�>YKS�]����I ?��$>�8�>%��?
k?�>�3*�ƙ׾�{��e�e���:t�=;��=LVI��_��j���P��վ���>��>��>�l>�,��2?�/v=���U75��,�>Ӆ�����M�L4q�>0����i�IP�3�D?�;��а�=}~?Y�I?�׏?qr�>�����ؾ&�/>����I=���q�����?z�&?�U�>D��K�D��A̾� ��f�>�6I���O�߿����0�!�t˷��}�>>쪾��о(3��g������J�B��0r�R�>J�O?��?Xb�Z��w\O�����\���c?�g?�6�>-M?;?�0������p����=��n?���?�8�?q>|@�=�fǽI��>1Z
?���?�t�?�t?� 8����>��;{,>������=�5>`��=g��=QC?A�?��	?����w	�II�)n���m���<��=\ߎ>� �>v�w>O��=�k=IM�=f�d>K-�>�<�>�g>9�>Ɗ>$ʥ���d]?a;:=p���T�K?ru�>�u�=`���!'�S�h>�j�������)�����,m>C�>>�]>W�y=�	�>�%ٿ��?��>�B1� �:?���C�꽘vr>rX�=Rq�=vl?���>ZZ?���>U ?��(="H�>��>��ݾV�D>�'��@"���P���g�ZQ����>�'�o�����!�C��R�h���z�ϻq�:ބ�O�G�X�Q�"��?Gݽ,�_�k\9�s�	=eZ?���>��B?:����g�<�k�>	�?Q�>����� ڒ�F⭾ߕ�?P' @�U>8̔>a6U?�e?,�h�i�;���\��Mr���=���e�bMH��<��������^J�a�Z?�s?f�3?�DA=�\>���?Z:��ZǾP��>��;��L���>�'�>#����o��ľb��D�6��_U>��^?�]n?��?w1���>s�!��.E? �e?�uc?38?9 �?"e�=WM�>+�>Ù?���>�pJ?	kM?�>N?)�o>��!=�X?��T���*՛������+=[p�=�Dl='�ؼ��#=�Z�=7�<8
y=.�=IƼ��ͽ�fG��#m��[}=3�>��>�Q�>G"]?\��>�v�>m^6?6��9R9�C����j/?�H=�G��d3������9��c�=�-j?)t�?��Y?�g>ԃB��@���>�U�>>�%>E[>�>S��B�A�j��=#>�~>�h�=E�Ԛ~���
�*�����<�>���>T:|>�č���'>'`��Yz��}d>R������S���G�>�1��;v��]�>r�K?��?���=�`龓����Jf��)?r`<?�PM?��?
�=̹۾��9��J�XG���>��<���¾�������:�)�:x�s>�&��
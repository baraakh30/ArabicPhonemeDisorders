`  �   Y3�>F�j���10?����9��s�_=�=�� �6/5>)�,���MeA���������~;�
�??��?� ?�[?U��,�Q��6&>=�e>K�?� �>4^�=�ڃ<�#>���>���!��׳��E??�T�?�@�uy?/�a��п���7���Dj���#<���>4�>���U`>M��=	���knc=�R�>��>g��>��>�u>s�A>��O>�~�i0�=ޚ�BZ���o��	��J�yv����c���1��e�=�Y��ܽ[��gG�<���H�a��ֈ��#����w>�]�>�:�>3��>A!>�f�>���b��B����d�������־���������h�*�9,"�oTv� �ͽ�������>C�ؽ�CZ>X��>�<�&�">R�>��=>"X>���=<J�<�S>���>��X>�+#>`��>*�>,�{>Zݎ=~ㄿ����ӻ9��R��N�;a�C??-`�����3���ݾ2�����>Ze?&RQ>�'�y����x��6�>,uB�	&a�/kϽ����p�>�S�>�z�=��������%�v�˲�/�= υ>��>�^�pȍ�)��Eړ=X`�>ƽ��y��<'U�<��G?ef?��<?��=�J�>v>
�>	��{	>~�>�g�>1��>4?�"?�d?̇h=�J>�0k�=��D<�D��
���TN���-��m>x��>�m=L_>��=���=�L>���=|v#;F��˩<���>�^:?�_�>5 �>��?�p�?���G��w�K2�=5�����>��>���>	��>���>ٽ�=E\罜¾�xϾA�>g�.>K6V�0Zr�%��T��>q �>�Q?��&?C�нE#o�8�=���=佽>��?q� ?۞�>�1?>t���!��8ҿ�P۾�?&��5 ��o>V�d���`��=�f׽׻���>O5�>��>�O�>Y��>�x)>��{�P@0=���>��^>J�=����B��=^{�=��'�Y��=5�,��J�=ZO�<5=�<o@ʽ��,� 2k�h	�r׮��yg��Q���[<?�i�>hi���>����/��R���?U�e>I��>d�@?.�">�{"�N>���Z����߾'~�>�W?�?d�R�S��>�=yqH>�(�>i��=A�м!�=��Z,����<��>�?p��>�Y�(�������'����>ch]=�#��Z�?�ND?I��~t���e(��eP�����=Q�P�Rfv�\����G+�)TH�����9��.z��ܴ=�?b��?����WH�=��̾��؋���[���w����=��>�&>
�u��:ž]���Lʾ��%���=�|�>��]V�>b?��>N_u?V�?�&5?ekf�N-?�Ь<.>>��K��?)H�>>�>p5>�>��<փ��W����|�y{���ug�l�\=��w>-�P>��=�>�$���4��.���dt=���2ͽ�Q=���=F�8>Y��=�6 ?EG?���BR|<�9�OͶ��1.�?��=��
��H(>�����@>�>��$?�c,?`�f>�v�_�8��cH�h���>��?�-?1?=%�=~��=.��olA�R�=1�>�����2� ��A\��o��DF�>�l�>Q�=��>��|?�,?&)?p�;��"8�=�{�Y��(����:�os�>���>%�a=۪̾
�5�k.r���a��+@�{��	�Z�n[=m��=�t�=�S>�=�W�=����$��Ʌ���J;�h0�Í�>��> �?�>�d�=������(9s?�𫾬ue�򠥾�*(��!���>��&>�p�=?[w �?2��FǿKwX���>��?vy�?H��?5���}�H|�=}e�=�2�=�s�W����3>���>���>�q>�_�>E��;6-�<&�)=wh��2�m<���H��}�>�����V���P>���J������g�׾�w}��v�Ā�'���3X���$��B�-������P!��c������땭?�ps?p��>�� �W���(� a�f��0\	���X��A,�IG��0��f?'�Ӹ��=��+0��q.�@�p�>��Q�4����yt�y
)��* ���7>�l2?;і�����,�=ܷ>�z�<U��G"�������<�[?�38?�i꾍������k�>�Z
?��>��C>�˗��������>��6?<�/?�(�;�=��<����ټ��?q|�?5O?�;�F�
+�����X>�I�>�M?jz得&$�Ǟ=1�M?�W?3k?y��捿�k��ׇ>(}?-]�e�>�t�>��O=˶�%���Sݽk̾ܤ�=f�>�����v<��p<��
=�	�=I?�o>��$&*���>%�-��*x ���B��J�󆉽�v�>��S����>r�\>�`C>�_)���4}���b%���S?��?�)/?{N?�e��AJS��܉���s;{��>�?}s>8&�=��>�� ?���%]�c����>��?��?��?l�$�^y̿����x�������>�?�=b�i>�[�V�:>�0c=��7<���=8v>p��>Ziv>�7>|X>%>�Z>�ۄ��+�;Ş��h���B�����w����
��e��I��q����B��P���3�|��1���
�n煾҈>��?X�?Ŧ�>)?G>>�=�+���q�;����jؾm�%ﾧ�۾�谾��d�Գ��������6�����0A�>��=u�>�L�>��<��=D�>�7W=�n=a�>Ƈ>x�U>S�]>�;\>��'>�O;>���=�|�>U}��7Ȃ�ʂ�":@����^h>_`a?���X���/���@��4ž�!>׷+?ȁ>$)�
�x��c:��"�>��&�籏�^I��|�޽G�>E��>�]3>�J=��<X?r��cA��z�WU>��w>{|=[!W�������C>��?Jɾ>����n���>�>�l�?��9?�̳�ì?9�>6��=Qe�J�=$	�>ҁ�>�#;?U:B?���>��?��=��� �=�s�=���N'�8K��bQུ�%��h��e���!>#ձ��\H=��(�	�=ǟ��2�'N3>q��>�&?�I�>M#	?����%���B����Z$=@1���=�{�>���>��>���>mAM>d�~<�䉾:���K�>�z|=!^����TԢ�U��=L��>�X?܌H?g*>��
�I<����/=�>�?!�?�J>�v��ao�=����kӿ$���!�\낽!W�6��;+�<��M�s"�7��-�����T��<I�\>�>�p>mE>�>�>3>DR�>VIG>P҄=�=*�;�;��E��M=���>G<��P�7u��[ Ƽ,�������I�L�>�,5�'ټR�?��>Ag�`���a�˾UM/��-���J?�Tn>Ԏ�>��?�؇=Y�,�c�R�<��o�~�>��a?u�>M*����>F)�=��=>��?�$�>𸽚w��(�`�w韾�m�M8?��I?�}�>�A�9<m���A�Na�$6=�0_=#�;;��?	rX?~���[����-�1�^��\'�3B��|����i��DG���^�>��c��\��4Q��e>�T�>�6�?�]K����=��4(��͉���꾍�:!��Fz�>�>�-�9^�6P�vl1�$X��E���rT<w�)��?��?��?J��?"ۊ>��>��`�oR�>�o����?.?;KK?-.?4��>T�O�9�N�H��������˽�~���3�=Cˏ=�G�=b�g=���>��<�=���=��<����<><?1<<s�<ټ2=.��<�>��>x?�X�>Q)j��0X��>�<M_�=�^3>��=� %��>�r+��]����;X1�>�8?�;?%w>å����=<Zپ�ϛ>��?��O?T?.������e�����ߘ�<��=�94�Mhy����PLҾJ[[��>�ĥ>V�G=T�:;�?�)?�?y��<B� �M���������!j��Ө!>�>�o�>e����qG�p^���\���f���Ǿ�腾�l�=OJ>D�1<���<(�FUR=��9>�U==[;(��X>F#>�k�>�D�>t�?=c>��B���Ӿ������Z?�� ���G�N���#&�o5]<r��>��>�U>�D�>K&Ľ��l�ǣ��3W�Y�>悭?V�?�Ӏ?�&<뭋�"�j>�>�<�����IK�T�������<G6����G��T���o>1�>~:��eؾ�H�]�":����B����>*ݪ��1���x��9�徨[ɾɎ��_�ހ��`ͽNX�� �3������mV�/�Ҿ'��?d?�f�>��@K?��u����XV>�6g��0��׾��2���Ǿ��򕢾� ݾǒ��dt�s�Ǿ�>l�Y�E=���|��(�ᯓ���?>^;/?o7ƾ�ƴ�(v�*�h=|!%>ϓ�<�gﾎ���횚���
�ZW?g�9?N(��� ����>e�?�j�>6S%>q����g��>f$4?)�-?�����6��G*���[�?���?[`C?B }�:C�=g�A�h����>�?��>���-~���>���?��%?��>���s�t���	����>�0]?��=���z>i��>=Ɛ>�ɽ�Z�J��E���6ϼ�S�>f�E��/�A_��O�p=\==�~>z1�>�6��U��
��>����j�Z�F��P��J��<��4�6?)�h�Y��>��?�O>�P�c������+<��?v�?)|J?��V?S��XJY�]=�򄚾;�����(?x��> �=���>��;?�^�g�Y����H��>���?T��?~`b?�5 �8Gӿ��������P��=�$�=��>>��޽�ɭ=`�K=uΘ�8[=���>���>o>7;x>|�T>��<>��.>m�����#��ʤ�5ْ��[B�� ����vg��{	�oy�����ȴ��񽾈�������]Г�j�G�Y��0T>���žf@�>�?N?k��>�MC>��=x|¾���o8��V}����ߜ��f��_O��=���7���+ľ[���-5��1,����>ke_��}=�=�>l���5�>��>�c@>${>��=��=�Q�=r�=ՕQ>o3�>���>��>ot�>��M�O����#���O@�s\����=j%J?V�	��s1�ŐA��_�~~����>�?���>#c�w����a��6�>�,j�W
p���޽$����>B+�>k2�=�G˽Mz���u.�`�=�M>i�>&�9�*Ú�ù��1����?���\V��=�?�|�?��?�i��Ў�>2�����>�t�>�ɾ�
A>���>��?m�?��_?�?#�C���+�>���>�P�C��9q�<�9�{����Ǜ�@�=�5e>���=��c�T���&�}�ս@p���.<T��>߈9?.��>,��>)�5�Y>�)EM�����>q{!��%�>��>�P?C��>�F�>_t1>A_i���ľ�b�>H�>��>>��^��w�����mx>�u>_O?s22?�$i�
:e����<6N�=L�>	�?m
*?;�>_=>�M��|(��]޿����E�������<��!�̲�����=w������;����p>0��>y�>�/j>�f=fa�=T�>uu�>��,>��
=>�[����=I@e�ػ=�">�)�����Hd�o ׽�Tʽ�'��"<{�=���<���=;�)?Ye�>�/���vV�@(ʾ�^�����D?5��=U��>� ?��>nCپh\\���S�E���%?Y�D?��?�>%�[�
>>}��_�=5U�>t8�<�݇�x��A8��U'W�9��y�>��m?1U�=�誾r�x�sx�O�9�Ksq>��=hط���?�V?m�u���a�&�ǣF��k�C >�+�� �DR�`b�WBG����	�xI��h�	>咺>�@�?�Ę�Q#��j��������c���ݾ��e=��<���>:�>�̽g��D� �����c��خ��7dW>6���_
?}��>�L4??|?�3�>ܻ�>�7��=?4%K�ח�=:_>�3?iy*?ĭ>qc=?+/=M�kw��ww�kM����=-� o<=b��=���=I�=��M>��v='��=�I<'���k�9=J�e=���<yޞ���=�->�S?1�+?*ؽ��:�Ks�3��;��<ҹ�=�>�����΁;�Nk>��?��)?���>5�A=�[�)z�;*����=3?*�.?���>$�E=�T>a������� =_�<>�PĽ�U��,�ᾎ���n��ɰ�>�7�>*�>%`:>���?q�>��?��=<��愿8�F�6>	��e�)lH>XC�>�=�>���sG�Iߞ�Eꈿ9�{��K����E�>8P�=�cl>��W>:��=�$>/xH=����:�2��Id�����>Ru�>��"?�Ԩ>��=~�p��!�a�Y?���ܗ0��r2�5!�.9;�?-��>*XQ>�W1?�Z��ȋ�HĜ��r�T�C?��?X}�?�Nw? �>�B���i>�n�<�~����>:�}>��?��T���=\s�=3��X���ӽ^�?ɬ>+%ƽ�ƽ0<��� ������<�x�>qz�̆?�Sr���"�1Pؾ�(������;�Ů����!�����!��W���T��־�������?<��?ب�>�ʽ@����|���D>ez���n=��q��0�(����������B���$��������֛>-�Y��'����|���(�����@?>�D/?W;ƾ|����h�>�h=�B%>�]�<j����������
��_W?L:?�9��.��p��Bi>M�?Q�>�c%>�5��Z���>�G4?�-?��r��*"������^�?���?ilE?�͈�hzB��������?�>ϵ
?-i�>��n�'��oͤ��8?pK'?��
>&��3�d�.���>'�\?oI9��=a>`��>㐡>�,v��34�L����ٹ�Y4��K�>�q�0��h���S4�oq!>��>g��>�_�q���N]�>2[���8�����G��c�����<�y?��]����>�>��5>��1��?������$����G?�C�?��h?�~A?�ܼ�dWq��˼�b���:
_=��>��>�ӽ(�H>�G/?������n?���?�E�?MR�?6ij?�:F�&Jؿ{���|$���յ�v�=�}=4X>0�޽<&>���=�6�=��$=]�>�Ū>��k>g,R>��>n�>a�%>����a��D�� ���q1����Y �]�;�iԾ]�G�����D����¾�_ҽA8�����MlP�z��@����Ǿ��>�+?��
?rd�>��>���<S똾r%Ҿ�z���	�'��$���Q��S�Ͼm���`����N��/���4]�=���g??����<.!6?�%�=菹=�,>��\>F�H=�WZ>ތ輾��=�%a<��>�19>�i�>-��>'�> �<t�}�c_����?�Pd ���f=Q4?�?��)S��0>�բ����$ҝ>ݹ&?#u>%�������g����>Q�����<�-�M�����E�>�i?Ƞ�>��q=�f�;d��������j��=�N>���H}g�J�����<>��>	N־H5�=)�s>�(?r�v?��5?�/�=� �>C!^>6�>��=�TH>ǚL>:�>7�?�L:?�2?\�>	�=g�^���=��@=��=�+GZ��������k�'���<q�1���T=�|=�#<�hH=�8>=��ļW�x;��=>
?`�'?-'{>�L�>����w���7m� �侾7�r�ݼ/;&>Hi>1�>G�"?�#?�T�>�;[�2>����L��>��<G,���������M>��?b�z?��a?g�>�Z)��Hڽ�9�(�_>\�>"��>ӣ>H��=�A������˿s�����ܾ�3>�����罐�����>�+�=��>�qH>�<>�!�>m!u>�|�=��K�S9���)>r�>��>b۝=+��<ަ"=��=�󃽷Ga�~ս�ﲽ��2�;��=�5:���g��=�#�Q<XcD���=��&?B[�>�X!����d�^��Wp�a0	�q�?�a_=Pu)>��?�.�>9���+l�h�F�!nr��c"?i�K?A�?[���X>ʂ=���=���>�G>�2�>@�p;��k�+��;�=�*?��Y?V��>:B˾��'R�h�3��ȼ>t�w=�b[�jk�?j�P?Z� �'�r���3N���޾��B>�]-�^�"c����!��?�x��9_	�O�E��4>	,?�?�@��9>�
��"��N{��3w�Oq>�yi=g�?Nb>\0R���Ծd9��霾����@�(>���>�?w�a�?6��>?$�>�@�?��?�?GN���ν>��j�~&�=��v>?�L?�U?>Lj��:�=����,�>�C� �z���=��,���=r�G>�޳=�� ��Sm>��=K!r=��<i N=,>?F>�v�=� �Zu�<wt>�?��?�FJ�Db!=�g=�Ļ����� W������*���׾�[����F>�$ ?��R?�*?�!S=���pB��7���WY>Jn�>w^V?]�?B�5>G����8�k�^����<��>�t��]X�a���}�u㬼��A>М>�g�=�%>g�?�c?�>$?++�H�FJO�߾rWY��ڽ�X�>��>:�>�\��7)�~V��I��FI�q���ؾ^�X=���=�-�=���>Ɗ��!А�54�=}2;�����	��<y�����=�ň>���>�f�>�q
>��:��-:�\?��)��;C�\vR��F��4ξ�Ի>g��>�c����>s��=�Փ�ʰ���a��<�>g�?(��?	��?�`ӻ�J��K0>��=WnL���>c���լ�Ό�\
�����@h���kJ����=z�>nN�=�?��n��ϣ�7f�"���Y�;��q�>r���L.�PY�PR�h��~�n��������(�������!!���\�ԷѾ&�ľ�O���z�?�^?ux>�h�<#T���\6��d*��d9x��]
�G���D�ڵ��E�p�þc;��ݏ��Ӿa.��q�><�[��I���{}�s8)�7�S��D>�G.?/Bľ�񯾝F��F='/ >7��<��羨q��,͙�\���U?��9?�U������｛|>�?SB�>E0>ѐ��J�齳%�>B�3?�g*??h0��I��3��0�W���?��?�??, K�c�3�֜���D��?�>fk$?9S�>y¾�q��6ؽӆ-?�|U?Mh�>���֍�|��o�>NJp?Aћ��ՠ>o��>��>LE���C�q��2���<�=�H�>��Ӻ��D���mn��@!�=d�@><J��>꫾�{��.��>B2(���پ(1���B��%������9�>� ���x�>�2^>��= $������
{�D���h27?6��?��?�Ł?+��3�������	U��t�<��?R->A���>��,?!G��ʄ���3� ?���?��?���?|���cӿ��j쵾�X���\�=�v�=�?=>��ě�=�}F=Sd���D�t>�;�>nn>�vw>��S>�<>��.>Ԝ��%�#�Ω���ڒ��:B������g�.a	�!Ay����&�������Xا�����X���jG�����=�L�.>!�%?���>,[�>�zv=�=����2���R(;p�ھ���n�о�pϾ��˾,������9��?�澈,}��T"���
?^�=�K�=]��>�^��h8>��>v�=�">�B>V�>��>�� >�H>��	>��A>;�=UC�>/�<�t��׃��.;��+�F�;��7?M�p�2�p�$�?���?���Պ>�0?�!w>ټ�0��I+e��O�>u�ҽ�߀���Z�C����ܐ>u��>\�N>���<�Ȼ�RH���ὑ1ڼ�^&>p>P��Q
4�q�����=W�?��\u��4T�=�"?G�?q�?�>!�>�&>	V�>¶O>�'T�A��=��k>�?+�e?�:=?F�3?��=�ټ���'>?u&>�ER�BIR��h�{KK�s�������>R�<�R>�>�+���S@�߽_���7=M%<(?}1?��}>�4�>�Eҽ���@�s������S��[��r >�Y]>���>`<??�!�>�=Ƚ�~����`�>u>sD9�⌑��F��ۋ/> p?��?w�d?��=����w2�zO`�I�@=c��>��>��>#^x>��=�+���kӿL$���!�S���ߏ��K�;`�<�U�M����6��-�����£�<3�\>��>H�p>��D>�>=3>�S�>PG>��=
��=�ʦ;Y�;F�A�M=8����G<ܵP�H+���.Ƽ������d�I���>��6�yټ�B'?F=�>"���sh����h�/����Z]���>�$R>��$>9z ?2ؽ>���+W�X�g��񛾖��>,]?�?%@H�-��>V��<�ɕ=�mX>UuU��K>��2�)9���+�0���I�>݃d?�/�>��Ҿ�킿����m#��>��9=߬�:�?_]?!�E�}��"���E���
���J=���=�V�<*��E!��Y8�t���c��t�pp�=Ҹ�>�?����}}�=3���1%��^t��^<���'g=��=Z�>�L>#\:�O ���D�8;�G;�L�=9$�>�H����+?M)+>�J)?!v?���>a�?��V>Qy�>��=BP�>W��>�/?c=�>�W�<>]�+e>�X˼�9=OBr�i�C� I�=�^9�<;AE=�L%=$����\>���<�M�=eE�2�;s!�۷^<�ߛ=�\f<��R=U�,>�?É�>G�|�B=s>�*�=᠈��'־�ʾ�i���޽ZWԾK����> �J?�`J?vb?����.��n�%��KJ>���>K�U?7T7?�Ï>@�u�P�@��G���a�X��=�i����AL���P�x��=�A.>uW>�[�<���>�?�F?e?�V�Z3��1<�x��L��\�>n�>�=?\�>����H�K�Ι��Žy���F���e�rO̾*�\>s��=|C->ә�>y`;>�@ټ���=EX�'���4W��^{���={,�>��<?���>��>pwK�i:���a?U���<�~S���Q�V�y�R��>ӵ�>̼��8�>��d>�j��{/��Y��S?�ǰ?$�?TJ�?��f�1܈�z@">k��=b��<h�r>z<=�0�Leƽ��s=d��=�V��&'���z=p��>F>H>,�ƉJ�P0˾/�>5�ο+���.?�l ���žPt+����?���JK>�d��tM�bWD��yT�ZȠ��tF�n��Rw'���	���Ae�?mr�>6�Y>�ދ������]�W摾9�!>�t���"~�(������;�G��b��wh���:ӾDa �c��7��ٵ�>�&[����7�|���(��d��,�>>͘.?#�ƾ�����P��:Y=9	#>r_�<z��W��+������3W?��9?����{�����8>�?���>F^*>����-���>��3?��+?�v�����w(���w[�*E�?ݍ�?��G?]����+������'�Ȏ�>��?BP�>_Ȇ�jB��<qc�X�)?�>?<�>��3��ό�n`���>��^?f܇����>n�>��>3`�Èɾ���[�����g=c�>�н�A�����1ϵ�w=�>a�;������g���W�>g����ON���:����^5��'���*?@�����!>���> /�>ӛ0��6��֊���}���=?�w�?�`?�V2?3	�uҾAU?����=�+�>Z��>ۼ2>�� ;�:�>�W�>?ٸ�>�X�n@׾l�?��?���?sS?�o�7hͿ�ٖ�=t��5��T=�=�dQ>:"p�5l=�`�=-��<�+�  �= �>s?j>��4>�=W�8>��>����%�Tp���]f�XO��*���<��Hf�ۻ����P���x��^.ɾ:~ �������YK�����׋�p�=?�l?�_�>wXN>��=���lվ�`A������ھ��둯�Ϫ��'��fH&�9 e�
6�����=�q־��?�=�=��`=�U�>�����-�=MК>E̓=d��>��>vn�=�=>�Ҿ���I>+�->{��=3>���>��=�菿����έ=�_!��cK�J<?Ó���~���Z�x׾�f*=�b�>\s$?g:�>���?������z��>��8=�n�ϬF�3��=��>B�
>glr>�4���L��N	��ýx+�Zn>�ܐ>��>ox�e.����C�>���}��=(Q>_#)?R)q?1�9?ҷ�=�]�>yS?>Q�f>=}k=³o>�H>�&�>$?�)>?��(?F�>Һ�=��O�-c�=�4=��,�T�<�(z����-<{�^���%=A�=d�=���= �L=���T�Q<.�<0c
?�r'?xԂ>;А>;䂾�D9�n�7�oi��Q>/�a=��>�p�>t�?���>-ɩ>uF�=|r��7����)ؾGR�>�r>�vB�����s�����>�q\>��W?<�8?L$��>u�������@�>� ?J/?��M?��>�g1�ː��� �M�ѿ#!�f��� ߺ��=S)A=�����D�s����P����������a{>�W>c�>`}ݼ%6�=��=�R�>/��>q�h��w��e�="�q=S��<iDG=?� ���=]ީ��d�=d[�p�o!���t��=�A�=[D��&.?j�->]�z�StE9���=�\�,w%���?�>?%	?n�<?��?��H���5���h�F,�e�>}rj?#�E?���T�=%yH���F��c�>�*�>�>�\��3����X�
藾 ��E��>�|)�
�����
��,d�������>U�<��"�j��?oLQ?y����}VG���J�уݾ��
�5�3=���p�4���H�;pʾJ��ʷ�Tq�={�(?�k�?���4�{�&�*�����H���]���9=�� <�u�>�;�>����������0�8��⾺\Z;�� ?��c<��D?��?�)�>�7n?Gf?�P?zPռV}>��p�{���� � -?��?�=?�>$?~<>h=��W�L��u|���)>7Š=�n�=T��<�~?>���G�>�	��<�y_�����3�=(��=s�D�MRP:�C>e�=�G?��"?�ξR���	����4=�➼��>P0��W~>R<P��%��-�>M�m>��?�Q ?��>�$޾*:�������y>Q�3?-D?��>*�"�}�t>o��Z���X�>�T�>��=�j������վ�񋾔c�>)��>�xi>kNm>;�|?
�>?j"?�q���,���u�f�,�*�޼���;7�>��>G��=�a�
�7��s�#�a�+1���o�E���
=L�=GO>�?>���=�E>��=/m��c�ؽꬓ;~�_�� �>�]�>�$?�X>��u=G7��g����I?o頾���H��D�ϾG��>��?>����?���}�溥��=�,^�>�a�?��?�c?�E����93]>@X>��>$�!<#-?��4�]���D2>:�=5Mx�9���;��;V�\>2x>W̽3�ɾq��cBB�f���JH�����Ġw���Y��~�����z4L�����s��ž*��9����:�I&ؽ���'���b��Ь���?�r�?n1�=�x�:�G	��Y�.b�9�>:�����M��������>��a����\���Ծ`D$��93�-R����>_�Q�e·�O�^��'O�?��ـ���?�����l~�C��>	/���@4$���/"��a���{?6=??qJ���1�|��\���I�>˪�>��	?3�<�뻾�>�Br?4?2�M>N`�6����J>9s�?�}�?j�R?7W��^�,!¾$ɍ��i>ID�>��>רr���N�~��X��>q`�>�d<���K��Տ�r'E����>>�?}�����>I��>�K>���=3K�<���=svȾ�׽N�>����ܘ��}+��i���g>�f�>]�%>�ބ�H����W�>g����ON���:����^5��'���*?@�����!>���> /�>ӛ0��6��֊���}���=?�w�?�`?�V2?3	�uҾAU?����=�+�>Z��>ۼ2>�� ;�:�>�W�>?ٸ�>�X�n@׾l�?��?���?sS?�o�7hͿ�ٖ�=t��5��T=�=�dQ>:"p�5l=�`�=-��<�+�  �= �>s?j>��4>�=W�8>��>����%�Tp���]f�XO��*���<��Hf�ۻ����P���x��^.ɾ:~ �������YK�����׋�p�=?�l?�_�>wXN>��=���lվ�`A������ھ��둯�Ϫ��'��fH&�9 e�
6�����=�q־��?�=�=��`=�U�>�����-�=MК>E̓=d��>��>vn�=�=>�Ҿ���I>+�->{��=3>���>��=�菿����έ=�_!��cK�J<?Ó���~���Z�x׾�f*=�b�>\s$?g:�>���?������z��>��8=�n�ϬF�3��=��>B�
>glr>�4���L��N	��ýx+�Zn>�ܐ>��>ox�e.����C�>���}��=(Q>_#)?R)q?1�9?ҷ�=�]�>yS?>Q�f>=}k=³o>�H>�&�>$?�)>?��(?F�>Һ�=��O�-c�=�4=��,�T�<�(z����-<{�^���%=A�=d�=���= �L=���T�Q<.�<0c
?�r'?xԂ>;А>;䂾�D9�n�7�oi��Q>/�a=��>�p�>t�?���>-ɩ>uF�=|r��7����)ؾGR�>�r>�vB�����s�����>�q\>��W?<�8?L$��>u�������@�>� ?J/?��M?��>�g1�ː��� �M�ѿ#!�f��� ߺ��=S)A=�����D�s����P����������a{>�W>c�>`}ݼ%6�=��=�R�>/��>q�h��w��e�="�q=S��<iDG=?� ���=]ީ��d�=d[�p�o!���t��=�A�=[D��&.?j�->]�z�StE9���=�\�,w%���?�>?%	?n�<?��?��H���5���h�F,�e�>}rj?#�E?���T�=%yH���F��c�>�*�>�>�\��3����X�
藾 ��E��>�|)�
�����
��,d�������>U�<��"�j��?oLQ?y����}VG���J�уݾ��
�5�3=���p�4���H�;pʾJ��ʷ�Tq�={�(?�k�?���4�{�&�*�����H���]���9=�� <�u�>�;�>����������0�8��⾺\Z;�� ?��c<��D?��?�)�>�7n?Gf?�P?zPռV}>��p�{���� � -?��?�=?�>$?~<>h=��W�L��u|���)>7Š=�n�=T��<�~?>���G�>�	��<�y_�����3�=(��=s�D�MRP:�C>e�=�G?��"?�ξR���	����4=�➼��>P0��W~>R<P��%��-�>M�m>��?�Q ?��>�$޾*:�������y>Q�3?-D?��>*�"�}�t>o��Z���X�>�T�>��=�j������վ�񋾔c�>)��>�xi>kNm>;�|?
�>?j"?�q���,���u�f�,�*�޼���;7�>��>G��=�a�
�7��s�#�a�+1���o�E���
=L�=GO>�?>���=�E>��=/m��c�ؽꬓ;~�_�� �>�]�>�$?�X>��u=G7��g����I?o頾���H��D�ϾG��>��?>����?���}�溥��=�,^�>�a�?��?�c?�E����93]>@X>��>$�!<#-?��4�]���D2>:�=5Mx�9���;��;V�\>2x>W̽3�ɾq��cBB�f���JH�����Ġw���Y��~�����z4L�����s��ž*��9����:�I&ؽ���'���b��Ь���?�r�?n1�=�x�:�G	��Y�.b�9�>:�����M��������>��a����\���Ծ`D$��93�-R����>_�Q�e·�O�^��'O�?��ـ���?�����l~�C��>	/���@4$���/"��a���{?6=??qJ���1�|��\���I�>˪�>��	?3�<�뻾�>�Br?4?2�M>N`�6����J>9s�?�}�?j�R?7W��^�,!¾$ɍ��i>ID�>��>רr���N�~��X��>q`�>�d<���K��Տ�r'E����>>�?}�����>I��>�K>���=3K�<���=svȾ�׽N�>����ܘ��}+��i���g>�f�>]�%>�ބ�H����W�>g����ON���:����^5��'���*?@�����!>���> /�>ӛ0��6��֊���}���=?�w�?�`?�V2?3	�uҾAU?����=�+�>Z��>ۼ2>�� ;�:�>�W�>?ٸ�>�X�n@׾l�?��?���?sS?�o�7hͿ�ٖ�=t��5��T=�=�dQ>:"p�5l=�`�=-��<�+�  �= �>s?j>��4>�=W�8>��>����%�Tp���]f�XO��*���<��Hf�ۻ����P���x��^.ɾ:~ �������YK�����׋�p�=?�l?�_�>wXN>��=���lվ�`A������ھ��둯�Ϫ��'��fH&�9 e�
6�����=�q־��?�=�=��`=�U�>�����-�=MК>E̓=d��>��>vn�=�=>�Ҿ���I>+�->{��=3>���>��=�菿����έ=�_!��cK�J<?Ó���~���Z�x׾�f*=�b�>\s$?g:�>���?������z��>��8=�n�ϬF�3��=��>B�
>glr>�4���L��N	��ýx+�Zn>�ܐ>��>ox�e.����C�>���}��=(Q>_#)?R)q?1�9?ҷ�=�]�>yS?>Q�f>=}k=³o>�H>�&�>$?�)>?��(?F�>Һ�=��O�-c�=�4=��,�T�<�(z����-<{�^���%=A�=d�=���= �L=���T�Q<.�<0c
?�r'?xԂ>;А>;䂾�D9�n�7�oi��Q>/�a=��>�p�>t�?���>-ɩ>uF�=|r��7����)ؾGR�>�r>�vB�����s�����>�q\>��W?<�8?L$��>u�������@�>� ?J/?��M?��>�g1�ː��� �M�ѿ#!�f��� ߺ��=S)A=�����D�s����P����������a{>�W>c�>`}ݼ%6�=��=�R�>/��>q�h��w��e�="�q=S��<iDG=?� ���=]ީ��d�=d[�p�o!���t��=�A�=[D��&.?j�->]�z�StE9���=�\�,w%���?�>?%	?n�<?��?��H���5���h�F,�e�>}rj?#�E?���T�=%yH���F��c�>�*�>�>�\��3����X�
藾 ��E��>�|)�
�����
��,d�������>U�<��"�j��?oLQ?y����}VG���J�уݾ��
�5�3=���p�4���H�;pʾJ��ʷ�Tq�={�(?�k�?���4�{�&�*�����H���]���9=�� <�u�>�;�>����������0�8��⾺\Z;�� ?��c<��D?��?�)�>�7n?Gf?�P?zPռV}>��p�{���� � -?��?�=?�>$?~<>h=��W�L��u|���)>7Š=�n�=T��<�~?>���G�>�	��<�y_�����3�=(��=s�D�MRP:�C>e�=�G?��"?�ξR���	����4=�➼��>P0��W~>R<P��%��-�>M�m>��?�Q ?��>�$޾*:�������y>Q�3?-D?��>*�"�}�t>o��Z���X�>�T�>��=�j������վ�񋾔c�>)��>�xi>kNm>;�|?
�>?j"?�q���,���u�f�,�*�޼���;7�>��>G��=�a�
�7��s�#�a�+1���o�E���
=L�=GO>�?>���=�E>��=/m��c�ؽꬓ;~�_�� �>�]�>�$?�X>��u=G7��g����I?o頾���H��D�ϾG��>��?>����?���}�溥��=�,^�>�a�?��?�c?�E����93]>@X>��>$�!<#-?��4�]���D2>:�=5Mx�9���;��;V�\>2x>W̽3�ɾq��cBB�f���JH�����Ġw���Y��~�����z4L�����s��ž*��9����:�I&ؽ���'���b��Ь���?�r�?n1�=�x�:�G	��Y�.b�9�>:�����M��������>��a����\���Ծ`D$��93�-R����>_�Q�e·�O�^��'O�?��ـ���?�����l~�C��>	/���@4$���/"��a���{?6=??qJ���1�|��\���I�>˪�>��	?3�<�뻾�>�Br?4?2�M>N`�6����J>9s�?�}�?j�R?7W��^�,!¾$ɍ��i>ID�>��>רr���N�~��X��>q`�>�d<���K��Տ�r'E����>>�?}�����>I��>�K>���=3K�<���=svȾ�׽N�>����ܘ��}+��i���g>�f�>]�%>�ބ�H���r�>k���P���I��;�D0�i�;�
?�!�Cu>�i>n7>�(�ݜ������z2��sL?�?��O?�5?�1�Ml����l$�=壣>h]�>���=�r��:�>M�>�w�A$s��H�r�?]*�?�u�?ݰZ?O�j�I�˿3a������Վ��"�f<�?z�נ>Z��S>X���[��l��O�=bj�=%�>�8K>�O�>C/�>�E>r`���u%��8���,���j��-�b���Ԁ����_���G�2�I�˾�8��"���'%����GDK���3���q�H��?=�3'?��?2=�>d��=��E>�о�.���4�!�ȾEk�����#T��ɭ�z.�e��<ao�;ax��z=qF�T??�=�=�	}>+�?	��YA@>
5�=�~)>�4�>1�f>�]>I�U>H��= A>���<
H�>��+<�?�ֻ�en��e���^D���W��J/D?{��#lN�?b����Q���ս���>�>1�b��$��񳏿��>�꽘��ʿ��r�=_�?��?u��>C�ƅ����ԾU�+�߉=p�>��>���=����Ĕ���=8Λ>�5X��-�>#�>:Y:?��o? �O?��U��e�>"�>��>\>ދ�=�l�=_��>6?��A?��7?���>	��=	08�hg�<��7;F����;�<U�۽bb7�����P>��#=3�;G,>k��;W��vi=��<�Y��xg&=��?�w?fB>�=�>��侟1s�����+q[�=E� >
[$?�g4?�V�> I�>)V�=u9.��ܐ�֔����ݾܒ�>ځ�=�/���^����`��|�>���>V�k?�!2?�����.��1j��!�&>��>X�??*U�?�z�=�7���^������ӿ�	�D��D��S��O:=�ǘ��7=�X������Ӿ>���u�˽�#��p>��>�C�=ڣ>>��>��>Z3w>H,;>yY+>�� <�p������K7�������=�;���=�;>4b�<Q�L=B�ὥ~?��oa�p?��?_����}u;ꣂ�so�͝;2��>�ڵ>�W�>��>u'L>���b_Q���J�ۡ���>��_?v�?ntF����=G���� g;���>�D�>�p�=�ĽRj�*�D�1�w��R�>6�0?���>cĥ�:aM�!�X���\q>S��<G�׾gǒ?�l?�: ��J���A����ŵd���j>3�t>��6�/w��/��Q.u�m��� ��)��EF��U;?�ʠ?�8˾����5��B��0����!����Ƽ��_>�(?L��>�d��(I���Z6�
����w|���(���u���?�(?���>�i?�;?2F?F���>?kǹ�):�<�n+>L ?U?��?��>��>�Y�>�|�=��^�W�	��=Y��;�G#>hL�:�Z>
S��=>��=a�(�7����u���W7=�X=&g_:� >PM>7�6>��?$=?�gt�oS���,>���<%�>~XԽ]��<w�V���:��^�>���>(L*?�?W�e>����ph�����`>�?�h?ˬ?���<��=F��E`�4._����>L�>C*���u�� =��(k���J>���>��=I��>�'y?|s3?�h(?��f:��#���#�TuF:u�N<�6�>��>(D�=3���@>��x���j`�-���G�;��?�-�	=��>�G�=��>��=�\�= �G=`��|��'��n��<��>��>�?/Xq>�۸=4���"&
�/gQ?��
��!�&�徒�徹�=[�=@^�>�͔�|�?�, ��W\�=���רE�y2�>�o�?U�?�yF?pH���dQ�If�>�[�>��>���9���c�=�j;�9�=s��=]b��K�|����`>�h>�H�<M¾�ɾ�s=�ǎ��~�k���7���3���&�ƾ���,���r��������Ͼ�	���K���,��8�{oW��#b�R�V��X�?\c7?��=���<�?���ھ9
���=)^ܾ�8<��P��Y4�b�_�.i��T�� ����2�>�_�b`�>�鬾�ߟ��}���8��25�@�!���J?e��O������q>���<�5>mw���7���)��|�z�.{B?�$?�1ݾ����E�C>�r=�<�>/ϋ>3Nq>_L���슾�	�>Q?"��>-F=R$��Z���Z>�j�?U��?�"S?����mU��I������`?�>AÃ>�+?Ѻ���^�+>3
?T�>/��>��)��Μ��pE����>���?��~�Oܼ>���>��>H�s:x��N��?�D��<�g>��7��	G<�k� o��3���u�=F �>�q��_K�+H�>z��9�O��IF����-� �R�j<|,?�<񾢻>{&l>��>�L(�.j�������]J?�1�?�T?��7?�����������=�M�>�>���=���V�>�(�>q��q�=�3�?�q�?��?�4Y?�lm���������:����D��дμ>G�Y�m��t�<�����=�厽k�`>~1�>4!�>��'>T��=.�]>vt�a�(��ߑ��j�x�j���1�ZrD��謾s0��yݾ6��Fa�����b1��<ݛ������t�|!ʼ����\p�=��8?��
?�K�>��#>��o>EB��X��IG��P	�4�'���梗�B��[ �<�-��*�>󖾦��=̓Ǿ�7?��>�>���>f��r��>I��>�ӡ>i.�>|�=���=�W��W�:�A>�SK>)F�=�� ;��>�f�= ���E��G$2�,��|,�[5?B9��Jf�{)�e�;�ۈ��ɤ>I ?�Q>�.����6�|��>�;�/C�b��Y�;���>�x�>v�B=���a��<����Y��=pk�>��>�n;=Υo�*�?"=�$�>�W3�t�J>�强nA?$��?�s?���� 3�>���>�'>��T�R^>��>cC�>ג'?"AH?#�)?#>�>��=Xn �lݔ<���o�&�<w��^GȽl����i�&@�<52�=nq>ѺN=#t�=YR =��=�e��U֢����<�?D�!?�9c>�s>EaC�����R]�:�Q�\�U>�b=��>E5�>��?�V?�>��>_U�o���k��>�k�>�B�̋~�I2,>Qm?]��>i�?��?�>�;ܳ/��O.>1s�>�'3?tT?�G�>��->��ξtt��>�� �nܶ��[`���6���E�gX������Q�P1��K�!�,���iK��Ah�>��o>��<���=��N>t9�>�U�>��G=SnM���=��>Iu!>Լ>t�>���=�H��@���BG�R�F�7�Y�˙�c�=V)	>l-K=7l?M�
?c����#�M$���c���ﶾ'O�>?�>���>�X?��>M���P���O�e���5<�>(�h?��
?�n0�-?�=�)w=���>_�>�X">vW�l�U��t��e{|<*T�>TG?=��>�$��<�O���g�M��"��>!��8B����?q�O?ڗ�b����$(���9s(�M�<�V(>�����۾SwB���C�kƾs2��j���w�<3?1��?�оHR��J&�����W�������a�=#���;1?���>h�"�����V:���&���|�#>�x�>���K�?�?B�>��x?�v&?�PE?Ⱨ���#?��Q=1��=�ܔ��h?6�
?��(?�$�>��?.�C>�0�xG��Rp� {�=�������=.�>��'>1�4�D� >���}�=��0���>��;��=G�=٥�=�/S>�{?�/Z?�x��?����a>��>
C<G�>k�㽓?�>����@�Pq>��>5�%?5�?���>��ԾLm=��"ھ�.>|�?�_>?n��>h۴�o��>:43�7č� ���"=�<M����<�����[~�>���>��F>�vj>�B}?��@?�v!?;" �L/��w��*�{�����F���>:m�>��=Sھպ6�%s�ˎ`�E2�|46��E��'=���=��>Z�C>H'�=>5T�<�����Bֽ��;W��ʄ�>�\�>�X?�a>���=%X��,�_�I?޹�����uU��m�ɾxW߼5�>Y'?>���4?����{������;�d��>J��?w�?<[`?&%M��@�̭^>\G]>pe>��:>bF�xI��^V2�'�*>���=��y�@������:~}X>Py>����,
Ǿ��߾v�h� )���X��j%���t��������k���t(�H设C(e���򾄩f������J��{Y��n�;��6��v釾�?�(n?��>{C��v$�����ľ�Z)>�
���������5g,�-΅��Ѿ��оn�������R����C6�>(%W��5r�o	]��lP�`�ž-)��ڨO?�D���p̾@���i~�>0��>�q��,����K�����S=��^?]�??������Q���K;�ى���q>���>�>�"�甝�v
>�J?RP?�V�=m}|��q��hb*>�ޤ?D<�?�|Y?�����:x��!�����͐�t4g��Q5?���=�5��M��>M�Q?f�>�X�wSR�Am���M<��>e~?�⇽��B>���>Ѧ@>T	�=�{+=2��=����W�I<>V1�/�!��FO�p�7=���>�^�>��(>��þ����ݳ>9��&�6;���A^�����sD�>̎�\��=C�.>tv�=�|)��v��[�������)K?'1�?�SM?:?}辮��p����b<[)�>�>XB��9��='s>�ݻ>�,��:j������_?�?�^�?��^??�b��Ͽ֟��m(���Ѿ��>�->܃�>�o[�]XM>�Ͼ����<P�j����=\�q>��=>���>�W@>(��=� >����
%�>Ѥ�g;��ű7�u��,��U�����������kQ�����s��𬦽����%"��WA�J���#���t>��2?���>�x�>/ֶ>���<	�������C 6�,of�S����	����ླ�ξe���z�������ȼ5 ��?T�"=cYF���>�'���^=��j>&{��Ñ����:>e��=�,�=�6c>
�>���>���>B��=0i{>��b=#��C��!F6�?�Y����<�@?�j�nk���1���޾�f��]z�> �?�a>�"�������p��X�>�4����a�{�ݽz�!��N�>$��>e��=�ٶ<3o��4�W�A���Fu=Y5u>@3>Y�e��,���<�u�m=���>�G־���=�v>�p(?��v?j�5?�ޝ=��>I�a>.؏>�L�=��K>�O>�K�>��?��9?ه1?߈�>���=_�ۈ=m�;=	J?���V�Yѳ�9-��}#���<��4�n�G=F�s=<��]=	�@=��ͼ1��;�( =�??*�F>! :>�?+���h�_��T!��Ѿ4v���*�=7�~>�i+?z�C?/'?8�>а�=�L>���f���>��a>�.d�������=_T�=lB�>��V?|m�>n��<��=������<��P>1��>�U?R��>:���������z���N��Q2�h,>�2>k�(>���G�T>��=�!�x�?��}ݼ807>���>��m>/�=3����|>���>p��=f=��=�Dq=���=`mѽ�ϐ�7�=ҕI>k&��(�;��=��t�<��xJC���6���{9��-?g�D?��h�? �e5=� �Q◽I�>29�>_��>E?S':��<�@�p�!�i�b`%�N�>)�q?��?�ƀ��Ϗ>�bJ> >\�>&6>	H=�$O���0=�������=�>�?c�>�����Fo���
��#�>Ȥ>M�z�mx�?䆄?cH:�r���ND��`�@�վ�����������)��겾|"���;��U9�� �Ͻ���=�L?j	W?p���;c�>YG5�������$�,�ﾽ�ͽ���>��?@V?Лs>E��������ߣ���dǽ��<Otx�C�>��? ��>�Mp?�9 ?�� ?U�l�?��l=|��>:m�>3��>YX�>�+�>��R>¹>oN_��}��C������A�<�Nh�4L�=2�9>�q:>��	=c�>�[=z���ӕ���Q<^t�=M�=�Zc=���=<9�=��>?�?/F��e���%6��E1����=��!>>	谻2\��,��nL>�?[�5?:V�>[�=�!ҾB�߾Χ�B>��	?I�+?���>���<؞�=]iž��2��^�=��>^ً�(g�������'��!�Ž�ț>(B�>�:�=M�@>v��?!�.?`j?�L�=�B�1�K�3��}=�����?*Y>��Y�cc�W�I�z���j��&�5�R=څ�����<���>�h�=e�,>�E�>� >�� ������GҽƧ�9��*��[�>��>>
?�f>��
=M�ݾ2��O�A?�L�6s�G�ľ�⡾���EIC>��>$e
���?���{�Ի���+��?6��?��?�SX?b�;�Rl���>B�=�p>#'g>-��
�ֻ�ڬ�[	�>�}�QT��x)���׽��b��%6+����qM��gX��+��?̵��"��c6<Q������M���)����"��-'=�7�=�j�����1���9X���;�����Y־� ޾
$����?A�J?s��>�"�=o�g������:����=gT
��h��ۻ�~�����t�$0Ҿ�о�u����b
�1�ھ���>$�Y�$���|���(��g���>>�/?6]ƾg��x�� �h=��%>̦�< ����D����
�;CW?��9?�D�c������>L�?�,�>��%>oi���_�LǑ>4?�-?��������#��4(���Z�?���?�,F?a�о�<D�L����h�!��=Ņ�>Q!�=�������3���%?�c? ?¹ʾ��K�n<��Il?[��>χ.�(�>�4v>c��=�����P�vz��pk���-��\�=�n��Y�����}}����>�:�>)Gx���=��>��>8D꾍�N���H��������3�<�?{��/>�i>b>>��(����ω��(���L?��?>�S?�l8?tZ��8��P����~�=U�>ˬ>֯�=���lݞ>y��>[g��wr�����?�I�?T��?[Z?��m���˿I���ˁ�����=6�>P#H>��ͽ�I6>5�$=��h:��<��=�]�>��y>�|e>��9>�aT>K�>�"��:*��q��~Ñ�u�Y�y��3����ލ����m��[k��C���촾�Pӽ��x�-�u��D�3:�������"�z��?�6>ђ�>���>'Z>QtþF�����L�ՠɾ�|�V}��)�e(���ξ�ʼ��-��r����<�	)�)?���N;>hP�>�����>�?>��=��=]�$>v�>O)R>L�N>��>pB>,�5>Y�> {>N��=ӟ����1:��wP��I�;.�C?��X��˙�HS3��D߾�T����>�	?��T>$_&�Ӥ��dw��!�>�LC��f�� ǽp}&�ad�>��>��=�������v�.A꽟3�=si�>�%>%���Ǐ������=���>������)B>�T=?q?|�D?�i�>�.?ؘ�>��>]D�=�v>m�=�%Y>�U?��;?�\�>���>ԭ�=�C�*�"=�(�<��X�>�G��|��՝k=u X����=���<���<���=/=9=n=�F-=�X�<ZJ|��j==�?R��>Y �>ڙ??����
�J�`6�b������R�H�R�>��>>
/?J�;?Q�>P>��~���=叾]�0>bB�>iQ5��=_��(��;>�E�>A?�(�>���=�����G��������>��?��@?�ӝ>���<~��=���YTӿ��#��!��h��E��;|�=�YeM��q��2F.��������<{W[>�w�>Wo>¢C>*>_�2>�v�>�oF>�m�==P�=0��;�OL;WjG�G�M=���$?<�-Q�쳻R�Ǽ����(���TH��t?�ҹ���Լ��?޹J?�[V���j�5S��%�
�U��t�>���=���>���>cFŽT!�3H_���a�	�j����>�z\?��?��i�fO�=������=���>�}�>��<>����������d��>� ?��?c��>���������ɒ��*��غ>svj<��l�"�?�i,?��%�����!B�l2�ھA�S�,.o�����n�˾�+��4��?ʾ�����Da�|��>�?v�?����M>?��)g��5��ɱ���7=�w��!�{>��+>R1@��վ�d���Ѝ��[���`;�M�>�&�=���>6�q<�_�>I�g?G�>��K?I�>��2?�y�>SDU?M��>G�>��&>qj>���>(�?s沾�~��W�����S��]=��3p�=5�S>��<��役6����:��⻰y�<N��<��=HJ<9@ ���=ٖG>�2>A?r�?,��L�<����J�O���;���=�u�=.(�����Q����T>}�?J[9?4��>�jr=y����Ծ[���W�(>^�?�`?�>=�)���>�����p��$>� ,>���s�� v�R����!-�;�>�/q>�Z�=�Tv>�6�?�e?��?�9�<�/��kC�|a%��������=��>!�?>u9#�����J�����.M{���D���f��ߗ��?��-E>O�O>�8`>!�e>��>�`�=gR>���B���3�;�ڡ>�͕>�?Ԟ�>Hf =eQ��r'���B?.S��%	�򹨾�ξ�����=�ș>R���ǟ$?�	��c���J��j3-�2�>���?�P�?�V?+
��ҽ�	�>�P�=*Qƽ+��=P���!~=8?w=�!<>H�>���&O��7}㽶���l��kD�R23� ��:}ν�ÿm<m��w>e��\����$ؼ_��B�n�:~���,��}���B�����������V�+����׶�ś��{����?��\?��>���<E�L��2̾J�'���8=+��&�w`ʾ�Gi�2���%��I�E�ϔ��];T;����k=�>$����_��J��SX�XZ<2�����>�ű������5�bX=E�w>x��>Ƭ�넿����$���΃? 7?�f��� 1�,">��K>�K�>�5�>��(��3��s=7�>� _?tj?��!>�i��rʑ���� ��?���?��H?��� �[���˝��ȕ>G�T>D->�۾w]��$��E?�/t?6?�<Ⱦ\��'-�p�%?	?�'��S>���>q��>�[<��ľ�:Q>�́�V�<]��>���=�M^�9�ڽl^�~��^��>[�;>î^�S� ��*�>�о�,�\1�j�F����w�r�>�W�I�=I>~X�=��3��k���փ��C�6BO?v��?�EN?�s7?L۽�����սE���1!>ڔ�>q��=��ي>�>���o��UѾ͘!?n4�?z��?��X?��W���ͿB���2W����	����>��>�F+=����~>�}2>P�=	N4>U�>�Q�>ec�>^I>�K>E�=��=>
j���v'��������BA�<?ھC� ����U ��<Eܽ���Rƾ�I�L#�y �H�w�=�̽�]�8��o����GI=�]�>%]F>�)�>):�>����G�=�۾ :�c/ھ�r���پ�q��G�<1þ�Gz�� {�r4���(=����9+?�]�=�U�C��>�&��Ō=��= !�<�N�<��\>�j�=jo�}�=�S�<ha���m>�ys=	�n>o=���t����4�޻>���X�R�E?K-M��ݣ�Ĵ2�L�ݾ���M�}>�b?nyJ>�#�8
��qyt�b�>��6���J��E��A�x��>>�>���=0&�
3O�۸}���@��=�v>�/>�~ݼ�ɓ�M���G�=��>�XϾ���=Yx>�[,?��t?=�3?��=:��>��e>��>3��=�	Z>�-h>z�>fH?�3?�G1?[<�>P^�=��r�6}�<���<n�B��L0��>������j��X�{;s����u=�=�=]9�<���=[ =c����q�<2P=U?��9?[	�>T?:jD�5.�=�"�\B==ný?��=W�>	��>G7?���>�r�>M�D=02b������ �>4�}>��c���|�Zy >��>$c�>־O?:%?}?������b#�����=��?^�>��?�X ?G�ʼ�sþ]�����ӿS�s�V�l�Ĕ!=�;(>-H���ʾ�B�>��>�g=gs:>���<bi�>4��>q�K>�N$>�0 >�>���>Rچ>��?=vQT=hK�5�<�.�;��>y:k=�������J��v�=O��샬��I�<��v�~���қ�:(?��?K�><���
]�������V�k�>vKw>���>�d�>�?<H#���N���B�������>o0c?�O�>[�O���>d>�=	���T�>)�>rHd�ۉR<�c��O@���o�<v?[�?N�>�/U��xv��e���
+��,>�>��ɘ? �K?����]a�x)$��+�h�7�ݽ��{���@�m�⾫lb��Z��!���#�%x
����=t��>{�?�>���?�>ٜ��B��[]�2�ľ}�=u_�>0?zv�=m��"����$پ�h[��u���T>%��>��=}�>�?u�?j��?�?E1�>�O¼x9�>��>��H?O�?��0?CgH?���>��<��=�>����c�	��¾�����d��Q3>��>�~=w�g��F>�l�/�=���=��˼�;��Au�=�k�;*2=b�>r��>�?]�I?�v���=��ѻ�{��s(l>�%�>"5a�%�w�g��J"ڻ?��>�?#?�p�>')�=:o$�#45�PJ��7�>�?7J&?�5%?$��=�M/=P_�'���?@f>�-�>��=���Oأ��d����F��L�>�չ>�+>%N�>lq?��U?��<?�s��b�"�;I�����,��*C;>m��>W�>E!>����9E�q.n�����(4���"Sڽ�q-=�%-=��>P2_>�C]=���=��.>Ys��������9>Ȼ�=hw?T��>��	?�� >�'^=X�Ծ���cS?���<��~у�X;A��Z��{?>���0���(>��T��pI������W;?�\�?���?*lb?��>�̋�UF>���L�`=�ۢ=�s���i�>�ʐ�Vm:�P(>�6r���[�e�z��7�>��>ܕ�<P��flپ_K<� ��q�>�-b���&������'ѾL�&>�G�<h]��	
ݾT�B�C�3�D$,�y|T�)�I��4��:���֙�A�?DT{?��x>2>;���ƾ% ���Q">do��jA��;����Z� z��x>��̿����YI#�&��t�־ш�>��Y�dߑ�֞|��(�Ӯ���=>�a/?{Vƾ�ǵ�@����g=�$>O�<{�ﾋ�����4�I�V? �9?�W쾧���,ݽ�#>O�?t��>�X$>�*���s꽱A�>�&4?ƈ-?J�����������]@�?W��?�>?��R���>������}�?�:	?=)�>f9��!�Ҿ���)�
?��8?S{�>�W����.q����>
�X?^J���`>u�>��>f���ғ��,�q3��@}����<>=�1�9����l�o�D�c�=��>��v>�W�/:��L��>�D꾶�N�n�H���|��?�<܅?ϐ�j,>�i>?>޺(�����Ή�,�{�L?M��?V�S?�m8?9[��#��X���(q�=��>\Ǭ>���=���J�>O��>�_��tr���}�?jI�?���?NZZ?$�m��^ÿY�NL��K+���>m¤>vԚ>� ����>�ǉ�ϭ������Y�=l�>��^=&�>��>~Ja>h�w<��s�o�$�j��� S��̘1�������>jy�
M����t�����閾u�]�MP�Є/�g:c�{�޽z�r�վ�r�>?���>?�~�>�|5>ǋ�F�̾o��������B/�����㾢�)k�/^�qJ�hIپz����uݾ\��>A��<� �=W�>d���ܵ=��>I��<��A>je>k	Y>�K�>t�>�Ԅ>�U0>��k>�^�=�g�>�d�;s����h��8�]���X��^�0?�ϒ�
h$�l;��쵾������9>f�?ڠ�>� :������~N�v#�>D�
���G�����=����>�ʹ>�Կ=J���6�`��
�ҽ�	�=��>~�>����dp��	�S�\=�4�>'`־Pl�=�w>�(?�v?��5?�-�=��>]$b>���>���=��L>|sQ>��>��?��9? u1?G�>ċ�=N�_�Ȉ=�<8=Q>��]U�̱��eݼ�\&��m�<�3��WF=ʫq=k�<Bq^=BA=�>¼Wָ;��<�?�ui>���=�X�>I5���3�F����@�E�][�>��	?�o,?�c?ؕ>�`�>��>@2~�l��U�1��ƪ>�s>�,��;���>��>09�>ޫY?Q�>F�N��Gо����f>c��>l�>��'>R�>���>��6d	��FϿt�6�$��6�$��=�8=<�(�Gǭ���X��}U����<K�X>��:>�*+>#.>��7>�5>���>ҝ>)>4=,=��Z�W=�2нU�6=`����`��v��q,;;���k��fa=�!����~*�;Ҽ�<��?�m$?H�Ͻvpp��K��+��켚>�>�G�>��>䮶>�<^���#O��Z�ׂ���+ ?�Eb?h�>��o���1>�O>v~d>��S>��>��=�M���4���~��I�:�*�>�1?DH�>���w�%����#�DKK>.�<�����ן?��N?Y�Z��M��0�]�	�w��r�m�1=��=���=JU�����t �[I�쥜�7�X�ޠ�=V(?l�n?f��	��>N����R���/@�=����G�=��>%�I?;�>X빽���W�ž�S��P���8*��i"�>{c�� ?��?��>�FX?3 ?r	?��F��G?:<K��7�>�>���>S�?���>��=\�B>�DQ=�MB�|� �5銾�zZ=�yɽ���<�aE>���>��<�U,>�G�<՟�:Y�"�Ac =�(�<d%�=y|>g��="��=�>;>��?�b ?��V����ϚS���x�4	�����=�֑=.q=�e$����<_;:>m��>mNF?VZ
?\�`=��侱ލ�bؾ~0`>���>e?u�>1J;�y�=A̾g1��_#��>�߄��䐾�kǾ�ɾ�.��i��>���>V�O�@>� �?��8?�\?�q��G*���Q����!3���>��>��,>J�<�w4ھ�L�Hҁ�/@R�wC#�Ƚ٠x�y��=��,>%�>Bx>�h>~� <!�z�q�ݽ�9��k��K��*1�>��>o�?�">]C<�,þ�7��K?�+��b6�cT�?�K�$5̽&��>6�>A�L�٠�>�mD�����G���0%�2��>:\�?�?�h?�S�F��5�z>���>؁7>p�N�S��5��=_���AA>���=�ev��rͽT������� �ܽ��I�〠�DǗ�ml4�ns���jZ�d�\<��پ��u��
�S$��գ�Ǝ���Z�����j�� ]����|R���n�� o���X�����M�?�q?���>C��=�F�i��q!���<�X�����똾5S��Y�Z��ʥ���Z��a;���b��N��c�>u\Z�+,���g|���(�Z�8�>>q�.?��ƾ*�������k=��$>�ߩ<M9��p��bŚ�p��ϞW?��9?&��K�����3�>��?~j�>:~&>r����ő>�3?�\-?(D�⎿7%���_��^J�?���?;�E?�C�ʻW�&����˽���>Jl?�?a-���v����{��'�>~�??�N?iEO� �e�(L�B$�>�O?W���ͧ>�֒>b�-="�{=�+����={vٽWj�=9�>�L�(������W_��-�>%�>겆>/n� ���L��>�D꾶�N�n�H���|��?�<܅?ϐ�j,>�i>?>޺(�����Ή�,�{�L?M��?V�S?�m8?9[��#��X���(q�=��>\Ǭ>���=���J�>O��>�_��tr���}�?jI�?���?NZZ?$�m��^ÿY�NL��K+���>m¤>vԚ>� ����>�ǉ�ϭ������Y�=l�>��^=&�>��>~Ja>h�w<��s�o�$�j��� S��̘1�������>jy�
M����t�����閾u�]�MP�Є/�g:c�{�޽z�r�վ�r�>?���>?�~�>�|5>ǋ�F�̾o��������B/�����㾢�)k�/^�qJ�hIپz����uݾ\��>A��<� �=W�>d���ܵ=��>I��<��A>je>k	Y>�K�>t�>�Ԅ>�U0>��k>�^�=�g�>�d�;s����h��8�]���X��^�0?�ϒ�
h$�l;��쵾������9>f�?ڠ�>� :������~N�v#�>D�
���G�����=����>�ʹ>�Կ=J���6�`��
�ҽ�	�=��>~�>����dp��	�S�\=�4�>'`־Pl�=�w>�(?�v?��5?�-�=��>]$b>���>���=��L>|sQ>��>��?��9? u1?G�>ċ�=N�_�Ȉ=�<8=Q>��]U�̱��eݼ�\&��m�<�3��WF=ʫq=k�<Bq^=BA=�>¼Wָ;��<�?�ui>���=�X�>I5���3�F����@�E�][�>��	?�o,?�c?ؕ>�`�>��>@2~�l��U�1��ƪ>�s>�,��;���>��>09�>ޫY?Q�>F�N��Gо����f>c��>l�>��'>R�>���>��6d	��FϿt�6�$��6�$��=�8=<�(�Gǭ���X��}U����<K�X>��:>�*+>#.>��7>�5>���>ҝ>)>4=,=��Z�W=�2нU�6=`����`��v��q,;;���k��fa=�!����~*�;Ҽ�<��?�m$?H�Ͻvpp��K��+��켚>�>�G�>��>䮶>�<^���#O��Z�ׂ���+ ?�Eb?h�>��o���1>�O>v~d>��S>��>��=�M���4���~��I�:�*�>�1?DH�>���w�%����#�DKK>.�<�����ן?��N?Y�Z��M��0�]�	�w��r�m�1=��=���=JU�����t �[I�쥜�7�X�ޠ�=V(?l�n?f��	��>N����R���/@�=����G�=��>%�I?;�>X빽���W�ž�S��P���8*��i"�>{c�� ?��?��>�FX?3 ?r	?��F��G?:<K��7�>�>���>S�?���>��=\�B>�DQ=�MB�|� �5銾�zZ=�yɽ���<�aE>���>��<�U,>�G�<՟�:Y�"�Ac =�(�<d%�=y|>g��="��=�>;>��?�b ?��V����ϚS���x�4	�����=�֑=.q=�e$����<_;:>m��>mNF?VZ
?\�`=��侱ލ�bؾ~0`>���>e?u�>1J;�y�=A̾g1��_#��>�߄��䐾�kǾ�ɾ�.��i��>���>V�O�@>� �?��8?�\?�q��G*���Q����!3���>��>��,>J�<�w4ھ�L�Hҁ�/@R�wC#�Ƚ٠x�y��=��,>%�>Bx>�h>~� <!�z�q�ݽ�9��k��K��*1�>��>o�?�">]C<�,þ�7��K?�+��b6�cT�?�K�$5̽&��>6�>A�L�٠�>�mD�����G���0%�2��>:\�?�?�h?�S�F��5�z>���>؁7>p�N�S��5��=_���AA>���=�ev��rͽT������� �ܽ��I�〠�DǗ�ml4�ns���jZ�d�\<��پ��u��
�S$��գ�Ǝ���Z�����j�� ]����|R���n�� o���X�����M�?�q?���>C��=�F�i��q!���<�X�����똾5S��Y�Z��ʥ���Z��a;���b��N��c�>u\Z�+,���g|���(�Z�8�>>q�.?��ƾ*�������k=��$>�ߩ<M9��p��bŚ�p��ϞW?��9?&��K�����3�>��?~j�>:~&>r����ő>�3?�\-?(D�⎿7%���_��^J�?���?;�E?�C�ʻW�&����˽���>Jl?�?a-���v����{��'�>~�??�N?iEO� �e�(L�B$�>�O?W���ͧ>�֒>b�-="�{=�+����={vٽWj�=9�>�L�(������W_��-�>%�>겆>/n� �����>���H�e��sz��J��[���Z ���>�����=`�>q��>�k*��b��H=��H�;�?�F�?�l?k�?����M�\��<���>0��>L��>f��/d��n.�>���>3��;�G�;���6�5?#J�?C �?�S�?�+R�<Gӿ����������=,%�=��>>��޽�ɭ=��K=�˘��Y=�e�>~��>o>C;x>u�T>ћ<>��.>p�����#��ʤ�2ْ� \B�� ��� wg��{	��y�����ȴ���E�������HГ�w�G�`���T>��V	��x��P?_E�>k��>4�>&�5>}1�� ����> m-��u�8ƾ�f�,�_��xbY�Ԡ��.���g="xJ��<
?v�fT>���>jR�=�|>��>�}�>��>��F>�"5���u=�R9>GG7>�}U>�>��=m~>?T�=�턿o����:���N�/�H<}GD?\�
���ot3��߾Q/���[�>&t	?��S>�#'�����yx����>�b@�2�b�e�ɽ��"�0�>��>	i�=���U ��Ew��j����=>_>1�#��O��0>�B�=ۑ�>�D��'>�>��*?�x?A�0?�M!= 5�>~�>Ce^>���=ֳ%>��E>Ww�>�?9m3?t&.?���>>^�=run��=�<��\=�u�����ؽ1%l��X��{�<�=m�<��=uo�=.!�<VɄ=�K�<ݣܼM���4�<ʶ�>A�5?�c�>5Z�>H�[���I�d�L�F ���(>S�����>X��>���>A��>h�> ��=̧��:޿�`XӾ;��>�nI>+�f��Z�)���{>~�s>��V?��2?D]���+R�L��; �=��>h��>�y#?rƪ>6>4=�;�	�L�ҿ|�"I.�h���j�=� 7խ���{�=�k)=�V��i�C��=��C>��L>��}>�<>��+>��8>��>�cl>���=�<>�	�=;�<�������� ��"=�(L���[Ӧ��{����􊽃�Z��T���xݼ��?�.?@Ȅ���]=��=��[
 ��??���>P)>��?GƽmI���4��|�J=%?�Tj?H'?���@?]<!������W>n>� �>��>,p=p/(��+���(=���>F�??���>b�F�]$G��@|�:�E��>Gn�9E�����?޽s?a�G��\���6"�f�K�4P���K~>����,>拹�����nN)�&��@H��R I�Ȓ'?dO�?�������F�0_���l���<B�>X7�UaK?��U>Zj�������JB�Ѝ��D����L=S��>��L=���>�n?��?&�R?�?�?a���H�>�ց<4x�>��>@?��?�}?b�>��h>曈�v㦽��,�����ⲟ;�z���=��!>fz>�)u���=�=jK=-�V<�b#��v<媢<��==���=H�>C">D	?�T?Q�-�֚B�Fj��`˺�	X>;v�>I�b�UC����L�e�N�D/�>ӬJ?�He?��?e�}=ϝ3���>���R�YI>�a?�-?��>&9�<\�j�*����<��E>#=R����Ҿ)�ξ�i:�s�4>ܳC>0��=g>��~?�wB?8"?�^��D�.�-Rw��q+�� ��#�K�ރ�>Z�>��=�۾j�6��Os�8�`�ڂ1�i<�q�F���<؉�=sj>��@>J�=�c>��=̼����ٽ5c9< ����2�>��>-?l\>���=�F��5&��1L?Ο����+�>�~�N�^����@*��#�>pY�=���>%xr�\�r�����m8�B��>9�?��?d�?����������,>q;�>��>l���a|��]7�ݙ`<zz�=�;��}��Ծ�����>�B�>Q<����\뷾�b���uÿ3lP��{���Xw��9��K�6����޾�"��r�=Yj�bCξ2,��De�D�A�vH?�R,��O0�����A��?��}?�k�>�bM>=����e�ؾ(�p�DS��rὒ����梻!�,�9�����`�����8 ���4��-��>��������}���.�w,I�g�=�/?lM��q#��=Gɾ��=߯=n;��������AZ����ƽ��^?83?�)Ծ���k咾��>��?�N�>G�C>�EA�U?(���>��(?�P2?�����w���vi������?�o�?0�J?�����6�A�/��`�]�?Ҽd?�?đW�/� �	ܜ���?�fP?�(?��d����9� ��"�>4J?F����>��>��r>*s���2����=&�nY�=��=���<���m�ԃG=���>�s�>�Eh>�Ҿ�����?��׾d�Q�x�o�jᅾ��"�`�ӽ�?�	q����>|��>���>_�b�,�������z۽ �&?۷�?
jb?�F!?�|����'�==�H��>��> �=I�=܅���O�=F>q�վ��P�����]�>���?ѱ�?�0?k�B��п9E��\�ؾ��ʾ�:=Q�>�z4>�~���.�>�'�;D�~��>d�	>�q�>���>���>2C>�D�<r.>�<��U+������0��b�e��;���s����^þ�����7��D�^ݾ 1#����.�Z���0���o(�]�	��g����H?��?�S�>n�>�5p�C���"^���d��i,�쭼���;ž��;`؟�J��:��|O3���>�IپP�?*w;�)�<�s?Ky�iV�>z5�>�o><Fr>B���釒��L	��[>�3>8-�>���>+�?=o�>ܑ=���ʭ��fP9�ƉP��i=�dF?NEe�Hn���O3���䙜����>�j
?i�D>*'��앿/y����>��Ҽ��`�t��kf:��C|>��>���=�ϱ�H[�:6p�d���=o�>y�>��<��~��>(��"�<M-�>�rѾl��=�x>�r'?|�t?86?�=W&�>��b>���>�M�=�RL>+4P>�݈>�?��9?��0?j��>�I�=I`��~=�JB=[�=��I�����A��U����< �?�cC=`e=�4�;/�T=�I;=n˼ S�;�E�<�?�>p�7?׾�>o��>T��OA�.!K�oP���'><;�����>���>'�?m��>�.�>�� >&&������3ھkS�>5�>>�.d�H-x��_�ׇ^>,�x>��P?8�0?m��}�^�t�=\��=E�>�9�>!*?�j�>k� >�͔�z��8yԿ�z4�Z�0��h��A�=ȥ�<����ƱC=�na��� ��a7�R;]�V>��>B�>tM>>Z�=:�*>�@�>��=>�@R=?4�=①<���<�S��V�=JĽzU��y�d�J�#C���������̽�b���cv��*�
H3?�H�>�w��=��=�%߾L�*�??��>���>8�?S����e��3���'��{ ?n�?L%?a���`�=����r����>QU�>j��>���ի���⪾"!��83�>�3c?���>g�`��J�/W�����D��>ӻ<�����β?rTZ?��S��Ἴ,�,�2P3����먜>,�X=�8��7ܾ�.�<. �Q]&���꾩�E�6~�=^	)?��?|��fJ��}�����6�)�(��<G$�>�E&>s�%?��e>�����pA�3���R���)�>C�?����0?>��>���>u�>-�_>�~6?䛅���?޷�>/��>��8�G��>yF�>��>��?�$�>k��=��<1����`�.�=δJ��q	=r�;��>�u�,Ӵ><�{>Ԉ�=��<�UI�[�q�c{K�E헼?�~=D�=�eO='A?�e?W���,j����z���սp��=.�T>}R����D���n���f?>#e?�$I?��>��|=[r�������Q6z>Y��>%a?��>;�=�-���������]O���Ȇ=6x�>���d�� ��)��=��y>M��>�g�>fg>�~?�yB?�="?�}����.��Mw�Vu+�ʗ���XK�Wh�>r�>��=�a۾'�6��@s��`��1��=��G�Ë�<���=��>��@>�P�=�V>� =O꛽�`ڽy8<X��!@�>]��>�1?e\>X��=�<�� �!T?�y��i����U��NM�sy9�g���՞�>���I�?zƊ=�c��ت�|KL��ee>?Գ?$��?��?��ڽ�j�@�>(6|>��>*D8���缤 ����y�;>���<#p�-Ӿxc�=H��>x��>e��ZJ��.⨾V.y�k�¿��]�/�v��w{��.��5�`��>��@a˾z�3��̾V��=�^=����6&���kU�wž�*�
�����ɸ�?=ȁ?���>��Y>��ؾB��B��2>�h#�-��w^��L�P��4ڽ)0���s��q���6�j��K��^�>�"V���j:����Aa9<e�j>or0?	��C��-	�ҿ)=C�i>lDv��x���r���Ԝ���h?�s/?q�ݾC��!��ef�=��?��?�{+>����U=#��b�>�B?�,=?x��=�����y����#��z�??��?�b^?��.��9�R�F�P:����>�\?�*$?���� �n*ݽ[�D>�:`?�"?׺��_ئ�:?W���>\?�n/��D�>Y�>��>�����5��,:c<Q�5�=H><��5�[sW��[�>�R�>��>ш�>��#�m�@�5(?֚�+Hm�/@����_�NZ��EG�[3+?����W�>�C�>S	�>5�L�囿�����ּNv?�~�?ݧn?S�?���E���k�l�>��+?!8>��6=�[��xF�<���>� ��,E��.�3%@?m��?m��?4��?��q��&ο���jJ���B����>bD�=y->p(�Q#1>�N>�񉼮EI�/��=<��>�ʃ>p�>�\>�q >�>����T�,�����#���3E�	�����j��i����=�b$	� o���ʾ��ƽW��+&H��q/���.�Ҹ��g��O��|�W?�4?a�μ���>�)㼯�<�'�>�����UF��EY�a���e!��\��侾r�Ӿ�&�N�=��)��>͜R��P>ZL�>.t����>�>�P>�iP>�0)>��=��(>�?�=&>�>Ju>���=>|>���=��� 倿�$:���O���;��C?V�^�f��A�3�R߾�2��l�>��?y�S>�f'������x�O��>k�C�ozb��9˽� �h�>��>}Ż=��ӻ����cx�5��}��=U�>�/>�L����p���=���>�̾�(�=��s>�~&?+�t?��5?���=�ȼ>PP>%��>к=I�R>��S>���>�?�9?�<.?Ώ�>���=T�j���=��D=�3��?i�����?ÿ���ڼB��<�g �k��<��>=8�ڻ�h=S�<v�ۼ:j::��<:�>�8?���>�u�>�]:�(�>��M����z�>"+��B�>�^�>ܼ?�P�>:0�>E�4>U�a�`þS���>��@>S{_��x���dTw>�es>\�O?˧1?j�j��"c��{�<�>�=��>\P?BV)?{A�>�>�$������lӿ_$�P�!�����w��W�;Y�<���M�A�8Ϧ-�������<{\>��>��p>� E>��>r+3>�W�>DZG>F��=�=��;l^;kF��qM=�]���F<��P�����gƼ����_����I�,�>�_�ޞټ-�-?�r�>�g����a�+���W諾�r��q�?�Ɓ>m5�>��?d�i�3t��,H�gW?��k�|+?H�h?�/?�m������·�+k�1�">ĭ�>��?�g�������;��e��>su?7��>��=�睄���y�8�/��L�>��5<,_��IA�?Xn?�_����t�@�� D�q�⾺��>MO۽�0�=@
��������"�� ��ᔾ�\ؼ�0?/��?�`�eɽ���@����&F���*>�Z�>��>.�R?���>g�Ⱦo摾��G�3�D��[�g>��!?���RM?���>�f�>8�^?ʴ�>H�1?��{��?�[�����=���K�?��>���>x�>�=>r��QY��qE�c�Q�m��=����w�=�V
;L�=��9���Q>DP>�ǿ=Z�<�ʽ~$n�o��=�
0=Z�0=�N�=��t<'!�>wZt?��I��	@��V���>���=�>E>r�5��S��Ա��`�ƽ���>,�Q?	\?�?S�Z;����֮�u�)���=CK�>��?�͇>��Իc2߽���fG�=�ݽ��^�=��;�8���@ܾ�q��V�>���>�&Z>��f>�~?�aB?�0"?7��� �.�-w��\+�K���qQ�f5�>���>���=oI۾��6��/s�t�`���1�u<�T(G��*�<D��=+>L�@>^�=�p>�m=2�����ٽ_9<g����>Ů�>V?PH\>�:�=0]��d�"�[?� ��Ȯ4�uG��H���P���~�>�>�_���0�=^K�>�nS�UԹ�E1Q��c=>�n�?���?�K�?�􄽌�5�eA`>�2>�o�>�ӽ_GS���י���Ѝ���K��E��*�fJx<�R�>|�6>�6޽2·�a�
��롼��ſhc��n�=%���ھ1���¾�Ѿ�BR�>2�=�R��J�,�5�J�s�����G�����9�Ӿ���{;�?=��?�w�>�4�>�3@�v�ž|��#\Խ�b��LN�f�ھL�P�}�{�!����O�2���z<�{4��_y�>B�]�ڂ�.�x���;�فȾ�l�=̦@?'OA���ҽz�y��\s>��ü'qQ;�e9��^��@&��?M�-w?2�@?Ԭɾ�[A����u&�>��?�m�>!�>3ҍ�3N*>?��?ǹ�<�՗���f��^B����?3�?�R[?2�$� W@�<x.�-\Ͻ�_?�d?��??��3a��(�<4�>S"]?F ?s�+��� #��r�>�_?ЂQ����>�i�>yo�>$�9���{��yY^���4>�ł>)V�[\X�1�!����=�Q�>ű�>�I�W㾇���X?oJþ��S���[�	�,��7��W���3?,>�+>6Q?�I�=�R��ͦ�����?�5��!?�j�?�i?�V.?ZF;Ԥ(��������>��?��>��e> <B=��>��>�=����$�w["�Ȗ.?\��?�|�?!��?�I?�o�ο�l��7q��>��9->{�C=�ҁ>F:b����=)܈�I���Y��(�=��>��z>�"�>'F>i1>X/>�����&��{���k��rV�"� ���*�|,ؾ�0�I��/�9�A�׾�;�?W��� ��ՠ�6�Y����#����!��!��cO?i�?:
<���>ކ,��+�����=gvƾ�|������i��{��]��,�d��]������c��=�{)����>�25�-�i>U�?� >�ݟ>uW�>�:�=��^>�<>� �=��>��� @�=}�C<1�H>.�>���>��=���ai���A�iL��r=vB?�+v�����4p;��`��vd�����>E;?!�+>��2������4���з>��`=8/F�����[����e>��>��=��nc�=hA�����k��=�<�>�"6>�Ե=�d7��rN��h�����>�ܾ]��=�ti>��'?Y�u?��4?�f�=9g�>��e>R�>��=Q�H>y"?>#��>
?�9?v;4?�'�>N1�=��a�PO=8�C=��>�#b[���������>�{��<Y�?�n�@=��f=+D�<|e=��0=��U�6<T�<�*�>��8?���>�5�>I<��9?�,M�b��f>�}�m��>i��>\V?qc�> �>�3>qd�LþT�㾂��>�SA>��_�egx��-�Bw>A�s>E�O?tM2?�xj���a�y��<g�=�:�>_?�s)?T��>h�>?ȥ�?���ӿ�[!��v �C�y�8�м�o�;��<���O�%8�:��0����<�g_>�>�Ym>��A>8>��/>���>�E>���=�U�=.C�;/A:�HI��>=� ��Pr<=a�nݺ�Ҽ�����C��3�G�f<��
����-?j@�>萾�þx�B�����H/���"?)? ��><(?�&�=
��[���:��h>�(?�??��ƽ���=k����	��>���>�p�>&f��_>[���Ծ������>(�l?T�
>� �=�_�d��w�z��>�@<�����t�?�fc?C:����:U���U�g����>A�(�n�����jJ����F�vq"�8 �������t<o�0?��?A�/��u�̲$�2���a�U�il?�B�A>��<У4?;�=�J��n��y*S�T����h��7>�>?[�D�CP?�a�>�D?yil?ʽ?��>�L}�(�<=y�o� �?>�9�>�>/�.?�F?��>���=ZU���='k���ƾ8��=�� ���7>��=Y$�>;�4=��i>c�2<��½ɪ<���{7u�>Z���<gZM=�>^�=X�?�a[?޵���*=<�<O���<ؔ>Vl�
�>V1����.>�[>��1?��R?���>럛����}2�z��uZ�>K�??��m?�e->�A�=��[�D1��T6���g=i�>�^�>f}m�PV��\���R�m�>^ݩ>OU�>a�f>��~?TxB?�B"?}*����.��Ow�1x+�~��,�J�1p�>�!�>)\�=iw۾�6�Ds���`�ӆ1��<�,G�S�<
�=٩>7�@>g0�=�c>��=B�����ٽ%�;<����u,�>*��>9?�d\>x��=�N��%�L$X?�岾��+�MW���꠾��$��F;=���>��l>G�?��>��D�i⧿tKZ�F:�=�c�?��?�r�?)�����0�.>�E|>Nf	>�R��<��+����|�(9>as>��	���s��V����>�~�=�x�0�g���ݾ��Q�����5�\��Qw>��2�옣�|놾�|۾V��X4��^g���5��ˮ��*���1��ʏ�6@��č��������?oX?�k>H%r>V@��N���2�d4��}s��Ŷ>� ~���<��B0��V���I0��3���,�]��u�>��Y�r��!z�r	.���+�ߪ2>�l-?��¾ w���(�d��=aD>I�*<Z���酌�О����?�X?t�;?�㾥�N����>?z��>e�@>�̅��k���Ś>j�/?*?��0�_W��x���/ o�2�?S�?�rV?Fe���`�`�=����=�?��o?�X�>�=q�|�Y��)n��?y�f?׾b>e��%����A��2�>�Z?����|�>�
�>�[�>.=2<�7̾��Z��D]�|���r�=�����*پ����3؃>XH�>�J#>	�^�M��'�'��?e8��'n:�/A��r4�u!��V�K�.?�5�=�P�>-�4?`VǼ�S�7���d���_8��E.?�=�?YFb?��1?���E��Y[�L��>�.�>�P�>�5/>e�8>��=$��>�|+<����J��>t5�?���?ߨM?��)���׿24��@禾�������=D��<boe>>9����=N�=��a�%&>{��>�c�>ʟj>T>K�B>�>MS��\w"�l皿F׊�s�J���"�����m�9�mE�����<��ʒ��E.f���Ľ�����G���
�C݌�����(��Z?��9?մ�>��>��.�M����XJ%=�&������v��*X�D7�b��0����þT8���=2D-��1�>vϽ>T>�H�>����d�>iF0>1V>3�>pZ�=�(�<m++>�o&>�N�=��P>Ǥv>�״��v>�ό=�1��1E���&:��0M�g�R<��C?7^�"k���3�����M��\��>
?�+Q>�'�FԔ��Ix��N�>��%�O�a���Ľ����>�c�>ni�=��M��o��F�t�/���g�=
Y�>ْ	>�P��쌾��S �=��>R�оo�<U�0>\�&?�7i?^)?^$�=s��>8�u>_��>�m�=P>�׽=��S>p?U :?�NA?Ș?]��=�Mn���^=� =��$�u��j�ǽ��k�Ľ~�%�����a�<��U=`��=c��=c$==�4�<�Z,=`;b'�>ߵ8?f��>�`�>�;�f?�MM�:"�v<>����>��>Of?��>	��>�4>)�c�7�¾V��ǘ�>�RA>>�_��*x��+��v>��s>��O?u52?��g��Ta����<0�=���>�7?�)?	��>=g>�F��5��OKԿ���Jn��̖����	04=m�c�nxT��,<�H�{� �&}4=�w>�$�>.r>��A>̃%>��>Z;�>�cW>�5�=9��=�})��w�%����ɖ9+�(��Y�!���gW�Զ�H��aiO�s<��Ykm��8�P1?G-�>�V��a���?Y=둅���m��-�>��%?QL�>ll�>a��>����n��=�� ��?�ń?�)#?�K�l��=�Mʽ/�4�1��>�-?fY	?�����犾�����2�i�,?)?p?l��>�����m��b�������>�
<=2��?]�?��^?�M����odR�(F���
���>J�j	I�Л۾���"���A��!���7�ψO��iD?���?�����`���8�����K�]����;ź�>�f�=��C?�	>vƛ�H��l�^����kБ���h>�+?��C?ɋ�>��>�^?���>�?��5���>[�=��{d>C7{>:U(?�#?a��>R*�>��=P�f��j�=��o�ƾ��=�+=&}>�5��PTp>vhX=�v>3��=Y2b>V3_<E���"p=j��<�/��;�;�Ü=�ڍ=�-?<�q?�y����Z8��ӗ<��4>˫�>�G���:G�.���l�v�`�>/�@?��G?��
?8b >�\	��w��5�D��~>��?
o"?ك�>�Θ<��8�ʛ��P�<�Y�=~i�=�SO��xӾ_P��{N�=�$�>���>��L>��f>�~?��B?RK"?�>����.�qQw�V�+�&䤼�nJ��V�>G�>�;�=B�۾z�6��Hs���`�ɋ1���=�\�F����<^�=̜>+�@>*8�=!N>�e=�$���dٽXE8<􎕼�'�>���>n2?�g\>x��= U���6��X? t��7@*��ξ�z�G�ܽ J�8k�>s�'>L��>��(>K�i�]U����Z�G��=���?Ȑ�?qY�?,[��N����=(�P>�#>���=����e�䀻J>�b=�Ҫ�L��Vݽ}��>B��>�ז�'nr�%W�����fp��+�]�3��=f���݂�Z���G#���Wؾqi��+;����hZ�fs(��d��g��<^h{�6����¾��꾟��?�َ?=��>��>|}�Bپ(&�%��������Z�����ٽ����������Ej��<2���:��
���>^Y��*��f�|�K�(�e/��r�?>m"/?��ž�z���A��q=�0%>��<4��b�������f!
�a�W?�9?��,O����ὅ�>'�?��>[$&>�ؓ�Q𽢞�>,4?U�-?��U���'��q����?R��?�(U?4��_U��`=�Κ��T?Ed?{�><�+OI��i%��?�#d?6{�>���1,��j� �yG�>��[?^�t��"g> ��>}�>Kƭ�`�پ7��ı����t��=����_L�(z>�t�>���>���>5��=T:�z��T��>DϾD�3�8I4����C�4�t�A�c��>(�X^�����=�[x=H�4����믅�����p\?+[�?�2K?��1?.Aq�,p����R6>�Ӵ>�3!>* *��{�����>@��>�9��z����?���?ǥ�?cvK?R�k�O�пQ���q羖���B/>ǣ�=�J�=�e<���Z=�n=�>3��+0�ˈ>���>0�H>�F>5 A>z�>���>z���6������X��X�I��i��������N羁3���i=�������ᰈ�8M������8��}0=�b��9���&!?���> ��>���>ꬸ>�I�󅜾�Ѵ���ﾫ�ξ0���Y�����ྚ���񈻾���� ��;�=��^L�>���=�:��^x?�u>d�>��k>���,��+>�F
��ޑ���u=$��=�*>3��>[͟>���>��=)�|�ȗ����E��1\�`��<N�9?fr:�,;���u!�$�ľz/�����>M�>l0,>�v,��$������u̼>�W��e_d�I���	_ּ9��> �>��7>{����D��MP�����9/->�"�>�^>j��;�M��Ϯ��=L��>j�־���=�Ё>�O)?�~t?�r4?��=�a�>p#a>.�>z��=v�V>�2T>Ls�>A�?�6?�0?tn�>Q'�=��`��Y�<�E=�>�U�?��5��;n��Tc��֕<Z�>�Q�>=�*_=��;�g=j.E=xa¼��;���<>��>�=?7�>�U�>�Rv���=�܎C��K��`*>h%��@�>NA�>5�?��>���>VM>�!Ͻ|�����P�>22 >!9\��4q�"���Mт>�h�>�"U?��(?�K��:�N�4�X=]�>��>N?��'?2��>y0>��Խ���d��U�K�P5	��9<_\��^�/��j���
K;�HX>V��W�����>dR�>��H>LB�=�ں=;�>Y_|>,U�>�@�>Y>�M�=�=�$�pU�]qi:*��:_�=�./>�f���͖������@&�s{ƽǽ9��L��t�?~�2?#kU�aZ������W���&>� f>B�>Ǔ>����Ǎ��Al��[�ނ��=��>cZv?��>�Ge�N�<4�>�*>y-�<F��H`>��1�����Y &�w�>��>�D1?�'�>q�=�����W5��"J1�I��>E��=dͰ�O��?8�m?�!M��hK�8R��a.�q#9��¤��ȾmѾ�Jپ�Z0�ŃO��U�^��.�rM�=�K?Y��?f̽���<t��B���>��W�;P���Wl���>��߼�8�N�������7�rv	>�P>/�>���>����V=?��F?x!R?ru/>�a>f޾>�@7?*�F>K�>A@?�;?��?P�y>�0��<yD={�$>;G�>��;��^��ڃ�h��=>M�>5>F�<`h<��=��.�),��雼�@=���=z�-=Ei�;�3�=��>�$?C�#?����7������x�;;> �>b�>�=;V=�S>!��>��>L��>I��>��<��������\��k�s�?Y�??�l?�Ӊ��_�<)�'�'
�]k�=.q>�=���þkb��g���A��>��>���>��>�?k�5?���>���F_R��<W��(�����>�3�>`dx>=6&����E�|�w�ߋ�k�y��ؗ�`����C=���=:9�6�VCM>� >U��=�"k>���Jj�=I�>Ur�>ܷ�>���>�;�>�ʇ=�����3��:M?���>a�H`�]98��G�>���@}���3��+~>Y=H���k�ƿ%I���m?���?K�?��?-'��j�2����>31�Я�uHm>�8�0�Z��!d��#�>�3�>��<ч��|��=g�=5!�=�r:�W���e�@��������Q��y۽����o���k���s�
�ʷR��ڽs���:p���1���6��`<���A�ǁ���ZԾ�f���?(�D?*�>�r�<�=�8�¾��Z�ə2��!Ҿv����վ�l��K鐾⪾�����쾿7"�9�2�ޟ��>g=Y�*��Z�|���(�(r����?>�3/?�,ƾڬ���y�_�h=<�%>�3�<�=�<���m������^W?��9?�f�B����T���>�?Os�>#M&>o(��"� �>�-4?,�-?������%��Y>��zi�?���? �??�[M���@������@?/�?�{�>~%����˾P��0<?��9?���>�(��@����ĭ�>qZ?��N��G`>��>��>�콺䓾��&�����j�v-:>2��{2�D	g���=�=�=��>��x>��Z��߬����>lGݾ��=�t�6�+z��/�窽���><����n�=}%�=�/�S���^���P���$RW?���?�oB?��.?�Ǡ�����CU�>��=��>r�<>��N<�uY��A�>���>'� ��������d#?�$�?��?gEG?~�q���ڿ{���ľ����Cz�=��=��;>v4�����=<ڒ=��3�i�Ļ]*)>�,�>:.l>5�h>�OK>��\>��f>��kN�����ǡ��$\6�2�
���
����y��'����!����匩��5���I��T�@/��S�<�1Ծ���=�?;R�>%}�>�h�>�q�>��>��w���� ���������E쾦M��s�v7����J�]�`�����ۅ=ϐ�ǐ�>{q�<�>�;!?��M����=��>��"=Թ�=gka>6b�=GJ>��>��>�!>��C>��l;�܁>5��=̊��EP����8��N��̅��6<?
�g�e͑��&0��辽����b�>U?��q>��!�#J��#~u��x�>1%?��ob�&�޽�OF�\��>R��>#��=e�s�Dd���V�b�佲��=>d�>g?��6�����VZ�=���>��־��=:�{>�*?��u?�#6?+��=���>ɕe>k^�>���=r�S>��W>B��>2I?g�8?t=1?a��>Q��=c`����<�6=��<�eeY�|!���/������;�<����OF=�z=���;�W=q�4=��ڼ���:���<�>��:?S�>�Z�>�J�jr?�H�C�N��8>�̺���>j��>�y?�u�>wd�>�=)>~���c�ݾZt��>��/>B�Y���x���Ի>�z>S�x>�X?�/?���9��B=��>�ޯ>b}?�,?�t�>�P2>J�����
�NͿ���Y����k�=޵�&`C=S�$�!�j=d�@�����bǽ�:D>���>⼋>Y�9>��>�kk>��>R�>��,>M�K=��=�dT=�2=�*���=wBF����Qg^�/�Խ����3�r`��G׆�mwu���7��2��N?M�.?�v��n�J����	����z��>�`�>�d�>���>�V�=I<��v�}�?��[]�� ?j�?��>ꏊ�f��<Q�K>��<>�%g>�h>���=o�Z���W�޽->�=
��>��K?��>�]��b	������"�2�w)2>�>/6ǾdĦ?2�x?`@���3��yɾa=�5�E������8�Џ��A��t�:��(c����u�:���)=9=
?-L�?�Ͼ�Yy<�s�9��4Ȗ��꾲�|�8J���i>����޾
�Ⱦ�z޾�����_+>oI>֣>��> �=��?c~ ?�	l?rm�=P�?x1�>f%?���>�?�8?�7G?�&??�A�>�73�vFf�id>Y�D>$>��1���l'=�1>{�>{>/>�x�<�A�=���=.j��~½)�<���G=V<r��S=�>eH>�	?�$?��ɽy����[���L��PQ=IU">��L>��<gg׽^W�=f�>`��>d: ?�H�>J��;%5�Q$�r�ZJ=�*?
�+?j��>���<��=C2���\R�`�<E�->�Ҽ�G�BZ¾,��%g��XP�>���>ԳA>�D�>�4s?XC?�i�>�ɑ�LHJ�Q2�f;�to\���^>��?�c�>���=c�پ�t.�i�/�z��h�s���7���I`���:>�ұ:u�=}շ=�u>y>O��=�ރ<Hܜ=\u>G�>��>�%�>N6~>N';!qܾq���8G?6#o>�e^��1C�ʰ����>q���&������r<�=���K��7������J?r3�?f��?�l?Rӯ�v��ǘ>�5��(Խ��Q>��L���= A>�>�>Bti>�->֧.��ѼȨ=�>N�Ig�d��c�h=�Ԯ��`�o����Y�U?��4O=.z��~N�<}�a��gȽLm��o�r��tW��O��{����z
��M�ݾ$�辗X�?�#?3��>S�=ya�ڴ޾�:���]c<�@ɾ�'s�f쾳���C�����Ⱦ����$���<I𾹼�>y�Y�}7��%�|���(����r�?>�0/?�Vƾ&Դ������g=�[%>.�<�Aﾽ�������*��SW?%�9?�b쾽��:�ོ�>��?�p�>p�%>�D������	�>�14?��-?��[���7���+��)i�?� �?��??�O�xA����ߗ���?R�?���>xÊ��`̾����.?^�9?܈�>�r[��	A�!��>vg[?��N���a>6�>�g�>!񽁐����"��"���Å��a:>W��@����g�*=��ڧ=?��>�Xw>T�]�����><ɠ���/� %F�4L�2�J��
d�n�>�P���y`��޽�i&=@�=��������i<�<��p?�!�? 5?m�/?gc~��Q���ݾ��>v��>�D#>z�Že\�;@ե>>�>b��t������k?���?�?��F?{k���Կa������iÌ�h�M>=X`>��C��E=ѡ��9s�xv�<�p9>��>|T>z>>�>O2�>He>8Ã�l"�
���⋿��m���x���!������F�����޾�bHȾ�h����U��_�M��(2�]`��,��K��>��>�$�>j�x>c�>���v�ʾ�Ki�,�ھM�
�u9¾+���`־7Z���nf���N�*�޾�=�n����>Ͻ��<d+?->�ģ>���>��%=h��=�~�<�+���=��8>z/�>�̦=�́>�k�>|>���=)4��x���:��
P��0�;^C?[g]�ޘ���3��ྺ�����>��?2�T>9K'�<�����x�;��>�WH�[c���ɽ��<�>E��>Ը�=�_ػ͒���w�[�� �=��>�1>^j�@���Э���=U��>;�ؾ�w�=䗌>-<0?;�j?R�7?�'>���>KAO>=��>M�>�x{>t�r>"{>wU?1?h�-?���>]�=rR�k�F9���<6� �Wì����@������Z<�Eu����=�X�=��<��Z=�
�=�l����*<+�=�d�>�;9? ��>�s�>��4��B���K���%�>0��G��>'z�>E�?=X�>��>#(>%2����˾=4��[��>�a!>P�W���o�u�����y>*=�>��Q?�5?,D��9�e�sĞ=�r�=t'�>v�?*+?���>!�4>-^�����oLӿ�#��$!�}�{��m��4l;�P<��%N��Ǒ��.�+����r�<��\>QM�>I�n>>6C>��>�80>2��>YH>3��=ٶ�=��T;,�;�J��YF=�����E<y�K��琻ޚʼª���̍���M�1�@�yb��� ���?G+?"'�Rc�>o����n>H�e��=��=H�>ypq>^!�� ��\xv��^X�t�P���>,<j?@&?>^A�r�#=+>�g�='�>e�+>��;=�R=�%�i��!Ti=i,?��-?��>1���e���ᆎ�Յ��PI>�i=��r��қ?�.;?�� �)f��9��37�� �+r:�05y�=A����.T+���S�Y ��+��hٽ�'>�� ?!��?1�M����p꾐���m���w�Uv�� ���<��>�%>@(����Ѿ<O%��׃�;�<�x>��C>�`>�����>8�2?��X?��J=�?���>$1D?�.�>!�?��5?�J3?ܘ?xx>J1�:�{�E�D��4.>�5�*l���*�1�B>�g/>�">�S>���=S�k=汎����������I=8�2=gg�<��;"� =��>(��>J<?t�#?$�ؽ��a��� �T�����<�3�=jL>��'���Z�[��:*�T>V5?�R/?�n�>8[k=� ޾������ ��J�=�?�2?E��>���;>��=<��=�z�l��=�KR>�uI�ԟ���.�}���J��H��>̌>�x�=���>"�?>:'?��>�|�� �Y�����e86�R���J�K>��>ʏ^>�|T=x�;@�C�'r���w�~�zB�&1Q����~r>5Z���,�>�y�=��=�*<>t>�=�2ν��k>!R�>�>
�>�'?��>ZYF>'���ib,�ƃN?n��>�ъ���o�{�J��?p�����&8��0?�>	��������6{��H^?�r�?�U�?969?��3>�~Ѽ��,>
�<!H�>H��=�Eh���s>� �ϖ�W�>N�`���K��yx>�g>�L>)xM�G��c���ͪ=��̿��k�ޚ�=��?��J<�3�z�M����нPRn�A�p��G���/�Խ0k<��;&�D;��[s���羳���%�?wIc?��>�ټ}X�:� �����}������W�I�æ��.'+������ʾD%�����:���>��M����>�zY��@��$�|�'�(�����:�?>�*/?�jƾkд����^g=jY%>���<�?�ث��$���F�
�\bW?��9?�P쾽������>u�?`n�>��%> %���5� �>G=4?��-?�u����Q=��[���!j�?���?��??e�N��lA�h��I��"�?m�?�8�>���[̾���B�
?u�9?#�>�M�+\��-=���>/�[?o�M���a>��>�
�>���z��.�Z;��α����:>(Y��K ��h���<�^ҧ=+�>�v>�5_�����T��>DϾD�3�8I4����C�4�t�A�c��>(�X^�����=�[x=H�4����믅�����p\?+[�?�2K?��1?.Aq�,p����R6>�Ӵ>�3!>* *��{�����>@��>�9��z����?���?ǥ�?cvK?R�k�O�пQ���q羖���B/>ǣ�=�J�=�e<���Z=�n=�>3��+0�ˈ>���>0�H>�F>5 A>z�>���>z���6������X��X�I��i��������N羁3���i=�������ᰈ�8M������8��}0=�b��9���&!?���> ��>���>ꬸ>�I�󅜾�Ѵ���ﾫ�ξ0���Y�����ྚ���񈻾���� ��;�=��^L�>���=�:��^x?�u>d�>��k>���,��+>�F
��ޑ���u=$��=�*>3��>[͟>���>��=)�|�ȗ����E��1\�`��<N�9?fr:�,;���u!�$�ľz/�����>M�>l0,>�v,��$������u̼>�W��e_d�I���	_ּ9��> �>��7>{����D��MP�����9/->�"�>�^>j��;�M��Ϯ��=L��>j�־���=�Ё>�O)?�~t?�r4?��=�a�>p#a>.�>z��=v�V>�2T>Ls�>A�?�6?�0?tn�>Q'�=��`��Y�<�E=�>�U�?��5��;n��Tc��֕<Z�>�Q�>=�*_=��;�g=j.E=xa¼��;���<>��>�=?7�>�U�>�Rv���=�܎C��K��`*>h%��@�>NA�>5�?��>���>VM>�!Ͻ|�����P�>22 >!9\��4q�"���Mт>�h�>�"U?��(?�K��:�N�4�X=]�>��>N?��'?2��>y0>��Խ���d��U�K�P5	��9<_\��^�/��j���
K;�HX>V��W�����>dR�>��H>LB�=�ں=;�>Y_|>,U�>�@�>Y>�M�=�=�$�pU�]qi:*��:_�=�./>�f���͖������@&�s{ƽǽ9��L��t�?~�2?#kU�aZ������W���&>� f>B�>Ǔ>����Ǎ��Al��[�ނ��=��>cZv?��>�Ge�N�<4�>�*>y-�<F��H`>��1�����Y &�w�>��>�D1?�'�>q�=�����W5��"J1�I��>E��=dͰ�O��?8�m?�!M��hK�8R��a.�q#9��¤��ȾmѾ�Jپ�Z0�ŃO��U�^��.�rM�=�K?Y��?f̽���<t��B���>��W�;P���Wl���>��߼�8�N�������7�rv	>�P>/�>���>����V=?��F?x!R?ru/>�a>f޾>�@7?*�F>K�>A@?�;?��?P�y>�0��<yD={�$>;G�>��;��^��ڃ�h��=>M�>5>F�<`h<��=��.�),��雼�@=���=z�-=Ei�;�3�=��>�$?C�#?����7������x�;;> �>b�>�=;V=�S>!��>��>L��>I��>��<��������\��k�s�?Y�??�l?�Ӊ��_�<)�'�'
�]k�=.q>�=���þkb��g���A��>��>���>��>�?k�5?���>���F_R��<W��(�����>�3�>`dx>=6&����E�|�w�ߋ�k�y��ؗ�`����C=���=:9�6�VCM>� >U��=�"k>���Jj�=I�>Ur�>ܷ�>���>�;�>�ʇ=�����3��:M?���>a�H`�]98��G�>���@}���3��+~>Y=H���k�ƿ%I���m?���?K�?��?-'��j�2����>31�Я�uHm>�8�0�Z��!d��#�>�3�>��<ч��|��=g�=5!�=�r:�W���e�@��������Q��y۽����o���k���s�
�ʷR��ڽs���:p���1���6��`<���A�ǁ���ZԾ�f���?(�D?*�>�r�<�=�8�¾��Z�ə2��!Ҿv����վ�l��K鐾⪾�����쾿7"�9�2�ޟ��>g=Y�*��Z�|���(�(r����?>�3/?�,ƾڬ���y�_�h=<�%>�3�<�=�<���m������^W?��9?�f�B����T���>�?Os�>#M&>o(��"� �>�-4?,�-?������%��Y>��zi�?���? �??�[M���@������@?/�?�{�>~%����˾P��0<?��9?���>�(��@����ĭ�>qZ?��N��G`>��>��>�콺䓾��&�����j�v-:>2��{2�D	g���=�=�=��>��x>��Z��߬����>lGݾ��=�t�6�+z��/�窽���><����n�=}%�=�/�S���^���P���$RW?���?�oB?��.?�Ǡ�����CU�>��=��>r�<>��N<�uY��A�>���>'� ��������d#?�$�?��?gEG?~�q���ڿ{���ľ����Cz�=��=��;>v4�����=<ڒ=��3�i�Ļ]*)>�,�>:.l>5�h>�OK>��\>��f>��kN�����ǡ��$\6�2�
���
����y��'����!����匩��5���I��T�@/��S�<�1Ծ���=�?;R�>%}�>�h�>�q�>��>��w���� ���������E쾦M��s�v7����J�]�`�����ۅ=ϐ�ǐ�>{q�<�>�;!?��M����=��>��"=Թ�=gka>6b�=GJ>��>��>�!>��C>��l;�܁>5��=̊��EP����8��N��̅��6<?
�g�e͑��&0��辽����b�>U?��q>��!�#J��#~u��x�>1%?��ob�&�޽�OF�\��>R��>#��=e�s�Dd���V�b�佲��=>d�>g?��6�����VZ�=���>��־��=:�{>�*?��u?�#6?+��=���>ɕe>k^�>���=r�S>��W>B��>2I?g�8?t=1?a��>Q��=c`����<�6=��<�eeY�|!���/������;�<����OF=�z=���;�W=q�4=��ڼ���:���<�>��:?S�>�Z�>�J�jr?�H�C�N��8>�̺���>j��>�y?�u�>wd�>�=)>~���c�ݾZt��>��/>B�Y���x���Ի>�z>S�x>�X?�/?���9��B=��>�ޯ>b}?�,?�t�>�P2>J�����
�NͿ���Y����k�=޵�&`C=S�$�!�j=d�@�����bǽ�:D>���>⼋>Y�9>��>�kk>��>R�>��,>M�K=��=�dT=�2=�*���=wBF����Qg^�/�Խ����3�r`��G׆�mwu���7��2��N?M�.?�v��n�J����	����z��>�`�>�d�>���>�V�=I<��v�}�?��[]�� ?j�?��>ꏊ�f��<Q�K>��<>�%g>�h>���=o�Z���W�޽->�=
��>��K?��>�]��b	������"�2�w)2>�>/6ǾdĦ?2�x?`@���3��yɾa=�5�E������8�Џ��A��t�:��(c����u�:���)=9=
?-L�?�Ͼ�Yy<�s�9��4Ȗ��꾲�|�8J���i>����޾
�Ⱦ�z޾�����_+>oI>֣>��> �=��?c~ ?�	l?rm�=P�?x1�>f%?���>�?�8?�7G?�&??�A�>�73�vFf�id>Y�D>$>��1���l'=�1>{�>{>/>�x�<�A�=���=.j��~½)�<���G=V<r��S=�>eH>�	?�$?��ɽy����[���L��PQ=IU">��L>��<gg׽^W�=f�>`��>d: ?�H�>J��;%5�Q$�r�ZJ=�*?
�+?j��>���<��=C2���\R�`�<E�->�Ҽ�G�BZ¾,��%g��XP�>���>ԳA>�D�>�4s?XC?�i�>�ɑ�LHJ�Q2�f;�to\���^>��?�c�>���=c�پ�t.�i�/�z��h�s���7���I`���:>�ұ:u�=}շ=�u>y>O��=�ރ<Hܜ=\u>G�>��>�%�>N6~>N';!qܾq���8G?6#o>�e^��1C�ʰ����>q���&������r<�=���K��7������J?r3�?f��?�l?Rӯ�v��ǘ>�5��(Խ��Q>��L���= A>�>�>Bti>�->֧.��ѼȨ=�>N�Ig�d��c�h=�Ԯ��`�o����Y�U?��4O=.z��~N�<}�a��gȽLm��o�r��tW��O��{����z
��M�ݾ$�辗X�?�#?3��>S�=ya�ڴ޾�:���]c<�@ɾ�'s�f쾳���C�����Ⱦ����$���<I𾹼�>y�Y�}7��%�|���(����r�?>�0/?�Vƾ&Դ������g=�[%>.�<�Aﾽ�������*��SW?%�9?�b쾽��:�ོ�>��?�p�>p�%>�D������	�>�14?��-?��[���7���+��)i�?� �?��??�O�xA����ߗ���?R�?���>xÊ��`̾����.?^�9?܈�>�r[��	A�!��>vg[?��N���a>6�>�g�>!񽁐����"��"���Å��a:>W��@����g�*=��ڧ=?��>�Xw>T�]���Zx�>��羷�;�+Z%�GS��W��3j��ʽ>��ξcw`>4T>�k<�w8��J��[�����C7G?ᙶ?�)^?�4?$�þ��~�����>�]>H�>Ⱥ0>W��#��>�>���i�t����?/d�?���?�h?b�]�q�ӿh����]���-����>]��=5Q>r$��o*>�B�=�_<�I}=V�,>�|�>�6s>�r�>k�>�d>*�W>r}���-"���d��}�E�	B����.�N�w�ѹ��l�J�������`������!h����Z��Q���#����\�>>�?���>�>G<><`0>'Z���=x�����|���� �.��ytžy x�$)�T�\�\W��6ն������?��.<
�=a��>	���
>X��> ׀='>lF>h�>�G>��6>��K>��&>w"Y>�~�=���>��>���E����|�_lؽ���9-P?vrh�������@�7F��8�#���>�h�>��p>E`+�����Pc��^Iw>ŷ=S�A��ô������;r>��?c� >k¬<��)��.˾7�P���>9y�>x^�>�� >���=_U��꛾Ρd>G9���>��<>�35?M�e?�^S? �>W��>� �=��I>Tg>�E>�{<>%��>1�?�TM?^/0?�>�WG=�`t��t=���=�nq�Y�4`ν�xk���=�mi=4����<g�=�`<���<ϖG;�����򼏿�=>=?a)6?�zF>�zw>Js���0�c�J��i���=�==]�	?|d?�Z�>+��>>�=�����ؾf�!,�>b�>Mi�m[��'��=���>0:�=�/#?i�>�#d�_�羨���P�>ƌ?��?x�R?Ҧ>�yB�G�Ͼ>���aӿH $�e�!�7N���+���;=�<�ĜM��zE���-��x���n�< �\>�)�><�p>�AE>��>63>-;�>�XG>�+�=ץ==&�;O3;�E�n�M=-��@I<6�Q��z���%ż�ї�H����I�.b>��y���׼�M4?'K�>_��x��>V�1g�M}��S�>lG[>ĈF?���>�XȾ�H��B����x���:��$'��hw?��Z?Ҵ��#T>F|��NQ��� ?.pP>��;�}>�I�n\���i�>�F+?���>��>��{=Xo+���e�9>$���t=�+<U �SE�?�wp?�l��/�=A�B��}���d����>1����¾Rչ�5�U�^�z���(���I�>�>�R!?^��?�"�s_�>؄־����R$�v۾3�>���>�)'>q#A�9|����)�O�jܾՉ���>�?��z�!�H>
 �>�V>�\?<p�>�[K?�3½v��>Ѹ���_�>���>�@�>�?�6 ?{�>d�?R:E<��]��L�@گ�IN>YR8<Y�]=��	>�u>��=y�>��>�ق���u=��ܽ��9���i�|��Y=�D9>��O>�?��W?��վ	����VZ=�^��,�=|�b>AiQ>O�ܾ�G����<(��>�5?��K?n$?��5>�]
�e�=��M����#�ݴ/?�KJ?�&�>�:Q�R:g�Rm��������l��>j;�;�|8����-�yi��$׀>ş|>�6>� j>��}?�1A?w�"?�2����/�}w���)�����{�4E�>& �>�6�=Q�ܾ�(7���t��a�ZZ0�Z�(��D��X=h��=8�>R+B>��=�>�V=ꏗ�>�ڽeX�<\@��c�>�Y�>�?�5\>㡅=�_��q@���I?���-������Ӿ:2�z">Zq6>�Q����?����~�XD����=�Uj�>֥�?&X�?�e?|�=��D�S�^>/qP>:�>�z<=FA��M ��tp���2>���=�v�a�����;Z\>Bfy>V�ýx"ɾ�x�,�E�Y�пX�r�VG�>	�\�ܴ��Z�L�n.�B��X���f� ��s;���1R�8ヾD 	��I�-x��C%��Gӏ��?�!�>dS�>��;�+����ʽ�/.�R�8=���>����Ӄ��2�.���FپZf��je3��@�����Û>|�Y��@���|�.�(�$���>{?>|6/?�^ƾ!˴����g=�W%>���<+>�կ��P���W��cW?��9?�M�B,���*��>��?�s�>e�%>�)��?�'�>�94?B�-?9�뼱���8���ٓ��k�?B��?TR@?��L�>�A�G�(e���?�W
?���>�Y����˾M��q
?G�9?$�>�,�/�������>`�Z?<_N��]d> �>�7�>�^꽼���Y)��4��I�����6>�*2������e��18�(�=�*�>�?z>�^�oU���;�>�Q�d��Xk'�t��!>&e3��{>/����>1ҋ<d �=��1���G��[��S;?�#�?�&(?��k?�K	�}Ҩ�%eʼ~�����>�Lj>m@�f�>ۡ>®>v��j�\�!� ��*+?[�?�<�?eS?��Y�Ԩҿ~����ھJ���5��>��$>e>I>9&H�ʄ�=��1=#=(�m��4> �>�Z�>�.>���=�֒>7��>Ih��ӻ$��ұ�Pŝ�q&��$-��-�R���~o'��o������޾2ҝ����=�%4�S.��܎���I<���:�˾yU>[C?�,�>f�>
�f>�9>f�L���u|���ʾ�C��;�1ƾ��߾���j~��o^��lm��,(<�0!�f"?�>-�������?�򽞥�=z�>�5>�;�=V)J>�]�c��=�j�= o>�bA>� I>�8�=�C�>�n>�~�*����r6�T�l��e1?k�����!�-�:T���{���C`>���>\B>�%<�飛���z�C0�>����Z%�:{�87F�j'>�Q�>�">lp��/����fk��43�:��<��>|��>��=�O���	��jw�3��>�Ͼ ��=�q>)'?`t?�4?��=�p�>_[>�`�>��=H�O>�L>�Յ>bR?��7?�80?]�>��=@�]��l=�)=�V=���V�o�������+���2<(�G�j�A=�^=�r�;m�T=�A=������;�x=��>A�7?^�>w�>8;���>�;M���{>](��@�>���>D�?q��>�,�>EH5>Q$_���¾�P����>�B>Bo^��w�s3��Dv>n�s>�O?�w1?%Rv�RPb�D�=:��=�ܭ>��?�(?���>Rb>M������DFӿO�$���!�7�x���MS;j�?��PV��l�9&X.������r�<>�a>��>�m>7yB>�U#>8�4>���>�_I>4a�=�B�=�ޱ;��8æK�"�H=�"�H<�S�2���Mf��=�������}M�(�=�����V＋T&?���>��'� �L��=̾��/�M|��7&?��?%?�� ?c�Z>�@���q��R�p��5��Ue�>�k`?��?�1)�y��>�v��i�@N�>Q��>�?=-1�p�e<3ꆾ���S!?��6?.C�>>鉾�#c�|����m4����>#�=�0�Q��?�]?���(m�/"�^RG�o���oK=���2�Z��{��� ��:�W<����DVu�陻=~�>�7�?��j�{ �=��Ǿ�'���酿v/����=tU�=&+�>��G>b�;��褾��WȾ$=����<�d�>�gL�U�?��/>-��>7R9?���>Q�=?��>���>#��I?�0	?��?3>gh=���=Ia;>�m?>}�L�"�=j�=C*?>A!q>GM>%7�� �=��;=�b��v��ݏ=���=!��� �C�=�]=!�:=|�?=�?��!�4o��X'�՜���Bջ�s>�=�=F�K�.=��G�<��>��>N�$?���>�Z��F��������L٢=y�?K�:?6�>�D����>�B��a��m�0>���>�<����2̾E䋾����ϛ>���>(�2>(Eh>j}?8U-?��?���I.���e�
Q�N�˼����	�>�#�>���=^�ھy?.���h���^�y)�M��|R���<u&�=+b5>	�Y>���={6
>wz=[���a���?��W�Q��> 0�>��?�nR>l�I=IF��&��"`?�,D�����n�=��0��$��N��\�c����TB�>~��{��L`�����L?/��?�ż?m��>��3K{=�4�>3aa��W;7�=,���?�=�y�>U�@>D�W�>t(�Z��<n�=:q�=��� ǋ�E�E�u�d=��ҿ�+O�eX@�qo���ʻ;J���þ����/�Ǿ83i�?���^�;U当�g>��=�+½�f	վf�&���n����?�W?1(�>�a�=6�2��dʾO�����<]����o���Q���������0׾T_޾'ɾ�����3��j� ��>�rY�U9��&�|�m�(�s����r?>`//?rfƾ�ڴ�ğ�Ccg=]]%>���<89ﾋ�����'�VW?��9?�c�2����5�E�>��?S`�>,�%>���O����>�34?�-?������D1��H��Ad�?���?��??��ؽ*?E���%��c3����>��>�j�>q�;�)I���Ľ��?�"9?k҉>9t��R����5����>QSO?4�R����>���>:�I>�ٵ�4�V�aŽ᳔�>���e���W��C�+�|�"W��A�M>���>�<I>�����
Ҿ�1�>K��}�����2;���>��n&�>N�ξ�C>�_<��=��*��&��,⓿�ý�G?,/�?b�+?�Z?~(�pJ�T&�=�v�
�>X1�>�ս�f��a�>]E>\�1�ow�%l��\<?+�?��@�rT?�p��5п'����\��m��-�=�d>*A�>㱽�r�<�����$�;}.�&>�>���>��d>�+>�o�=Rb>�"��_=$�ܪ��\ד�o�R�y�=�Sn�ԃ��*(#�!��8���h��(����&u�1�d=��ѽ�'�����zV��M����<>%B?8�>0��>�@>7A!>��f��1�|h���̾_��%��s��9�\���_���y��`&����=Ge&�"�?�`�=x��m3?ЕQ�w�>��3>�3>b�>n:�=Kf2>�z=�,�<��0>��=�->u�=H
|>la�=�&��Q􀿒r:�rR�S��;��C?)+^��t���3��$߾�\��m�>�?�8S>��'�������x�;��>��H��bb�h�ʽ^���=�>���>x��=�wܻ���Jw�o�R�=Z�>ă>��g�TƏ�xU�h�= ��>�!о0�=��r>��*?��t?g�6?���=���>��j>��>���=(U>�,N>���>;�?
�8?�0?ߪ�>ҁ�=�k[�z^=�/=i[<��|@�٬�Y�߼���O�<��U��R'=CI�=9��;z�N=�U=n��ٙ�:���<Z��>�I9?3�>�x�>s�4���>���L������>[
����>�v�>k4?4��>A#�>r�/>a�y�΋¾��㾽��>ڻ?>��]���w��d�L�>�x>Y�M?�N0?�5`���e�T}�<��=�H�>��?~�(?�l�>Ȃ>�����B��j�ɿ{J����~��ط�g���(`">�M��2��=������-�->���>��>��>�<�=$A�=H3@>�c�=���>}�9>�˾<�7E=�R<9�`=�LȽD�=���=X�[=9νE�*�W���y5>��2��H =zm�	;�_u��)?&'?8���̸=�8d�t^�Q&��Ա>祉>9 �>��?v�o<W���\��9�Z�挾�w�>-�k?��?��"����>���=*,�4��>x� �µ=a����G�=Wb�J7E<�0?��2?� ?�yW��c�_N���QQ����>ll�<'=S�ak�?{�M?x	����4�jG7��?���Q=0EC��n�/ŷ�3@>�I:a��� �nG�ľ�I���u"?��w?�%���O>4{��c��э�����=�`>��>��=[�<�-���������]�߶k>�P�>e��=�?���>�h�>�a?
�=�%?�y��a��>eo>��
?b�
?�z?dY�>�>�u!���Y��`�=~K>	���9�J�ܳ�=��Q����=S_?>{�a>RZR���\>j��=�q���ݼk�=���=R���=E�=*a�<z�=?�,?��,�V�]=/`���������k1>-yw=T��k�潘j�=Ț�>=��>.X&?�T�>�M���;� ���m���4= ?��E?W�?ꥅ<��=aƾ��d�ܛ�=t��>M��;�r�h5�ǫ�Xt۽s�>�>��v=⃳>��?�\�>r�2?,��w{���e�&����F��{�G���?�j�>��=E-E�������f�Id�����9=�χ��w��� >�DB>^=A>fm>lm�>���=���3�ĽC�>��=Z7�>�j>��?Ai>�}	=q�1뾆Et?bc�L�@��ƴ=nJ�c��>�w��<V?��9��\�>��,��"��쩴�з�4W/?n��?' �?��1?[h����5h�>��d�uށ=/��>�����6��>�>��0WF����>�nb�K���oM
<}�>�If��B{�Cpk=�OL��x��%�2�� >� ���C����Ѕ���F��u��E�����MJ����������D���L�+ט�p(޾?�ݾ�N�?�؜?c:?t'>t�	��w�#@;�{>K8о�;��vRվI�|����R��������X�?�2��h��2�Dg�>]Z�����ɨ|��(�A����=>/?Y{ƾ����Ź�Se=ɒ$>���<�R𾹚��4���ޛ��V?�a:?3����ߴݽcf>��?{��>Nn$>Lȓ��R�e��>)�3?Q}-?�' �5�����"���v��?T �?Y�??^L� ;A�7g��;���??p�>]싾Q�;���R?�\9?,ɼ>��y?�����N��>Ma[?@�N�Ba>ĭ�>�!�>��
���+9#����p���I9>Y~��Y��Me�j<>�2ܩ=���>q-x>Q�\�>��L��>�����Ѿ� �kK�q��=��&��;��tߌ>��A�s���W�U�Jg���N��_ɇ��L?���?�=?try?�*�&&��y0<�Ͼ[�?M�=��[=S��P�>��+>J1����N�=�I�x�?�:�?�/@W)�?��W���̿b��0���NFվ;��=�&�=��~>Z8����I=e)<U�=�1�;�}P>V�>��B>�#w>Y>x=>>�U>�R��^)��j���Z��XI��&��f	�Ԑ��P������<H�����.��� �����q~Ž|�@�̈�6�g�?%����>�&?Y�?���>�����
>Z?���J����y����`�����������V�ľϙn��^��.������=����W?&�;�d@��o"?�8��I��w��>�|�=��P���1��}<�З�j���B�=�> �>_wS>ɂ�>)d�>a���&���F7�?c��g���=�`?@�ڽEɾ��5���Ⱦҭ�n�>��!?��'>��-��ޝ��ʎ�2��>&l׼�����Y�P+�<���>�ͭ>-d�<v��<'�I�َҾ����O#>��m>ȯ�>�B>}�l���St�����>H�Ҿ_u>�u>fH*?۞u?<^6?6��=>�>oC]>�>�ڹ=><Z>8�b>t�>ne?��5?�B,?���>Xs�=�5g��p?=�h=��1�d�!�?s��V��� ������$�˧y=�15=ek��ab=q�G=�����;�T=��?�EN?Q��=�e�>N���iT�H=h�6��=�K>��Q<}]�>C}�>[��>o�>���>Z�"�������	�5���F
�>*��>�Y��Բ���ڀ;�>�?�}Q?�-?��0�Z�ݾ(�h>��>�#4?�\m?V�<?��>@������	�ؿ\���jF�D�<=n�-<H�>�����V���q�������c=�A�>�>��>�b">�i>;=D>G��<s
�>І�>7>�>�K������� �iў=�В>Tg��%�Lf
�"{t����=�n�������/�*�e:r ,?y�?�F���d>F�ؾGU �'�?��'�>��.>ވ^>��?����W=�ɍ��x�;�þH-�>�f?��2?a��
�>d�[�򾲾�=�>�=�NA=]v�<���>�`�x*N>�`?]%=?�e?M�+����=���_��M�>uL�<	
��J�?m�`?�t����=����H�h���� =���ng������!�k�>��>����L{�Qj�=р�>���?!�l���=glξ���t���9���^=M��=fp�>4�%>W�A�?מּI��OA;��G���4=��>�(==�>X��>��=��O?��>C�5?/�=#?Y 	>�?:2?���>c?��?Jw+>B�Ͻ�0�>�>:#M�@���j�>$���/�=�G3>T��=O\�����z׼��`=�R���v�=�5=0������<٘�=��=H��=�
?OU?k���W���V��T4��ȧ����>[��>����'�qw>?�>I��>�;@?7&�>N��D��	��y��W���91?�J.?���>�J<C�>��Ѿ�+:�A0�=��>�=5)޾,����믾�G��OQ>��>>C�>�]h>Q�~?@,A?C�!?,����|/�7w�-*�K옼��=�!8�>d��>w��=Ԑ۾��6���s���`�F1���+��'F��Z	=T�=�A>��?>��=�>*$=����^kؽ��$<��`��'�>n��>=�?��Z>)Ά=�����;a?-�+h߾��q>X�Q�Ű>��g����=��(���?_���c��渿�푿-O<���?9��?���?���Z���q�>��"�'4>�f>%���:d����>M;ƚ���+w>x���*��48\>a�>�����ܾw���ti�=ܷ�;�E��3<��G��zA�]3�
����ך��7��ձͼ<�Ǿ��Y�� �N�%�����\}m��bþ�����?�o�?g�x>PR$>�� ���&����D_>T$�������վ^l����I���j�V�[D ���1��Z"��>�_Y�Y?����|���(��֏��a?>1/?%Qƾ?ʹ����lg=�f%>֏�<�0ﾞ���&���'�RW?P�9?#[���K��:�>��?�b�>��%>"(��$�콐(�>i24?ҟ-?���G��F5��=쒼�m�?���?��??S�N���A�=��w�<�?��?��>�M���̾Nq��#? �9?�μ>���J���9�9��>�j[?0�N���a>��>8�>������S�#��,��𻆼s�9>��e9�Y�h��>����=	ؠ>�Vx> �\�𼮾�T�>9������=���;���>ն��^�>'���{?>�}��\��C*��S�������??��?]�?�im?ߕ���'�%�=ƅ��3�m>)��=X���%�ҽBi�>��<>�~���*}���d�M?�?��@Ȍx?&#@��	Կ�Q���a�7���]>/[�=��>� 1�}%6<B�>�L�=R=�=Aq�=B��>}f�>��>�]>�@�=���>�y���L"�op��s�F��� �5l	��8���{*�3�Ѿ�g���r�'�����-]B<�;�=�״�1�L��=�ɾ0P>��<?uܣ>|�>)�>{5P>���y����ľ�����+�%
���>�`��.���^դ�����u�R��=��!��w?�1�>�����1?!�� ��>:�(>�!>u�	�I���m3����=�=�_�=��S>�z�>��5>z�>�Z>o�r�}��)2�@��T��rC?��u�-eɾ��!�7g����R���>J��>Ը >�t@��P���wc�Ɣ>��������.�����o>�S�>�= >��=�Z���U�gʽ��=Z�>�Tp>#W.=� _�C>��X��@��>�Lо��=^�r>()?	�s?ԫ5?o��=Ρ�>�X>�,�>��=m�P>�KP>.d�>a�?�6?�y0?D��>�L�=ɭ]��=��&=sN9��Yb������B+��x�<�M-�<~==�zW=�A2< �T=~C=�M����;�q�<���>G�9?\��>/B�>��8�P�>��vM�����>��)�׾�>��>�?���>�0�>96.>���U�ľ�M�U��>�3?>q%_��v�]��?�z>Ѽr>O?/�/?�5��FSk�t&�<��=���>Qo?Fa)?�]�>��>[����e��Uٿ��ɾt�B��ق<��5�wy>ˎ����|�sB�=�f:�wW�=Y3>��]>�|R>Ә�>�r>>x�
=�&>nU�>ߞn>�P=޷"����;�=Ҧ��7��=��=�5D>#m�=�?=�7�~�k��d���,�yL3����J����.?ud ?z8T��Ë�\u���.%�۩�����>�U�>��?�?���=�����Y^���E�ܙ����>�s?j:?���ۭ>��'��h׾/*�>&U�=�Z�=�o��8��#}��_.�=/%)?�u??�O?�	���=g������[���>�<�A�j*�?f\?��5�����n@��q�T�<�,�+ ��-|���f(�T�@���.��uɎ�� >=J�?xS�?�Bg�V3�=i�JA��i���.���e=��=l��>�8H>�k0�Tɯ�+��G�¾X�d��=��>��J=���>�FV>-Z>dWe?"��=-� ?������>�:�r��>lM?$�?�V�>R{8>��S��D$�hU#>���>{�~�M�y�>��i>`!>tr[>!���8�=���=�j/��޽��=׀=댛���d=�-�=�Zo=d�>P�?�.6?k��Z�̼����L��Ϝ��{�p>��}=������a=,��=ňx>h��>U6?�Ot>��H���>�۾��U�����?�L?�?�O�=�OK<f��� ���J��=[��>�G9�b��yh�J����@�>)��>�7�=��G><�{?f$?���>�[ҽ��'�;#Y�t���cѽ����#�>�"�>ɑ�=�/����%���b�jAd�Z�1�.#���:��9$=���=��3>�C>��>@�M>��>X̽z#���ѽR�׽��>�k�>?.`�>,�T��ϾyY.�{jk?�(���	�w�>&�@��o.>aϏ�.b8?�7>f^0?��&��5���aĿ�ʙ�Z`*?ґ�?���?�[?)(ؾ�
k����>���%��=��>鑱�S}�=E�>�>��b��fu>�ļ؅�=2�=I�	>."a�V���c�BU>�5��15�>j>�9�,��~�پή����ަ:�����g7��ȓ,=�J �e"���Eþ����Q��V�����˾�Y�?��?�~�>�D�=9��4�����so������3^����پ{B�yC���x۾���� ���Ih+���7���?�>� Z��e��|M{�د(�8:ݻ�.=>g�.?�7Ǿy2����GL=�!>K3�<��e������o����T?-�;?�[�:���Ծ׽�a>�??��>�m)>�!��`��e�>�3?\�,?�������pp���1��?�4�?��0?��=� kC��q���p�|��>�}�>���>ѿ� ����~?��0?���>C7Ǿkm{�z�!�j�>�'[?�]��F>�
�>�$a>�*������࿁�v���͝�=�À=ȋ׽��z�K��=��=8�>-�k>��^�<Y��%?�����R�#�n��KO��,z�n�%���>���>�	>i��=��>@�}��#���%���̼��c�?���?9kB?HI?N�������7�ӾZ���?�Q�>�4��:Z�=��?���>�9���96��و��p�>uN�?�`�?Ci? )h��ҿ�<���d��{���oC>%��=^�>�f�@?=o-�>d�:=ɲ�!(>�ҳ>�*>ω>�F>K�$>�c7>)���<!�@W���u���3�ڨ�F2���z�����~Y�q�
��Dݾu���N���ɽ�+����v�n@%�%P��]�fE�>�VZ?D��>cϚ>�n�=3>0���������0%��ce�@��#���2��V�����Ⱦ4.�)-��^.>9,��p��>x�M>=�<�?�b&�P-�>�mj>�!Y=�>&��>��]>D��>?��>�>��=E!>*��.p�>}�=�����.y�U�4���o�zB��hvF?��C�i`��2@��쮾$tT���>{�?ߒ(>�9�;��([s��ٲ>�FR��OBb�m?<��>Hu�>`�>�Lֽ���]"���Q�]�=���>��>��=�{��C+�m\�#B�>��Ҿ�2�=��t>�.)?�`w?��6?vƙ=�`�>E"Y>_��>���=�.P>}Q>FՉ>��?5�8?]?0?��>�+�=K�_��=q�9=X)8���d��껽z��T!4��w�<Md4�&�D=�[k=��<��h=�VY=fD�Ͳ;?�=J�>x�7?V��>���>!w=�U?�u�M�i��!!>�ܼ���>/c�>B�?50�>=��>�'(>3K���{ž�?����>��D>N\���v����>�i>��M?�-?h�k�8bj���<?��=�"�>��?��*?�N�>y>X����1�.gݿ�>��o6��w�=���=5@V<R�Ⱦ��Y=��>��>Q&�d�=>,�>ޑ�>�+�>G��=�=�=-��>�g>�>w{�?�6���;x��=���=��=�u��Ķ��m@<���½������i=Wρ���,�z?�<h�%�1XD?kuO>���8>T����[��Q󾵎[?۪?Y�>I"1?QT�>�!����J?��q$�s�>vaS?��E?C�I�=DE��\%=\)�=�#'=N`�= X����=��=���S�>�E5?�o�>I���I�b��N���.�G5[>|��=�kϾ���?�?�4���Y��oM�ȁ�o�e�����6�79���F��q}�\H��b���/�x4���Z�=�|G?gJu?1���E�i�¿��H|��F��������� >�>�~�>�;��!�R�.�j��j�=��>9E?L�ݽ8h?o?Ɨ�>ATi?�wW?�5]?�C��]�>�PU�7,m=%�>�
!?��?��?@�>E'>:�
����=�*��5l���=�H��VzW=�>��:>�f����=��=(�=Z�x��8@�������(p:C��=�v=�Xd>�a?
/??V�&>�{ =�|���0��h�>mh=y��<�`��d��=DY�><�2?�?ò�>E���7��N)U�9d�y�@>/e?�}B?`?x��=���>e&��=d#�����f>g�����B̽���b�:�{�>^`�>\�N=�5i>%�}?n�??�# ?����/��'w�+�)�#������t�>��>���=�^پA)5���s���a�Ȇ2���D��F��+=�0�=|�>͗E>�k�=��>��&=;���#p��Q�;�D¼���>>��>kk?/ze>9�z=
Ӫ�h��W?����K��� ����6�j��J�����>��?��*�>��>�
=�tާ��U�TӉ=�L�?���?���?⯂�Ap��a>I�>���>hG�>ݠ�����9^�>�7">�Ĉ���@�5N���>W/��'��>��\>QZ�_�����=��A��d=ѻ��lS���ȾB+��8ݦ�6�¾�l�ϙ��"6����� �CWT�������Lƾ����}�?T��?5��>��H<mF2��T�?� �!g�	��/������t�E����zf-�:��LU�Ƕ��e�>�<Y�Nr��|�y)����ͥ=>H/?{tľ�A��q��]�u=�'>�"�<�ﾘ
��"��������W?Μ9?/��!�������>��?��>��">�M��F1齎��>��3?��.?^�Լ3n��G؋��ר���?`l�?�nG?�e���^�Í�gE[�բ�>���>K��>����v����r+?�XV?~X�>���>����1�ss�>�hF?��K��&�>�z�>��V>B��<�"Ľ�0)���L��o�(��=�(�
2��_	}�ْ�<*�>?���=����)��N?�{ԾV7f�����^����$倾���>�"��z�:>H��>��>�\��I�������h���v)?��?��3?W�?f��H��.0����=ת+>���>�R-�&���^��>���>�� ���u������>���?lN�?�ml?���YNӿ�V��I�^��6C���>�h}��E=�f��OQ=���=�!��i���@>?B�>Mw�>I�z>���>��:>qcY>䢂�w������⌿�wK�Ȏ�C�)�{�z��畏����󽻾�����ɬ�^ؼ�m{��x�̆d���N�ȃ��ퟺߴ6?%.�>H�R>�,=��4>�i���������ʾ�H����8�/���4����D�ƾ,zξ�K> �;����>d3�=<ɛ=.9�>q��;,w?iZ�>�..>" =��?C��>�6>$;>>���>(a�>��>�_H>���>A��=́��ց�J35��n\���:�҅A?�U� ����$@��I������y�>@y?PU5>�l.��B��P��[f�>���)D���A�E{�#[@>��>�ZB=�k��ϓ���f�����h=��e>D�Y>�P�<������)�b�<O��>X�Ծ�?�=!�v>�.)?�w?'�6?*�=���>�_>��>���=�LN>u�R>�V�>Y�?�k9?��0?c�>�e�=�7`��=��<=d�>�pf�͍��C{��j'�\��<Ø$�V<F=(�m=*��;t�[=�!G=��ü��;� =|�>la7?�m�>��>�?F��>��CO��{���>��+��S�>���>��?�[�>�0�>�� >C܃������۾���>ũH>ϛc�Oz� ��m�v>��i>��L?�3?�u�z�f�/�;=��=1�>$-?,�'?뛺>v�>�㣽^���oؿ��0�A��y��f젽�P;7#��8z���U��h}�����ڔƼ�a�>o�>G��>J/W>�xq=$6(>�_�>��J>'��<��)><����7�=Q�P=�i%>�pχ�TK=2I(�П"�����0�����%�;�6���J�E�w�6?N�>����} �1Ts�'���6Ͼ��?�M8?36?h,?.��>p����*Z��:��$W�n��>;�-?�u:?*�ؽ�6e=_�h=U̦���m��FW>U�Խf����g�>*��۝�~?:Z+?g?D��M������}N��g>eq=ǣ��%Q�?(�u?8�F�8���ޢ0���оɺ?�`#�>`�U=���x�A�.,U�� �!T�/3"��s�>ke*?*�?H����,��!��+��T����(ý�,>H��}�>�̶>k琾����HN�'�<��Ͼ�m�=v��>��w�)?�)?�q>N�?�[?#Qr?V���_��>p�=�L�<�+�=/?		?:�?
v>-��=0[)����V_*�ıu�j��<�<��Ȟ=�};�S6>��C>I=-�={��=y'��\�ʽ�Aƽ�h&���=���=A�>�9>��?�F?l"��P=����8���T�\>��&= �s���۾4�4>^��>��F?xi?�x>�,��g8h�Gb���.>�_?W�6?/��>&:>�In>��MR���>�o%�>�-���BF� <j��G��4�v���>��>I>�0]>�l}?�A?�n ?�x��-���u�q�-�:Q�"w?��Ӯ>�Q�>�?�=;۾/q6��4s�D�b�av3��hc��E�S�=��=k>3~A>�۫=,o!>H=>=#+����何��;	��k��>��>�x?n�`>��=PN������vc?Uʹ�'�C�!���se�Dn~� @�<ۘ�>�*��v��=Z��>o�-�z�����Ʉ>�b�?�?�B�?�5�"�ӽGo>ɛ >n'?�m�>^?=����n=���;��*�U�˾����n>�b�=���>@��<����sy羍��>���\�`��� �,0��5��j���|tϾȕ����վ��ڽ,i�� C�O����ҽ�'�g�����(4��_�b�9�?��?A�>�`��^,�Y@�D�%���Ǿ��û�ˊ��N���o�������� ���I�ٓ8������9�>A�U�`��?	|�k�*�F쎼�>�/?߀��b��c-��[�=��9>_L< ���j��'��M�	�=\?�t3?_�ҾP���P���G*>9�?�#�>��>u���.9��yI>.�:?�=?,��<�㊿��������P��?U�?�6P?CA��8�H���6���*�8�?Ѯ>7�>�	>]���~ľ�L?:l?�??�!�����wB"�V^R>I"'?�HS�g��>o��>�T>�`��z���#�`�_?5� -�����>�UU��(�����#>
k�>�\�>ӪW>%���e"����>���k)@��(E�� D�4
�pk�='m!?9�¾S���?{��>�AE��w���"s�2yC?�|�?L<W?�y?0O���a	�q�ؽ����&�]> ?��J�:����>�+�>C�a���x�B.���?��?�(�?��r?e�T��ѿ2J�������A�B�˳�΄�> ��z�>�"�=b-�<.��<�KL���F>��v>���> >>H>��>�C��:������OK��`�j���(������0��N����jʽmd�dF��r�ھ�$/�W��ʏƽ,�<��z˽N4蹽���,>�?��?�9�>�y�>ݕ�>7���󹬾�`�T����U���Q���g˾�8��#�@���I�á��Vo�=S��{�;?:��=g�=!1�> ,�n	�>�M>�#�=��>W%@>
m`>>�>k�+�O,>M��= �R=��0=܃>z�=t���#��H�5�y�8���滂�D?X�s��ɗ��5��V̾_%��^�>XG?'�Z>�e*�k&���{�ʨ�>>u(�j_�#������Up>�\�>���=z`E���M�����~��+��=�؆>��>v(�<_����~'���'=�X�>X�Ͼ�j�=7�>�3?�Sl?��?���=Q��>X�H>
T�>���=�4>X�!>$��>��?�R;?�`+?��?���=y�\���|=\�{=�7>���~�ႎ��)�<oh��5
=�v�[Ƣ=��=��4��&�=(�]=�d��\<�'E<�Q�>z	7?��>"��>l�.�� <���N��;�b>��)��5�>I��>��?��>��>uO7>�l���ľ�zݾ���>U�@>��\��t�v�!��i>�r>�O?��0?crr�T�a���=a�=L�>�.?-�)?�׹>��>�������帿c�Ԓ��>��3A�Wl>q���_�>��>��<������Y= �]>˧�>!%�>�E�=��>���=���>UD>�p
>��6>c>\>����#�`炾�t���_���r�B�.;��D��p���C��R���A�w��:��3?:�z>�%K�Z�y���`����)��{M�>���><B�>6�?">���^0U�~���i�Ƌ�>G�Q?kG<?m�����J>Y�=J�L��P�>Ǿ�>�̽���*<�{<���پ������>�LX?�L�>!�<��@�gz���|��Q�>�V�= &�)��?ʩM?�+��XO�0�E�.Ͼ��=��!\>{�
<�۾�RL�X�ʻ]�1쾌���怾�t�=��A?T��?�#��Xu��!P	�Y�����{�F-�=��z=�����R?���>>找OB��E�s��4�~�*z>i�	?��P�{�Q?]�/?}.?P�y?A?�8'?���QH>�X��^>��@>�-?��e?9�*?[`Y>&�%>2�L��� 5J�����vX<��Ѽ���=�G>0�e>d2�r�]>���=;��=W��bJ�ތ�Uof�C�>NF>�����=7b?{l4?fG��-����=��D�󓍾�ͬ>'*V� ���B�8�?>���>�?��]?�E�>�}�+�U{9��!�J>
��>ْ=?9�>e�<��{�=t{ɾ��;��X�]w>�-E���A��Z���:���LF�>Y�>��>��g>1�~?4SB?
�!?�����Q.��w�O�*��F��<V�ǰ>�l�>�X�=��ھ�(6�R"s��`��1��b?�vG�:=f��=5>>�@>�=6.>�W=���ٽ�H-<����>��>n4?�]>�B�=J����L�V�M?p�վ� ��<�э������>�>zֽ��-?���=��H������iV���!>v��?���?�#�?����p��h�=�04>s��=�O�=Y��-�N��n>4��>��7�1��t�s�>�17>��m����1쟾.�ٽ�4���E���$�����}��:b��6�f� ���8�$�Q���W�Ͼe>������ Cƽ�� �o ��(Y|��3����?�\|?�}>֥�<��1-ݾ��;L">#e����8�`�˾�*��1Lݾ��ؾ�_Ҿd���|'�-%�o����_�>��\�����Ɣ|�RA)��ѼS4>G0?6�ƾΖ��=��p=pe">�N�<A���)���|��M"	�-�W?P�9?�e������U��]>��?��>_4%>;t���������>5�6?h�)?�
��掿*[�� �R��I�?�?DF?�Oν�����H�
\�l�1?(��>���>Bx�������/
�`D)?��Y?�w�>�w���ܞ��V���l>�3?Ҫ8���>qA�>��l>YH�����
鳽.������Fr>E<v��l=��ڽK.�=�p�>	�?�c>��Ӿv^�+?�Z����9�|?��$�Ɛ���粽a��>������=f�9>��r=@�M�c0�� ��!�;j}[?� �?��F?kf$?�ٻ���/���[��v2���%;!��>Y�>#�A>R��>�?9�!���X����xw?��?��?<Kc?�)[�S׿do��n=���VO��J�=]�<��>�pr��\>(�=w�X;��=Z2>b��>bu>��m>�'>��$>�2>L���*�g����|�}�F�N��/06�fk���r���ln����&i�]{��W�S�ҋ��ѩ���"��J��=iz�DO>�r4?o�?$4�>�
�>76�>XXھ�b���9��sD3�*��t��/c�����Ȅ���ʾ����,>xnA���?�F��R��>�:�>��=��>�>�ט>g�=�>z>�}�>n[>���=z��>Jw>d)�>�ӼW�> ��=�̄��d���#4���,�����yE?N�g�N���	9�l�;�j���Č>�s?�R3>��*�#��G|��>y1�s�\���]�+�%���y>䂳>@�=$���mjB��{����)
�=�rc> � >�`B<�����`���=F��>"u־	J�=��w>[�(?x�v?�86?J �=�w�>��a>Ϗ>��=jwL>&(Q>U؈>��?��9?��1?|8�>((�=�n`���=�/;="�>�C�W�������&�#�<I2��(G=�dr=�<eg`=~yB=wXǼ`��;���<1J�>q�8?;_�>b��>��9�[�>�#>M��-��W>a����>qq�>�?���>+!�>�O4>0�b�T�þ2��5��>&iA>9E_� x�s��Pex>��r>{�O?�1?�h��Qc���<���=�u�>q�?�1)?�&�>�>�n���� ����K����=l-4�t[�*�����2�r��>�y2��!�8n�>G���7�>-��>��>7Ѥ=�`>���>���>�5,>t�C>lY�=
������=����M ��p_�{$�6����:U� c����:���#�l���3�n�=�i,?� �>������O㗾v��}��_
�>�a�>m�>c��>��"�}<ܾ�!9��%�\y]�y�>�R>?]�?����'a���ռy�Y&>�ٙ>�N�<+��=�L�>'��n<��?1�b?��>��ƾ�e{�Nڔ���i�K�>.w=CK���#�?!�Y?K�����6�,��y�>�R�`�s�=`8�V������c ��jZ����I���ҏ�z �>��;?��?����;u��^
�'R������wY��ak;�&���ף>e��=�þ�	���� �k}�����=�u?>�˜>�h��o�M?;�	?�!�=�Љ?�|O?F�?�v��1?��N��I=d!�>P?G L?.?����zf��+����=\��)��/��?�=�Z�=���=Zb�=h�Q>�>{�ã>�h=��i<�������J�=N!����ݘ�<���=9�H>"U?�rS?[i����Z���=���=:9��i��>MT=H��ǘ㾴�K>ݦ ?�
?��v?�˅>�=����iN�_�3JR>~I?5�4?���>I�$�&)o>�e¾����;$5=��>�:=ٴ���ɽ����+�}=�> 6�>���=ѵc>�_~?ЗB?�`"?׿���.�P�v�V�+��㷼������>�>�{�=4�۾��6��t���`��2��&?��DE���=e6�=c->UQD>F��=T�>%�=pݛ�Xؽ�o1<<��<�>�V�>�A?�7[>Ao�=����}���Z?���*-�h�o� 8���+���?X&?YO���Z?Z?�8K�a��}��m۽a��?���?���?�Gu�~:Խ_dc>�a�<\^�>�5>D__��ۡ��@����n5������� *����:mK>!��>E|����]��^x�>6�:�n���I��">J�㽷�o�K��<�þ�@��ѱ�����2��������@i��w���� �#�_�%׮�18��|祽Nל?�=_?I�|>_���|�����yܢ�M�>>�P	��Z�������)����0���Ͼ��(��_B�� >��ྪˢ>UgW��A��AI~�~C&�B���$)>E .?�䷾W򴾿��K�=�+;><��� ��X���e!��A\?I�6?M������a��� >��?^�>I�&>������a|>c�9?n4?�ŀ��	��3��Z���M�?�Ӿ?5iL?};&���Q�0�[�N��o�?�A%>��	?����f˾���� k7?t;�??v�>e룾�ܗ���9����<��L?T[�����>�U�>hU+>�_��\�`=ԡ�>ؽ�'����>��߽	I�S����->��>�U�>m�S>�p9��%�8��>�ƾ�L�Z�i�#���;��=��?j�p����<沇>��>�D-�S[��5䃿��὜�<?~u�?V�o?s��>���?��}�y���4�!>!�?��>�i��Zp?�?����l�3����?��?i��?=5?��}���ٿ�����׾��ܾ!�>���=�qL>H�m�G�<b�o=j4�:���y�=
��>���>��>v�m>W
>�C>�Y���h������ď��7�n��,��	b����m���'��njþ�"���Ǽ[��H��!�3��"�� C�v�о���>�8??x�
?o��>�I>\?>>Ω���޾<�J�Ɖ��e�D�{+���־�7�����R���-�� ʾhv>���:?ּ>��[=���>�;�?�~>s)c>�w~> 0>�^z>n̳=$��=���=��>>��=�r>ӳr=#B�>��= ���7҂��3��)���ϼ�Y<?�,Q������"7�^YԾ�C��Nݐ> '	?�>>k#�w��V|����>vc-�D�N��碽�ɼ���y>�̷>6> ��O}��
r��Y ��g=*�>��I>q�E=8���=���=��>Ԇ־e��=A<x>��(?Y�v?y�5?���=���>��`>F]�>���=@�K>��O>���>�?��9?�1?��>���=B�`�Fw=�<=�>���W�����޼��&���<s�0���H={�p=�j<��a=ԇD=���	ʧ;%�<�x�>��0?aݾ>��>D"K��h>�V�P��ҽk4>gЇ�j��>��>X�?6!�>�q�>�g�=��н������;f��>!�S>�se�H=x���f*k>�%�>JH?��7?ѐ���e�c�=ٱ[=���>�U?��'?���>3>�S������ʿ�G^���f�J��=���=�h�>�þ�퍾�2y��*�����nt:=)u�>��>G0�>Ar�> e>��6>`P�>1�9>m�=��W=�ݽC�l��e�<)=Q>DG���YԽN�Ͻ���~��=p#H�"���1��Vν�F�=��g=�	&?2+�="�f�%�l�+��M�1�c=�?j�?â?4a_?��>���0�I���h�zbʾ+/�>�JX?�Z?5�ǽM�$>N��T�=��]?�J?��b��ξ���=�Ծ�y����a>]�?�s�>����}^0���u�қ���>��=O��w�?ɐ�?�������;�I��[��FO����>��;qWU�k����� ���F��:ؾ�G��>��x>GF?�-�?$���52�����KX���Om���Խ�zT>�%���>Z?\G}��W���NZ�#D;���G��"*>��	?��V�J?�'? k?Fd}?"M?��>!י��fy>\�t�=�u�>JRI?�0/?��?Ħ�>�s�>�QT=^ڧ���þ4F��JCϻ$�콦�(>��=�s>�5��&��=��=
�=D�ݽR��<g�0������8=N�&����<شG>m?L5*?_˻������L�=���=#��Z�M>�H�=yQ��5�龉� >9|�>Q�?�Z?�w?}�q=���F*.����o�=f&�>��X?�1�>|k��h�=����P������i>O�!��YϾ�	��z�ƽy��<6�>9�?x��=��q>�hz?��;?�?��{+��y�Us.�_�;���>;=�>��=y�ྟ 5��q���`��0��䭼�eI�GT�<_��=t�'>�P>��=���==��<E|��e㽖7仳���z�>��>��?��g>Aϩ=4$���+��I?���(��!([�}e��Xl�;��=As>dG=���>���8�E�a�R�M�^g�>��?M7�?Q�g?Q߽w 1�ۺ�=��S>]�t�� p�t!��L!>^��=>���>�g=W�Ӿ�f=��>��=l�7�Sá���8:�澻�b�;�]���L���#9�ϋ�ʦF���i�&���7G��̾�z�̐���n��.D�
�,�)T��8���Ln��4�?�͋?���>>N�>#��˾��v�� ����Ͻ����M����ᾆX��|޾��Ⱦ?���A��O�Y�>�KY�ύ��}�u��a*��`��>*4?}ʻ����������=q>ϟ<u���U����5��\��a,Y?L9?!�۾���[Y�˛>�?L��>�}#>ăb������>,�:?��!?m@�����4���b���5U�?5��?�D?�罻t:���Rq'�J��>��l>�t>B�X=��ξj+�I�?��1?~�S>��	�N��/" �(�,>�0N?
UD��e>6�>�tc>XU=P���jϽ���*,��c�+>,D�����A�ζ��>��>j��>�[���#����>AK澙ON��LF�l�7�&�ٻ;ɨ?*{�#@�=�Hc>�q>��*��ߍ�r�������N?�?�R?|�7?`h���A�����=!�>6i�>���=\���>�>�|�>��mr��'��?���? O�?�DZ?B�m�zzԿXʦ���¾/ƾ��K>�>�kd>ex_���1=]#=��8=�>=�G>�m�>%�=L�J>��>K�'>S]*>ʼ��π!��Θ�����7�;�J��H����O�T�G$��[Y���^��Ե�FE���$���D�s����+��8뾩�=W�K?�I�>�͗>��><R�>���_K��j���.�@��c��y��ro7��d� �߾w~��;B�M1c>������>�݌>|w=V��>�SY�b3
>��=�l�5tA>k�<~�<�f��p�=�,3>j+_>��>�������>��>���9��,#?�ono��@���H?�l�n����r�Q������צ�>k	?�1>-Z2������^i�]l�>@��f�q�./����!=
�><��>�~�=34�;Ug"�u�b�0�<�`�;>��>u >ڳM<�q����A��є��J�>�dԾ7�=٭r>�|)?3�v?f7? ��=(��>�fl>�>���=nS>i]Z>#��>P�?��7?u/?xz�>��=`6_��=�S9=��7�*�?��Ӧ������#,� �T<H�<��5=��~=�o<e=b�D=W�����;ެ�<�/	?�@?�'�>� �>�圾��Q�\�d��"����=^����>�$�>T!�>Z��>B��>��>���j�������y�>��>�{�|���ɹa<�WX>�->�2X?�;?w^�󧍽4F>(�>ń�>�0�>��#?oH�>Q��=V�H�ݶ��� :,�/*?�t�����=���=�W�L]���&��&����8��+M/>#��>�a}>�>ՠ>w�>{>��>@.D>9j=3���]2�t
=��C<��=s[$=|R(�K�'�ϼ.["��,=>(h��V���ż��l��$<��?��?;��A�y=X��D���
�9�>/$>�?[q>ϝ~=<��0�O�q�����R�/I�>��B?�[?ߥ#��z>89Q�TF�]#\>ǯ�>�WP��;�`�����ߛ�>k�?�]G?���>U��mik�	��0:2�F�>R">	Z��R�?�ɍ?s�$���8�����XL�O*<��U�Qҍ������_�?�m��Ҿ��Ⱦ�L��=S�?P�?'���:�1=�оz���ң�i�#��>>Y ��<8�>�>rV�F��*���1����9�=�N�>^� ?�al=_��>+�>��z>�`e?ͅ?�O4?7{���>?��%?m F?�9?�)?y15?z��>��2>Y��=O�ýX��>Z���c��T����"�=wV�>�o�>_��>�m��&�<�Ľ�L�p� ��=�e�=�*���&>~�=���=�]�=��?�;?��I��cP��8�=���|e��3�>�2
>�%#=Q�ʼ��>���>�q?r5?���>q(���o����>���	��Q?�8?Z��>T�<�@�>�n�2�ǽ�G�>�Ck>�_��쫾�J߾B���B�|��>�+�>��?>��e>��~?1\A?�H ?a����.���v�x�*�,d����b��T�>�-�>9��=�پ�6�s��\a���1���C���E��B=���=�7>�uC>���=�>y=q<��mB�U!_<��i�]��>�	�>X ?jO]>��=*ͩ�l��wc?/�ʼ�YF��Q���d�	����Υ���.?��>�3>Y.*�P����8�K���>���?�l�?,�?�0�X��jt�=F3�=䴦=|M;�R�\}�=���=� ��ď>\��s������=l͢>��>��X����H����Te��,��\�A�;�[<��������� ��I�N��IS�a︾�N�����𞘾�{-�lS<��>������촾w�پf������?Fw�?@�>�'��B9�,�-�ӡ� �<!I��v��h;����M����ʾ����N���>��A�.Z�N̛>�JY��A����|���(��㐼A?>�9/?Bcƾx���Z����g=Wo%>�S�<�*�ެ������[*��_W?��9?�:쾥<��$z�G�>�?�w�>��%>G��v���6�>�C4?]�-?W~꼛��,3������`�?���?�??�H���B�[W	�Q��ֻ?ͣ	?��>�����˾d���?�F:?'�>��������%�li�>�zZ?�P��8a>��>`F�>��޽'�;,������_w�!�0>������`�(�9�Q�=(�>��x>�&_�r� /�>�⺾�9�M�3�
��S�� 	"��!?眾��nPJ>��(=�u?�qg�������-�=�c?�z�?{II?��,?c}Ծ�
���~�f>��>^b>�HO>B.*�:��>	��>��שa�����>A[�?�e�?�3i?V.���.Ͽ~?��E%�V0���%>�N>�qP> "��%>�G>>U�)>W=��^>�d�>���>� %>f*�=�~K>�Yc>"���X#��v��t���
�2��񾒫�� ��Ig��(�Ͻk2��"�ž���x���(��v�������~i�{`���~=?���>��/?�^�>o�>��/���F�k��p�!�?c��0�ݾ���у������׾��&��T>�����g>!Q=���<��z>�i1<^J�>�q>�tƼ	�>}д>g�S>$'C>}R�=��{>XM�>�X�>e��>!��>�P�=-��私�R7�d�b������wE?�7N�+Ӗ�@�*�ľ����N�>��
?E ->[�'����A�w�R��>$@0�9�I���ͽp�t�rc�>��>��j=���<nS��Zw�E�ݽ�`�=�>�0*>���<��¾'�ҽU<�D�>��ܾf�=�Tm>�g$?��r?�6?`S|=���>��P>�C�>���=4|\>�mj>��>^t?�0?�l'?%�>���=&�d�5ym=;m2=r�f��:��=�ܽ��Dw-�ǵ<�	���=�K�==T�<$D_==e㐻�$�<	T(=ͩ?��I?Dg�>@i�>���a�R���_�$}�=���=Kǳ����>M��>LG?��>�
�>�C;�V����˾Jd����>�1�>��a��dy�'�=�~O>k�.>�Y8?]+G?~ۣ�� �@$>)�>E��>7}?�1/?���>���=Ac��3��Meݿ͇W��Z?���!=��>��>>&����ӻ�n>G~&����_�m=@m>�(�>��>B�;=_>��V>6 �>���>�][>:�\>vk�=�GY=�,{��*���m��p��n-��3�fK���j�u5��p3�P'i�@���m��qD/?zb?��=[�)>� ���=�}���?27=���=����k�<��.�y��������(?��S?:�>
�pR
>=U��,�(�>3Sq>�Q�=���!�ʾ�3��^��b��>�v>?�a�>���<�������R[U�N��>�F>2j�Zѫ?�i�?z�C��������k /�f&�.���ᔾ$
��Ҿ�о�!7�ا׽.v�P�����>M�?K��? P3�Z��>���Z��_ॿr=��>t�&��>
�����'��h�R��$A�5Cx>s~><��>t��=�{�>�э>7o�>�]?
$?�J?7�L�L&�>��k>�!?o?$v&?d�?�k~>i�>	�>�⽠�>ʾ������:���t��`h�=U�>e��>�i��6:�<�/N�t�_=�2��{D�=�i#>ut�=���=,�=���=�u>��?��M?�# ��]?�pM?=s�~���̽�l\>ܘ�>�j><\!=��>�>�6'?Ml??6�I>'@�"��#�ݸ�� ��=5*?o�F?� ?�=>!Ǩ>�� �z,ս�ƈ>iX>��C��,�KX׾Q#r=�n�>���>>�w>�'u>���?gL9?/?w|�2�0��x��� ��e���J��>[R�>w��=�mѾ�11���v�~i_��J3�$�&��I��5=� �=��	>�N>SV�=`�>4i�<�4S��@νi�a<��z�>�J�>a�?�m>��=7����
���\?���U�s����҂�+�m����>��m>��>2)a���g�n`��tdk��뽞E�?B#�?�?�{¾�N����:>b�=MK�<�� ��ý���=�`彾�.>�>
~�� �ǽd�%�s=��>R��0����Vz�$�c���n^�2OŽ���	���t�'���fξ��ƾ�i&����hþ�b��������=�������l�ξ%ԇ��F�?�݆?��>���=�C����@4龤��=~c��;B������xw��K�ݾr׍��|վup޾@�+�\-3�z���Λ>jY�#8����|���(�0���5?>�?/?frƾMȴ�����h=#h%>�<�5�
���i���7��dW?Z�9?�"쾌=��.��-r>$�?LK�>��%>���X�>GD4?K�-?A>輜���3���x��B[�?D��?�0A?)��RIE����$���>bS�>���>&Ȅ�xRƾH���?��??Փ�>:M���*��N��ۉ�>�Q?��W���l>T�>Y��>j���ט���+u�����v��<aA>�Rb�h���74��� ���>E�>�.t>u9t��bҾ��>Ō��d�W�����E˴��Bi=6�>�!�׿>-�>8E >�/�K3��O�v��齟�W?L��?� I?�I?L���Χ �Q'��谖7��=A;>YD�<�9��B�>�n�>�L ��ӆ������?e��?�+�?P�F?��}��Ϳ$���L��bخ�x�[>�">���>��-�=�>�|�=�?�=�M>̑�>�:=>|�F>�F>lF;>L�#>�p����#��V��ϣ��l�$�7:
����d�Z�.n�ː��$^��
��$��Vp�}H��ѳ�h%�h��"�2���%Pý�^7?�?��?f��>��>�Ŏ�V.ݾ�`Z������E񞾤�գ�c���R���Ҿ,^��r�=q�/�b?���=Bʅ:���>v�^=N��=vc>�G=W¼��4>��=%��>寃>�!>�+>��>'w�>wN�>�Q===χ�u����n3�Ka��'�I��E?7(C=D���*������þ�y�>��?���>fO�v���=�?����>�����"����u�,>uN�>!��>�M:>s�=6�
�����[~v=m΅>��>�`�>%Fu=9�Ǿ�g���]>L��>ǰؾ���=�?y>�Q(?�Zw? �6?�u�=c��>9-a>-�>���=y�M>�P>���>��?��8?}1?r��>�?�=w'_���=W?=ޝ>��HS�`ڱ��'���{7����<>5*��.L=I:x=�v�;�Aa=�EI=Bt��2<�Q=-7�>�I8?@�>k��>��D���>��J�e��h�	>�G	����>�X�>4��>���>@p�>�%:>9�׼N6��]�⾼S�>ZC>n�b��kz�Mw^��O^>4`>w�N?�b3?sq{�c�\�"J�<�T�=�;�>] ?��(?w��>'2>����n��Z�Ͽ��$�[�"��s�;��;�m�=O�=��.���N�=��j
�<���=Rc">p�,>��:>u�(>U	>�/�=H��>�Z>��=��=gC��Z��(�����<�t8������罘���ɼ�;�������EE��������np��P�?��??G����:��H���7�ศ���?%�>�/?Ti,?�[�>IE��=�D��'�)˂��E�>��f?M��>9mB���=����U���X�<�F@>�<�>��s>������=�>�3?��6?� �>��վ��}�v�x���޾Z͍>!�U<ሾ˞�?�-o?
��!����ܾ)I�5�'���=��F�����{��v�%60�{���޾������V>��?��?������=�W��pj��;C����پFҽӉ`=���>>�
>�o��ߏ��ߚ��W"�@�3=/�>��P>i�=��>��?�n?j�b?�^?w�?�)���?{��=��>$b�>�?�
?���>�a>���>��=� /�2��(Ɋ��x<0Y���*�=z7>��'>+d^<��!=��5=	�<s%>�o)��:�<iu5<��=훉=���=p>��#?�B?)p�	��������|P��4>��>鱑�U�
������:>tK?��m?��'?S��
� ���I��s��;!>#�?gM?9F�>���<��.>z�,žC�`>.P�>�Z�=|o=��w�P��֌��kٙ>��>+(K�g>��~?�?B?O�!?� ��P�.��w�-+��i����3����>�y�>2�=�T۾��6�,Os���`�&l1�o5<�b�F��6 =Z�=Dl>�@>���=|�>�=\8���ٽ��0<U����D�>���>N)?_\>���=����%�Q�G?�~5���$�ت����C��J6��ѝ:=i��W4�>��L����~��'K-����>ͳ?YG�?�$a?m,��oj��>~�[�(1p��Y���;��.��1�=CQ�>��ս�y�����9�+� 0�>T�>O�=GԾ+��o����ÿ��E�����л��Tޅ�y����
�Є<�!7���y�<�1f��*��yiH��d���v��m����Ⱦ����?�2�?\k�>�>�|ξiy���;���"��+����ٟ���3Oݾ��ɾ:�ž��������-�B&7�5B����>c�Y��%��G�|�5�(�8�����?>$A/?�<ƾbx��7��1�i=��%>4��<o;ﾛ�������B�
��]W?��9?�'쾀���ὦ|>��?`��>��%>�:��Ȏ�'(�>P;4?��-?�m����(��ާ��0`�?��?��>?e����C� �� �g����>�Q?Jd?4i�g���Dn�5??�C?aS�>(���,����$��Y�>��W?��U�"�]>F��>s�>���Qke��x*<�C��+%
<�I>�V���nx:���� ��=���>��V>�7u����q��>�S��7���B��]�Hg�IV�<1��>������=��8>���=�52��!�����1�����Q?h�?��L?��C?	���)i��
����="�n>�JR>��H=�z+���q>J�>p5��
w��\��?o��?'x�?�'G?��u�f�Կ;��T��������j�=~�K>�~>��#�U�p>|^=>f�==(�q=�.�=��n>\V^>dK�>��9>�F^>,�2>=�����*�����hb�%j��	 C��X��ic��o*���{�࠾$Y���������H��>5��^$;FԻ��缛�B	?��B? z�>���>�=hʐ�Q'$�%���a���D�.
վ�8����5��:5���b������`��=
����?�S:��`2����>f�=u{>�6�=A۫���Ͻ�>��>k>q��=�	'>6��;�g>��>��>B�8>��������v=E�h����ｸQ?�m�����(o<�ý;L ����k>�,? �>�&�H�����_����>��!�8���H���J�>D>���>��<vX�=��9�ZRȾ�)�<¢�>:8�>jhz>�8�������޽ ��=�=�>�׾n�=��{>$2'?5x?�6?U;�=V��>ua>K2�>԰�=ʊK>�K>��>HF?C'8?��.?��>��=�j^�=�&=�2=abL��v4�a���-���J�}�w<,>���G=r=^B3<�a=HmE=,�ۼ A�;�/=��><�8?d��>���>#5���<���M��@��>�E����>���>)�?3\�>��>(�8>a�=��¾S�ݾ=[�>�+H>�[�2�v�z����>#5m>|DP?d-0?A	�ȗf����<C��=�̠>��?{8*?���>�>Q�ɽ����ҿ$$�8��ٕ�mߡ=�y��M����A>i�X=��(����gk=U>	> )W>X>�K>Ѫ>7��=�j?Ap�=��=�,�>�.�=T�3<��<���=Ռ���^F�P2>�?��$l�������0��hV�������0�t#?.0?�S��z�k����k_�aC��f^4?<ː>�4?���>��>?���V���'���`���?�q9?H�>X�y[><
�����v?>a�o>��>Z%>�A>���JWZ>�?�.?�`�>���٤W�W��� d�2�'>�1=�/}����?�\>?Yw4���Ҽ�����?3�t��6��:��������;��'��$C��r�΂㾤 �"`c>ѿ ?���?m����+��������B������b'`�ṭ���>&-=�ȯ��
��x���O�f_�<'C�=�Z>�%�"Q�>�J?��>y�l?R�>\�a?� =��?���>��&?�?�Z}>:֡=7֌����;��y>�U��1� �s�=L��e�������{p=M��>Tg�>��彾���!W= �>%����&�;���<d^<��=��->���=׮>6�?+�F?ߝT�;Z���g�<��}�,����>�9%>����5e����=��=ĺ�>6?���>s�����l
�SX��ژ=l�3?�eU?
D?S������L�^�+��@I>��#>���qP�����z�������.�>�$>[�/<5[>t��?�O:?K�?K�<0�:�Fd�'/��Y�=Q=Tg�>?��>4�V=�!ھ/51�Jj�	>\�G�<������q��V�G#C>\T�>,`f>O/>R�>P��;��o�B@Z��ۡ=�Y�=9�>	��>��?�qT>Z�=��X���ɾ�Y?�ĽT������}��,L�k�Y�M"=����b�>��Ѿ3���Y+��W'��6?r��?g�?��?�qO��B=�f�>�U�G:��������W��^�>k��>P$>vߣ�u&��@8?��b�=\��>��=z%��N����˗�!�����j��ý���A{R�NC����ɾ�S��{1�#��6pr��{��?�i��8�/�8�xa���q�}L��I�ɾCc�?t%r?�65>{M�=!7��6�(﷾���=�#���Q���ڡ�{J��$]���O���!ξO����&�K�9�x���Q?�.�~=����t�T���о�w����>�}�Y���Vx��T)��1 ?��>8�>��L�?���w�,>-�?f�?��0}��{�����H>�@$?�u�>�P>�E�(�佷��>�7V?ׄ]?�v�>q��K�����н%��?�t�?�d?�8@�V�&F#���� A>:�>s�t>a���4��Z��9n?1��?ͷZ?A��@f��(I7���]?� �?�mX�)T >j�>��>��0�o5��5��W������>gy >9RH�u�������a=���>�q�>lf���ɸ�f�>�k �/5�Mo��$���ᑾ�M��
�>����ٙ=^
>��};��0��О��ꃿ��Z���e?�Ѽ?��6?�IT?n���Ae&���P��}>V 5>�k�>G#�>�ΐ=m��>�b?P�$}��َݾ��?���?��?T�n?nf_�:Gӿ�����������=
%�="�>>��޽�ɭ=%�K=�Ę�QW=���>}��>�o>;x>L�T>��<>��.>k�����#��ʤ�4ْ��[B�� ����vg��{	��y�����ȴ���K�������5Г�S�G�J��U>����dh|>Q�?�>�>w��>\1�>���>-�ؾ��	���#��F���!��C׾��=#�hPؾ񫡾o:��ܘ!�1p>��-�,��>�.>c;>=:�>�˽��<�=��>p�n=�cq>گ,>n�b>mMz>V�6>��=-[%>.d>�ψ>�ϣ=뷃�-����B�HR��c<�sE?ƍ ��yx��-�1�ܾ�~��3^�>��?�"M>Q�'�X<����m�O�>Z�$��v]��0ƽ*3��D�>���>�xn=��мB�����_��9ȽH<�=��>� >����������� ==&�>��־���=��v>��(?��v?$6?��=���>�Jb>g��>K��=��K>qQ>4�>R�?v�9?�z1?x��>��=A`�2=��:=&P>��uW��=���㼑�'���<��1�&�I=�
v=�<�`=A=naɼ爛;�s�<�?V�;?�>��>>�B�n�T��T�~��=�`>�.&>�{�>�e�>	I?e?�>�'�>I8==	�+�7ᴾ�˾j�>��>=v��j�y熾җ�>���>��??Ӱ=?�(̽I=2���&�-�>g�>;
?�x?�
�>�=��h���-Uӿ $�!�!�%f��M����;��<��M�S��&T-��O��ΐ�<"�\>��>�!p>m�D>��>�2>I"�>fXG>��=r
�=><�;��;��E�$M=U��N�><@Q��z���Ƽ7G���u��tmI���<����̽ؼ8�?��?�~�=���������F��Fh�>a\�>�Z?to�>l�">�`�1!N���3��Fg����> 6d?fw?��0�Z_9>����gu�$�3>��">7�=�.,>�(�=t�[�> ?I�4?V�>�H��<�~�R<�S#�A�>y�!�Q�˾,h�?�vx?�FA�4���Q��TQ��<�I��>�q�[�w���4�/�9������^e�l�>?�4?���?�d��U�>:��z���󌿊�a�:�=ɣ�=y*�>�I�����@����F<��4� �>ض�>���H��>�?�?h�d?��>-b!?<��6?m�>��&?z�?��2?���>�v@>u/���R�;��_�A�&�����{����{������>x�%>$e�>q�<5����K�t��!$�_~����s�����
����=��>�G0>��?�?�DN�N��q���������>.�>�e<�x�;�8f=��.>{�?��:?8��>�Gr<j*���so�Wo&�?�>�0?^�3?b%?����2o��=5׾/�龚�
��5�>�cT>-8����k�$�-2���"�>Ǳ>��S=*�	>���?Z0?�9?N���#/���o��j�	�>��F<�D�>I<�>>�n>�
:�`'��`���J�xT$�]J��E�����y�#��>���>AT�>��M>�&�=�"��礼q���H��e�O��>��>l��>��I>�9g+ʾ�L.���h?���D�Y���վ����R�7k1>�}�>��{=��?y�h��؉��۴��a�AH?&�?O �?V�R?�p>��t�T9>�3>����*籽O�=�g�=M�;�U�w>=4>�A��X?�����<-� ?z)	?��>G��3�2��;�=u���WS����2��Ɣ���ŷ���+-�2����W�r�޾�T�!�o��'�����i�J�D֐�˄��m,��H�?!�z?θ=y��Of2�� �-��V=�=q;����ҽ䙺��%3���Eg��6 ��1����**�aT&���>�Y�e@��.�|���(�,����?>�5/?^ƾ�˴�����g=g`%>��<�5�˭������"�eaW?}�9?�L�k'����[�>��?Kr�>��%>�)��GI��)�>�94?��-?|m켣���9������k�?���?��>?��0�� C���
���(�@��>g�	? �>64~�~�þ$½�??�9?*s�>e��w���j����>)�U?g�[��(g>��>l�>���ĉ�� ��Ƙ��4��q�>��������Yj�Ke6���=�T�>��{>|Y��=���0�>�˻��A��3��1���T���)>h%?:%徼Ӂ>�>mh�=��-�fŖ�S�s���;�/OW?�r�?8�<?G�+?��s-־"���i�=�>g��>��=�c=�H.�>�i?�ߵ��`b��� ?���?b�?���?��R�}Zֿ`����R���m�[�k=�=V�=�kd���F>�j>�S�<��=V�1>�:�>2Lk>�e=7��=<V>�>&�����$�p堿�ݖ�YD1�o����"�^B���蘾�M���d˾�����U+<�Ev�G\�,h�Xu����<r������c�N?�5�>	 ?��>��� �J�k�޾�4T������g��:п�����+��S��_꙾�æ�B��;@c>?ھ�`?w鄽�x���/R>��)>ZS>��>?�\>��=���^�=U�D>��~>ؕq>%2>]Į>W�>�>G�,=���䅿�9N��o��\�=w�G?K���K��[G;�H�龚�����>�Z?��t>!�����E�i��.�>��维�J�)���� ��R>��>i��=���F�	=���<�e/�<p�2>V�=O�(=�mU��Q=����<��>��ɾdM�=��i>r�'?�:z?k�(?�>�v�>o�]>�̘>UD=:��='/�=�N>��?6�C?ν;?�E�>I��=]�U�q)�<^xy=��D�����
��������1�~8��o���x<h�6=�x�=�7='ޏ=��>�=����2;%�?`X�>:J=���>�[+�5ѓ������b)���|�0C���F=��;?#��?�yZ??��>F�=T��M�t������>��B>	�V�J,i�����ɫ >�(�>;u?��?���C��:��>Q�>�>�@�>,�>_�N>�4�>����
�ۘ����!��B�K����D���#���t���pj>��<>鈵�k�;Ym=͋�>3
4>W�><"3��p)�=*�_>��>S	�=A�>��V>�b<�D<+�"��[�=e���=�����=D-��u���ch潝�;�����+�#���X�c�?М?I��O^�<��Y�5#�{x'��h�>"m�>��>�c?ft��)
�ȊD����j���~J�>\�Q?H�>�����\>y�<r;>nD�>�W�>_��=�j)���pm���>y��>��?��a>3}�no�=6���,�Y $>j5=������?�~*?�\�2�@���Q��&P��pM�����B۾����r	\��v��%i���z��I���� *>t�?��?�?��h=>�о-��V�����:���e<�6�>�>�U>2 >������W������I>����o-?a"�>�'�>9uU?=��>);?�^G��p�>��j>Bp�>��?�e>)�>�?:>8Ǽ�u�/��� S>a���ݾ:�*�E�1�D�>�n=^�=��<�Ƽ(��=F%��!��>*P�=9`i>lFӼ����h�=Z�=/�>$?%?�}�8/�=�y<z��W�>��=	e�;����I&5��_���?����>�?+�?��!>E���6V��e�O�>��>��q?�E?p��>TB��.���`戾�Il>��,>8�L��2�K��&44>D0�=I� =�">�.�?��!?"�O?��n;n�پD�b�m^�*�=a|2���?�>#��=��]V��{��y�y�\�"{�V���88>a8>y=�<�r>�B>�Q�=���:�m<��꽣�Z���ý�s�>*3>���>X)N>
�[=w��������f?�ϖ��(�Р���c¾��&<i:�>d�?kGC>LE�>W�d>@�p�-���F	T�0��>�r�?�K�?j>�?#�����ج8>��/>7��=2O=;Ћb��X�HH�<CF->�
�=$�<���Q�\���%>D�>�KD=9���?���i�r����	�e�?hO=����[�!��G��;�\�-t��ـ�=AY��*	=�&\�I��4����O���>Ǿ3�����%��ܖ?�e&?�q?$�=�꾗����Ӿ�,>�P�Uv������������ �]Q�Q����ھ�@�о7ͦ>s�d�4��h�v�\�'��G���^>Z"?݈ݾ�7�{S�f>J]z>[��="ʾ�������#꾽exT?h6?h��V�����9��o�=;�?	��>�dd>�{��Y����>��?&�?����w��EB����;�?!�?-7�?MHF?������Y�1=]��O���>/4?D��>Lsѽ��+��y��%c�>U�L?}j?_�zu�Ӫ!�]�>g�o?�:4��E>�r�>f�=�����7���>�!.9̭>�w?
-��Q�#�����1f>y,?�j>�2�鑩����>3b���N�s�H�G�����DP�<�x?1���J>��h>;>:�(����ɉ�w3�H�L? ��?�~S?�w8?K3���������3�=r��>��>X2�=.��Ǟ>e��>	��ter���Ť?J�?���?�QZ?��m�~aϿ`6������ ����V">L��=:V_>=%���4�=L��=��<V��̼>�>�j>��Y>�s>�8><2>�݅���(����������I����c	�A�f����YW�?:��྾��������2Щ�e��'�3�c��f_>�G�޾�|���Y?K��>�^	?z?^�	�>���+��މ�M��]*����� ����𾐕�����%�B��Lf�W� >�a�����>��(>ȄB>��>׽h�A��=��='�=��>
�h����1�=��7>WL�>�\>[��>�<=Ϡ�>\b`>DL�����":P�`�:��=`� R?("�&6��� ��Ǿ5�M�i�>���>��=�8����C2�����>�=��eh����;��LF>W��>���[�=��[��c����=�%�>Z�/>@��=�X���6��#�y�>��ѾE��=w�c>	++?�q?�o?i]�<Y��>��d>/�p>�\=K�D>a0�>��>�% ?F�7?gi ?���>��=d�f��&=�:{Xn��ܽ(�<�>k=�"�z��<Q���iE=���y���Q=���=�j<ޮA<|^<��
?-�?!��>�;�>#P9:��"�v�#{��!�*���̽6��>��0>��>C�-?C�?�O�>�K<^�ľ����Ը�>G
]>:�O��
\�G���f&�>l�X>�O??C�?8C�2�!�'�a=!�5>v�?�4?0�?�ݜ>F�=�^�;Ұ	�u�ſ�W�qH;���;��T=LH�=|,:��/���<k��|���	=��s>�H<>�>n�>zY�>Fe�>Eq�>47'>(OU>7�p��8�=+�^=��><$��=I���M�0X��/=^�Y�:�@T�����Q����,�<�s=m"'?C�?�D�t7�=m��V�4�A-�'�?���>��>)6?��D<��}Y��Q`�����K��>�Ԉ?��?D�`���	>�����v}�;q�0>Q��Y��>��C��5	>-M�>�(?1[?���>��>���c��i���f)��|>��{=�ٔ�e �?��c?�������}�(���J��v�Y�E<qGD�K������	)�o������F���*��,�=n&?���?La��(_p�����:��B��$����k��~u�u��>�Ř�	ٽW�������tؽ���=�#� E�>諁�I��>�u�>o�?[~6?���>o�??D����g?��>o�B>E�2?��5?���>�?OC>xs�=�o9�Q�=����޾n�Y����7�b>��9>�>Ba=X��=���=b�ݽ{��Ķ���U	�YU�=2p>��=Fk
>?_�>G�>G9?�lr�ͯ��?��:,¾�(>��=}t>��E���>�I�=�:�>ܬ!?p�?���>�V����bE����SW6�?R?!C5?�D�>ʔ�;(�>�վ��=,=����r>ݠ>���������И��u�>���>�>�.b>��?*�??3�!?��1�.��]r��;)���� ��>�n�>�[�=�-׾ڄ5�Vdq��`��j1�Aj|��"N�nI=���=�>|�M>nj�=�#>b�==Yf��̽:�r�8g��	�>1��>� 	?��T>�x�=戥��  ���J?ᗕ��!�%/�����Xh��:�;�;N�j����$%=ύ��@���x��������>.��?���?��J?��s��gG�_��>G��=��>��������ڀ=$��N�=�G����/�����w�]޼�����~��Uc������?Q;�V��%�Z��A�<�
������.���Y��IG�����=�ѽ������EVf��� wM�3��G,���]d��X��s�?�E?,��>7��=e�1 �D�����<]1��"�Ľ�����7L���¾4�ھcƳ��� �)PB�`A��,����>Y�Y�!A����|�'�(�����?>�5/?7_ƾ'ϴ����g=Dc%>0��<�:����𯚿|�ebW?6�9?RR쾏*������>��?�s�>��%>y(���5�I&�>X94?4�-?'M켈���9��ܙ���l�?Z�?�D?Ɠ�e�Mx��x��='�>{�>�3?G%����s��X�=(�? :8?�ҩ>��l���$S�LA�>�a@?�x���h�>���>�,f>�E"����R1 ��M��LV�<��K`����DB��7�v>���>�k|>8)ݾ����>�v���N���H����%~�}F�<�?��oO>��h>�*>��(����ǉ��X�D�L?J��?{nS?Ww8?�1������Ӧ��i�=.ɦ>���>?��=���]��>V��>|�辙mr�����?iF�?Y��?�bZ?�tm��ѿxd��}�ʾ¬Ѿ�R�=L��='N�>r��<x��=�,d>�p=�5=Oc=�BD>F�%>O�O>7]J>��4>��9>�����%�h���K㓿4�5�v������eJ�8ܾK���A��\n��Vľ0�󽏌���D�MyνH�%���a����"��g?�t�>@��>��>%P>��I���F>�Y�ܑ��>�
��V۾�۾���Ka�����=)>����?� >
9>�" ?Ն=ǊV>W�S>�P����=���=�Q;=0�N>�\>O�>)�>D۝>��<>:r�>9�=���X�y�O/<��j�t��</@?�YZ�{��j5*�Bw߾N%�����>#?<zV>E�%�'T���-v�gM�>�&�R��,ǽ;0�1^~>0;�>:��=Lɹ�b� ��!���I�L�=�ԁ>[>�*<�l����g
=���>
�����=
@r��a=?�m�?�?�>M7�>�)R>G7W>H�>^��>/.	>)L�>;c�>9�=?�?�D?|y�=��U�$P�<�5-���+���i<�;����������=i:���>%�{=d�*�Q_<B��<Oio�QȺ�0��=�P-?.^?d�.><�>�@1�"�'����>���u�^S��Y>[��:6?@d{?ٟQ?�A�>�����`��*K�=�N�>�g�>JU� �Y��T����<��>�vO?=�?�Gw���p�������O=E��>+L
?�@?xɚ>�_p=9�N�����+˿�&�L)R��H�;�7���a�g��=�4>6�>��л�6�=}rO=I��=�5>.>�:>z�=^6(>�_�>�G+>"�1>��=s_?=%g>�<^�M���WٽCo#>#}�k4�F-��H*��޽��������{��4M)?y�0?��P���l>e7�s�=�2ŀ��l�>��?2-?�,?b�����*w���x�������=[1�?|-�>nU�\,b>Z���-�ٽ�Ö>�H�=��=�	>��>�P��P�>��?[�.?#P�>[=3�̥d�{z����?��
�>��>�����?iWm?���P��*��M�=P,�J@� �Y��~��� ��J �M	�����FF-�=?I��?�9�3S�=-ؾ��Ж�"g+� y���ȸ�v۸>����;�=�=jM8��҉��ދ���=��>�Ó���>���>I-�>�)g? ?��>��8=f�!?߉C�7�=�?�H?6Ɩ>�ׇ>��>�-�>��w>(�>�1���8���	<��;��h�=O��=���=z��<��G�0�=S�I��f�=� K=�mZ���6=���=Y�=�g���	�=��?��L?\s�����="*��GB꾵��>�0�>��>��%��M�=��S�[�A>t�?A%?e��>��2>?���&����Of=o<?WE?�u'?�hD>Դ�=���(�G��n4>�'�rԽ�b d���þ}f���������>]��>���=��>E�?Ǐ?��'?r�o��TA�a[Z��J�S,J=].��$&?��>��=�GԾ:�?�Ƴz�'}}�X]@�ן��JuS�;��=��=\S.>��>�u�=�|>{. =c9Խ� ��1G���E�=���>�h ?_?��>�1>�Lھ�v�!�e?��C��!�d�9����w�O����=�׽Q]̾bH>���t��ba��w��0�>��?J��?%>?c����<�A��>��>�r�>�����a��:�=�9����>���<�p�<-�]� �a��t�2$����߾����/!�<�#8��:��;�Q�DB�@� �'.3���D�t:�����&t���[�=�!ľ^�����++i�dGi�
��oWؾ)����z���9�?���?ZA�>���=���>�����K_ҽ[T����O�����3r������1���`��W8��/�`�$����>v�Y�A��G�|���(����Q|?>4/?�aƾ!д�9��(�g={d%>��<�8�����ԯ����~cW?J�9?�P�[+����<�>��?t�>��%>�'��j8�&�>�84?O�-?�4�?���9������l�?C�?�A?&p,�o\G��e �q�+����>�<?X��>�G����ھ"$��Vl?��6?uϻ>h~�ք��j ����>>�R?�aT�cVj>l�>��>`����������@��ɖ��V%>�۩��� ga����b��=N�>#/�>eJc��j��&��>�A꾍�N��H�������Q�<�?��5>Ii>�A>4�(�����ω��*���L?�?`�S?.l8?5^�� ��9���闐=���>�Ҭ>~��=����>���>�f较xr����?�J�?���?�[Z?�m��zϿ�픿�#��aR��I�=	:t<U�c>�=�
�ڼÎ�>{��=*j�=F(>9�B>��>�Q>�UT>�>�A�>�����)�Z����J��{X�D�=���?nw��t���ټv�hh��-X�� C���߽Ë���j���-�5V�)W���qH���Q?_��>��?L�>S�>@���0��֊�����F�˾�S�w��C�Ⱦu������P����K̾���=]������>�Ȁ=�~>��?$5���== �>�5Y=طj��L2��:>�~>��>ؼ5>5o >i��>�8=aM�>�e�=}.���<�j�>�S�M�X5�<�|N?~eJ��'��M�$�׾�h�����>T�?�6>>��*��&��#B���i�>�y��t�e;ֽc\�S>\a�>���="�"=]ʪ�(Cs�Q�edK=B�|>��4>g�)=��M�<�
���w=�
�>$�;½�=E^�>%S$?l8t?��8?2-�=&:�>��C>��>��=�eI>�^;>$w>�?�=?��8?��>+�=R�c���~=��=�QL�+�w��X��őN�����O�<�k<��%�=3^�=�/��z"�<��<��;��C'<�;$=s�"?���>�>髹=5�+�����삿r���/���y��;��7>�}J=��?R�f?��?�>>����Ծ����~n�>*�>Ka��-��B��f��>a��>�d]?=J?0���R�GH�����z�?�O?�H1?G��>�����#��������],�׬¾
Q=��$����'*�҃����M>K�ڽ�0>{��=���<�a>��Z>���=}���F1>,��>��>c��=� >N�=>�Uk<����"��=�V�=�ܽ�&�����=�}����/��zѼ�����⽏�F�_Aнe�$?%?���= >>j���@���<Gp�>�%�>��>�?��=�󺾵^��x��=b����>��?c/?A����>s� ��w۽�Ƕ=R��;�I�)Yi>琘��]�=e��>;H�>=�:?�)�>��d�L\������H����i>���=W���V�?�j?�k���z�=U�@�d�g��4��-R=/���������s�%����o�or��h�=��?]=�?�
���;�=�ݾ�헿Z��>��œ��!�����>��ܼ�Cv��m�cc��[�0�ɓ���a�=>@�>t\��C?��>�*�>oV?7�:?o��>�ˤ�,?���v��>�"?:H=?R�>遈>��a<.��=֚ʼ� ��-��AƳ��>B�<���P>��s>M[=f���_��H��=o	�=$O>qr�;����k��<0�==[��<�&��zG=>�G	?�T?�ȶ����<5�:�D����Q?=���>Ǫ> ����!N>���<��>9�?�q�>m�>̲�V���e�������g>���>�:?�F?��];���=Y�#N��mJ���q>օٽ9���!쾛���z�Z�Ji�>Z�>��>2�c>��?'�7?0�!?/���;1,�el��{ �(�J9a⠼'l�>1Ϡ>��=�qϾ�{5�-q���^���)�\K�4�\���<�N�=:�>,�V>�O>�|>��<���������4��H���>��>aJ	?lW>z�@=]������&G`?�,#��;���/���)�-8꽒�>���>>* >�k>y�������H����j��g�9?��?���?�>?�*7��ﺽ��|>L�d>81?��=[<�p�;>�Ă��'>v�3�!�=�	>/�#��Z�֝�~,;������h�=����.���̉X�
�P��3���K����ω��5��}�)��鎸�g=.;��訾hp�T,x�������bq��X��?�G?���>^��DC��5��G��#�U=UWݾ����N�k��Rоx��������-�+.��X3�|'��#��>�Y�HA���|�g�(�]�����?>6/?k`ƾϴ�-��a�g=�b%>e��<�;�Y���"���r��bW?��9?ZQ�s+��}���>�?Rt�>��%>�(��?7�{'�>&94?p�-?�C����):������(m�?G�?�A?>]+���A��Z�F+9�E�>��?��>n̅�DS��,u���	?�d@?f*�>�x������%����>��J?�-L��Kt>N��>?ʏ>fƽU�m���=��m���ڭ��>k��l#�S� +�h��=H�>��x>򊀾��о4��>8B꾻�N�W�H�%������K�<݅?��p2>^i>�@>Ի(����rω��*���L?ƚ�?@�S?�k8?�[��l��ꪧ���=���>bҬ>6��=����>3��>�e��wr�C�n�?.J�?��?�[Z?K�m��ͿJ���~������x0>c1�=d��>D����;�=���=�l����=|?>�>�Gi>9�P>�;>0�+>�9$>����(������#G�q��S�
�����s���S�r��_��MY��#k���"���ý�Qh���Lu�$;������!F?9z�=lW"?Y��>��m���0�#Z�2�N�3.���վ��yM2���2뾦9��ş�����R��;��%���?��,=ҟ>t1�>��Y>`�=4��>�z>���>��8>��>��y>�##>K5r>���>fn�>۳S<���>���=�Z���l��h(�2j���\[�(,?�?5�������B���!������>~$B?.�>���H���'<��O��>�<	h��q����;y�w>���>J`>�z�=�r��*��L���ֽ��><��=�V�<��.��<\����<] �>A��A6�>0�C>d�9?���?�+(?���=`��>�^�>��p>p�	>+�I>���=�W>��>ט-?�--?d��>J�>��]�Dc�=�J�=�ws��
�:Aj�D����V��g�����<���=��<�Ҥ���= �h=y�k��j=R��;}?��?�">A��>����-��Ld�A��F�"�v���o>�->�Ժ>b:?��#?�J�>��*�8���z�2��>Ls�>�b�븓�r��@�����>�i?q�H?xzǺ�̬�Q1;���u=��>a>$?�D?��>g�j]>�����̿�,����q%=��r=��=�s��6�=�s=�
�n�>)ry���/>D׈>:�>>�.>�>=R�=�z�>�F>?>S�=�j�<���=����Y�a����)����Qϸ�u�[�ҽ\��������,i���N� r?�?Z����S>�Uݾ��[L�=v�~><Ul>�	?�>K��=k=��	[S��Lj�B����>��?��?��K��aּ�ve�Wfb��K��5�<)�Z=_X�>��Z���+>�u�>��>��J?7~�>BT'�	_W�?���h�t�>�f	=�������?��m?C���F=�.��5Y�!Z)�ǹ�e6%��	��Ə���| ��_���վ3�˾Gͼ�Eػ�n?jK�?s��Ň>V������D������jr��!�H��>.	/�����ݐo�f�f���)��)<?9߻T�W>�.��'`�>�
?@�?C?��?��A?� ���V?!�">U8�>?m�>_xC?�R?��>�>�JO>t�O=�s��
yU�������M=p��)L>���>�^>���@�Ե�i1ɽ�Q=�y��&���l�=�&�=��ü�m�=�>�?�]:?�t��Omȼ�:�˜ӾM:�=��>�1�>�^��k�0>��J�y��=��	?���>r��>sK�>����CU���S��d�=$0?8F?pX�>��">�J�><�ȁ5��<L5�=Rv<>�8���]�r+��ͥ�XE�>�\�>��;=5d>�2?�n=?�"?����/�qn��%�
Z�l�><�W�>��>���=�Ҿ{�6�i�q���]�[[/�[]M�=wS�;�=���=��>��H>u�=� >��=����������޻�l��aܴ>�"�>�?�Z>$^k={B��s��RI?iך�M��9��ƾ��1�g� >�y>N�����>d���}��	���\6����>��?��?Δ_?�;�W#����j>��<>�>��I<]�F�u���g��{$5>�H�=�&s��_��n��;^�d>��z>Q����tľ�E߾�T*��G��r8W�\�ͼ��ܾ�7,��4'�Qx־5�o�e�:�)^����ӸW=y@���ۨ����~���[�Ӿ�	Ѿd;��!�?$�O?ز>�@��DE2�J����9�|^3>8�����a��xC��yľ����:����>���:�?����>��Y��:����|���(�J���
a?>`3/?�cƾ̴������g=[P%>7a�<B����h����9�QaW?��9?�^�0����X�>��?�m�>�%>�+���0��>�.4?\�-?�����j8��h����e�?���?L�I?@��gN� =���7�����>?A�?�H��)�U�+��=jW?a�U?p�>�?
����a6:���>	��>�/a��~�>;��>��Z>j��.3�o��:
��E��=�*9��<yܽ�g�l�:��>���>�ʩ>��|��f�f?�����^�{;C��E�HA
�5���?���;:�!=��>Sa���
2����x5���I�u�8?�b�? ٌ?��@?n�ɾn$Y�^lX�K���r��>&�>6zc>���=}�����>���g����d)�W�?�?62@���?U�o��Fӿ+�����������=�7�=��>>��޽��=�K=������<�D�>���>+o>�8x>˸T>Y�<>��.>t���a�#��ɤ��ؒ�[B����(���rg��|	��y�o���ȴ��ｾ��������ѓ���G�I��H`>�G4��}X�<�?���>cY�>�(�>x~E>)h��� ����#�����ݾR�þr~¾(տ��t���b��g��L����(>��E	?ݢ=)�=�l?7�>��D>�$��>��}>�U>�Z>�>J;)>݇>r��>l��=��{>!��=R$��z���t:���Q�l�;|�C?��]��N����3�+^߾����G�>��?�xS>ќ'�-���6y����>BG���b���˽�w�{T�> ��>�y�=�˻2u�P�w��b��=���>�X>�k�(���#V�EU�=��>��־x��=�Xw>~�(?y	w?�?6?ꨝ=c��>R�a>�ď>��=>L>�P>�>��?;�9?��1?a=�>C�=��`��5=B:=�>��W��Q��D�㼩U'�eU�<��1�\G=(�r=ۻ<gr`=��B=�AǼ���;���<���>�9?\�>�^�>_9���>��M�}����>�����>fL�>��?o�>���>�4>��c��þe��ؤ�>
�@><_�O�w�W���w>��s>�FO?��1?�g�v�b���<���=+�>1�?�r)?wM�>�>������tտ��*�2�/�7B>�z�=%<*>,����K��b{e��?[�n;��4?�=jY>$�p>g��>=�>�fM=i�>��?��[>��=&�>l�X�c=��������=��=���=Ȋ�=��\�H�5�ӽ��]�S�<�wQ�ň����#?�?	Hn���*��žW��h��E�+?�F�>PH�<��?��=#9�Zc���u�������>Fl%?�#?�ç��0=z�w=����1@�<G%�3����=�)�=��:���=i�7?�f?�?
�c�gƆ��R���%6��l�>�Oj=���P�?��:?8	��w���N;�1�)�3OC��w =��>=�(t�gT}����o�7�t�
���U�U���=�.?�j�?#��.�����Ѿ�v��$�v�������>��~>6��>~K뽾�Ծ"���{F�bξ�S�q�K>̵?J 3��e�>ASB?9��?�0�?5�>Z�d?�ҾqhO>��>0�>�-�>�{,?��0?���>�Ѳ>A�,>_�������%��������(=\=A|�>:��>H�M>�.�=�B�<(�Z��>�D������Y��0��wG>�`>D�?>�!^>���>��=?��=~A<!G�=ꭲ���<��0����=���>���YdY>۸�>��3?�EX?�`A>�3～��] ���rꊽ&��>ZGY?�?�%;
^�>�빾9�o��[�<� }>�� �#}��� ������=�6�>�0�>�5>�>�i�?�w"?���>���W��̅����Ǭ�=jBw>���Ɋ�>���>Jh�	< ��g����y��
=�wс�Q�۾��5>[�Y>k�\=Z]�>!�!>pyL>bݾ��1�ah�>-k��S�*�l��>�`*?3gB?n�>���=�G۾
�%�;�g?^�{��U\��<��S �bas>P7>Ui�>[�=C@='�C�M}���^��@u�.�?��?ȯ�?�̟?�3R�Nz~��*�=�fG>��=��=N����oսN���g*�T�Q�u��E<�z>�	
>��@�����B��J�����C�`���<��	g��������zV�������B�,m��2Gٽ#���"ʿ���%NE�ﰟ�Z뻾S\����?�"L?-.�>���=�7���ξS���%Z>Yݣ��C��Ç�h;���;�l����J��������(���4���{ٛ>ZMY��5����|�]�(��B��_2?>'Q/?	ƾܴ�|d��mh=�+%>}"�<�x�����������wW?#�9?�R쾶F��9M��>-�?�e�>�U&>�����(�%p�>KM4? �-?1�����_5��8F��Y�?���?��??�zN��sA����KX�.�?�y
?U�>Ě��o�̾;d��?J�9?�V�>���c���N��-�>x�[?�dP���c>R,�>�D�>`�뽣���~/2�5۔�7���<>z�Y�l�g�c���8��@�=8��>^�u>0(^�����H�#?���V���=D���d�O���%�ؾV?ln��vV>hp$?z�ھ�Ds���2����}���,?�?΅l?��
?�%�_����I=�-���>|�?e�`>����]v?:�!?�'�Bw,�Y�?!h�?���?��o?�;v�6�ۿ�;��(�����վ��=Q�=<bF>� ˽�)�<ZԼ��?��9��e >VL�>�Gy>�xx>��J>�v:>Z�:>0���Q���J���ݍ���>��P�x~��pb��b��o��q��*Ҿ����;
��b���~���0J���6���%hþ�<!<T?�%?S:>w�>�,]>�S�Ov)�>�k�'6���þE?������S��b�Ⱦ7������[���F�>po;��7�>�3�=��{��"?��<f��>E%?�Y��OC�:1�>/ g�g��7�M>��>Z%]>8�>�Y�>�"|>�0�=1�{���0:���Q���l;2=C?"^��a���4�O߾ǯ��Ey�>E�?�TR>�'�Z���Hy��]�>�H��#b�p�˽�0���>/
�>)	�=Fp�7�LIx����uw�=7�>��>*<h�tC��k��=:��>T`ʾT��=��o>;�$?�t?�;?0�=���>3�\>�>q�=PyE>�G>��>FR?R-<?�1?N��>�a�=�z�2��<nڌ��Q��#k�������E�`%"�hx�=	�q�d����=�4�<G&Z=�� =��Dg�r�ۻ�`�>el;?�s�>ٗ�>e:�w�<���O��S�y>Q���	��>h9�>�+?�	�>� �>�T&>M���@˾�D����>�8>�Y�}at���+�Rp>y>�cM?�\,?X���j�a2U</��=[ �>@F
?C�'?!�>�>0�ɽk��p�׿����2�ޤ��!���=�z�ˈ���R�7@����b�d�=ײ>���>�\>UcI>=w�=PU>���>�>�}s<�^>I]n�����3��c��="���">�K@=B\�>?�~=�ż���v��*�P9��,���'?��?Q���K���F�t����t�'�?5[�>�k�>5�>�gA=�����l�`k^�ʔ��>CPp?���>����[��>�e���FE�ԤI?���>
z��c����l�,��tv?���>i�S>�>ag�������L��>��=��ھ���?��x?֋�/�9���A�O|-����6���(��t6�߀��]� ��XB���C���ƾ���=?���?D�׾����D��ĿJA��-w`��ɻ%<<�?g�>c����B��|8�#e��˾���?�ރ�[��> �,?o�>GT8?��=?I-B?|�ӽ<(?t���ȓ=6N�>	�?��?v��>A�	?6>���=��>�V�lP��4�N�r�������=C��=�r�==�<#�J���=t,=������޻"ݰ��(�<H��3an=L�A>I��>�xM?/
_��m���l�>��c�(Da�z�����j��;1?����l ��?=>.�?d�}?�t�>o>ƭ/��t����#F��/�>�T?�q!?�>Z:�>�I���N�0��Q�_>�� ��Lx��f�����͐�<Da�>��>��$>\;�>��?l`?�v�>�7����!��:�)��~Ǽe֒;��<�[�>��=�s��󾧻s�_�}��!F�ܩ!�pKM�%��<�F�>�_=��(�SN3=u� >�e��>�U��n�>��q��� �(?�U?�&i??>4|K=�%򾮖4���h?Yӻ�c:��▾�h0�����XM>�@?���B?�E�>���/<��MQ��p�l=�t�?��?<q�?��w�r��g�>��g>��A>af\>�j�Qι�>F_��1�>�#=������h�=q&>�X�>\��=�2��`ܾ	���jU�䡺�]�X���{ꆾ��������j��Bہ�\����������7(�5�#�x�4���"�������y��ݠ�����c�?Ͱ�?F�>2K�>u��A������K���b�0�����{��%H���䎾������,��3�h<��9�>�*�aa����~���1��j��i���j1?L���Y!Ӿ�l��S��=��ƽ��� ��윿�d����'�n�?��U?�#����S��ޔ��~N�,ò>`��>(��>�7Խ�
�љ>;[?�*�>Ov���
��.���7=��?�? �??�L�/�A�A��es���?�l
?�*�>�4���v;�3���
?K�8?Y��>�&������g��>J�[?|�P�fIc>�\�>�O�>`���[���:-��-��{���ę:>�ƪ�n�f��I=�C�=��>�w>��`�\-���� ?�1m��#U���_�ĝ����0a��G�Q?�(���ֿ=���=�YV�!K�������㭽��Q?`��?gMJ?F?b����e�v����f>�>�*?�7>��r��ֻ>�9?����ޔ�<Ӿ�l,?�x�?��@GF�?����!�ӿ���ۉ��<���R�='�r=�R>8�s�����9<�H=#t�:�>
l�>��l>))�>��Q>�>��p>��� �
��8Ə�S�S���+�|��Zx��r��_3=���þt4�M��2g��4|=�)��?��ֽW���;�|�H�?�"?�@�;��J=ϸ<����-��t��� ɾw��&@վx�о\����/8��%+������N��xt:>�N1���
?���=,�C��q?9U�W%M>�_<>��)>�g�=��>d�>�w�<� �=�;�>W>6�>�Y4>���>n�>�}�ũ��K�;���L�ʳ�w�8?����M��"
3���ƾ2���8۝>#_?ls$>�.�����4����>E����/��d	��
�<��>�W�>�/�=*�ڽ0��<a����2��>!�f>8�3>jI=`I��.v�A���H�>kqվ���=,Jz>Wh)?�Rv?�l7?6�=�)�>�`>��>�v�=� P>�R>痈>�W?Zo7??�/?��>��=�a��<=�%=�r@�d�S��6���餼�8�l=4<�]�
�U=:�y=sI(;��V=!�5=d켃I�:>M=��>��A?n�>�ޯ>�U��w=���S�X���>�"z�O��>	��> ?D�?5�>��=��ʽ6Ծ���cy�>�N>$�J���~��ʹ�ˈ>���>IZP?<?}S����)!�@�=��>��?9�,?x�>�>�1�=*	���ѿ����������}=6���E1=/%���=ʰi��y�<�M>k��>�:P>-Y�=I�%>
l>t�>��i>��<�>Z�s�'���R�=���>��>"�==ש�{U�t�韘�r��Z����︽�}N����=�7?���>#.����ͽ+yо����᫾��5?��> '	?AD]?lO!>�ݾ��T�z��D�־��>m�Y?�m?'��x��>��2����<v��>�	c�L�sp��SE��8^s���<o?�?R?�_?����ᅿ1옿�tq��k�>��=J�Ⱦu��?t�9?ZT#� D%��Y��R�2q$��}Z�0���j��B
�v0�$uO�n��g=�}�;�	/>۵	?�f�?4�ӱ��R6�����O���H�aԼM]��Õg>o>?>~���q�l�8�jz�'�g�t��=���>�&����W>wZ5?M3?�M�?R:?�gS?�S/��?
�=dIV>�~�>4�?9�$?+O�>�`�=R7�;�'�<�Q>>�뽤;K��<��=�&�ڽV�>�J=�r�=��=��F���&>n��n]�;m����q�z�F=���<���=;�>���>/hf?�[��:yr���>���~�׽���O�ܾ�+?��
�ڑ<>v�>�_4?��O?t�o>50�i{"��)��x��[*��f�>v_�?WH?��M�q/�>�Ͼ�D^��҇>���<�u"�x�������w����`W�>[�>��->��>��?���>���>Ҧg���:��+4:���=S۞��?�i+?�(B>�@��#@�0B����v��VB���\�l���>Ҙ>]B��٠<ط>h�=*������&�A�@��$g���>=�,?�T?ٽ�>ǚ*=��о��M�:��?�Co�D����5ﾏ���#?��3>�3V>Z���@-�V���K9��@�̿]��zK�>���?T��?M�?Q�w�9����<��n>�&M>Q�L��E׽o�=Q/� j>��4>��=E~U���#>�:h=�|=�lZ��QǾ�e��:/1= ܷ��,_����*��l+������t�I �=�_����J�x־�ڽ�����j�o�P���>��Q�ɾ��$��g�?�x?{��>�>;sھ�!;���,V&�,�ƾ��_�oY��m��~&���T�ᵾ[_��Q�W{0�c�0��؛>{.Y��$��Q�|��(���!�=>�N/?��ƾ���_��d�h=�$>��<��ﾫ��������@�y�W?:?+o��%���X㽱[>��?z{�>k'>������e��>�4?��,?A��7��9��M���-|�?���?�??O�I�UB�,��\Q���?��	?���>�����/̾���.?��9?�>��VՅ����>�[?�"Q���g>�T�>2��>�.�:-���	8��)���%���K8>�S��=�<ne�)<�2�=9̠>��t>��a��䯾���>R���E�I F�k�����������3?m�
�_P�O��>ȓ�=�D�nף�8c������Q?�?�?ѧ6?��E?NZ^���^��딾��>h��>���>��>����r=h;�>�x �����G\ܾq.=?[��?���?Αn?fgz���ο{����.���mʾ@�(>�m�=B�k>������A>�8��q�<�@���>0W�>9_�>��f>���=I��=��=$������������;11�l�����ZO"��I�����0�!Ѿ��ƾs�4�+9_�HU�:�l�D8<��Ƚ.r���\9![?YD�>�0>%}�>2߾<g�þ	E�\������\�8�ľ!����$�Q��X#������E��:��=y�&��� ?i��;��3>���>R�8���=i�U>�~�=�^>�oN>�Q�;cN,>���=!�h>�.�=E7�=9-�=s�>8��=�����|��ߪ:���F��6e;�>?5�r�����5�2��6޾�h��ap�>^�
?,\X>p�'��_��bcy�WO�>*2U�>�c�5�Խo�߼�%�>�D�>|ל=
����4��jz�44�?ʿ=�y�>$�>��/��������i�=���>�S־���=�_x>��(?�Kw?;v6?��=�@�>�Ma>*��>#��=:uM>�R>��>w�?�9?�x1?���>�<�=��`�
|=ٽ4=��>��Q�LC��o�߼}**�L3�<��2���G=Q�s=~�<��_={�B=h3Ǽ��;�X=���>��9?�r�>j��>��:�>��{L�X���>����:�>���>1?ې�>�z�>�.>�/v�Z�ž��澵p�>�.@>��]�fw�t��wCw>��x>*�M?:�/?3Pc�$�d�}Q=V	�=��>�~?��(?@�>�n>�#��ŉ��uÿ�����$�%�=3�Խ��o�,��<f̭<�X�F������N/k=��Z>���>7%z>��I���q&�>�~�>�A>4�=�>Tэ�W����a�Ri�J������>�=ܽ72�=��9:�p�����Юֽ��ּ����)�>~Y"?Yf?.p��e�f�O��@��(̾'?K��>��>��>~��=p�������W� ]�[��>��n?8�*?�*����>]��=���=�p?D|�=��X�:�%�"|����y|���>�0?Ǽ1>4)�,"��T���8�zIz>>��=�6��Z��?�dU?�����6��G��;@��`�5��=�0l��p#�{�����>�Z��e�P��#����'>,A?�>�?A��A��_������O�s�Z`���>=ܝr����>Y�h>�MܾS����/����ߞ�[��>}�>�*=��>Q�Y?�-�?x��?o�>�rz?G��p,?|�>���>�c?��>?P�?ݽZ>̲p=(�>�'>�(i�H*�������=�]"���=7(�>0�>J�=o%=��7�rN=������?<e��7�;.�>�u�=���=�ȭ>l��>��M?@������=9��H�>rN��B���>�o�A�>�d�>?˵
?Y�>-��˰
��T���оϼ��>�S?�?����:�b>؋ؾ'�==��>`
����p�Z ��Q���Hڽ?h�>���>5�>|͝>��?-�	?s^�>50X�Z}6��p��f�3�,�pw�>p ?��>e
 >y�¾�k"��1~�f�f��L�,]�
T�%��=��k>wv��H<a��=�ͻ>W����ŝ�5�=��7=T��=J�'?�G?��?�X>��#��(þ��7��pu?8���j�t�%���,�##�>j��{���9�:>C�(��߾�˭�~���
K�@]A?�?v��?��h?�ϼ˾V��K�=���=�q#>��j�b�Ž��s=�F���	�>��<>J>�.���w.D=�2�=ZА= ��Mɉ��'���#>E�����K�}Խ��ܻ־��ȾO5��� �����M�o�־SsP������@��/э��í��ə�.���?2x?��9>�>�S(�U����<����
�p�H��
�5ra�)�~���L�%S��_(�w���t/���>�Y��@��g�|���(�Iˏ�ق?>K5/?4aƾ
δ�H��u�g=6b%>iı<a9�Ю������a�qcW?��9?O쾰)����,�>��?Bt�>R�%>�'���4��(�>�74?��-?�H����K:�������l�? �??�??��L���A�G�����QW?��
?E�>���j̾:���?h69?�E�>n]��w��yD���>A[?�lO�3:c>K5�>>�>v�⓾��1�OU�����zS;>��˻��&1g�`<�F �=zD�>?!v>"B_��{���v
?ϙ���Yv�;�J��nH���
�N��=6�j?��T�e�>X?�2>��T�nϙ��K�V��J?��?�g?��!?w����� ��f��z���ST�>��?��=�ᱽ��>A��>�T�|��M���>{�?_��?��?�5t��+Ͽ���*Ǿg���g�f>�9>A�J>&g^����=ׅ9�v������3�>�D�>h�K>���>�E>�,>q>�=�������tː��>� �1��` ��=�=�9���}�������f���HX���%|�� ���&�9���\��纾k�R�*?�>!j->"�>��T>�ue���b��a���q��Q���W�i� #����o�dx�B��ns�
:>����%?v�>>�����?�E��x>M��>�S'>RҮ>�%�>��E;��=��T>!��>�,>�>
�=&|>��=gꄿ��8:�� Q��u�;E�B?��_��ŗ��3�]�ݾۋ�����>0	?��R>��'�T˔��x��a�>r�G���a�0eʽ������>K3�>~��=�r����]sw�$D�W�=<��>`�>�+`�}A���c�Z�=�\�>�����>X{�>T?Z�?C�?��=��>{)">�#�>�	> @Z>T�O>V��>��?��?xd?S<�>��(>���ߢ�=�v�Ѓ/��Pܽ��	���8������=ʯ�<�H�<��>������9�z�<I'��	s<O��<1��>oe9?���>?��>�ND�qz?�h�N�`���L>���C~�>���>H?.N�>w��>��>!{���ež�վa��>>�H>��c�'�v��~&��&Z>�K�>��T?1�1?�葽��_���=��=_��> ��>��$?��>9�$>�	��U���w����������-Z>�	<7Rb>��~�F9�7y��+' ��Ծ��^>5³>��<�S�<ۄ�>��>�����>�1n>��>��<>1����=ŗϻ����V�=d&V��p���c�n�d�[�)��� ��zW��R��w=��=�1#?��7?�Xz�uy��� ����V*����>���>$W�=؜�>�X7��`3�� h�S�<����p>�#P?8-?��1��>� �=�+��$�>p��>9Y�����J
\�Z�I���4���>e!5?��>�mʼv:s�;u��fF:���>&��=-|�<��?MP?�%�10S�g�D�<�.����=�!>i���(�]V�	��������d������=�?)�?� $�F\f�o�־hZ���h����D�Q��<���=U��>c��>C�پ����2����g���|��=���>H�=W�>0�@?��t?��?}:
?�x(?�`��Q��>��A=Q�4>Z��><(?(�H?�*;?Ok�>��>�)]��Ԯ��u꽄�P�S��=���=v.B>~y�>Uc>�=ɣ4>� e��F9=��`�۽[0<uԸ=�^�=f��=��=�0}>f?,%4?x^[=����b�=�v:����=��q��š��ˊ>G'��Sh�>��>�Y?�`?�"�>Ԅ���M%���,�}���� ����> `?�?��:s;�O�#���i�V�b�=��d���>��r}������_�>v*�>��Q����>�H�?�?���>J������[Co��1���J���U>*O>t	�>����ӡ��ᾔco���v�Y�9����=��`�A\=��I>!>���=ڝ�=���>�uܽal�Y-"==�q=n�\><�>�	?d 4?�ה>�S�=dt龖D1��3[?��K���@�Lg��y��� �8�>�1�>��>	L?Ջp>��g�č���=_����=��?���?�͙?�[�9~$�&��>�V>�ߚ=?�q>��&���`�Y%Q���>��B�VӾ�Z�khW<�1C>�A�>�zͽ�H��M��h���,?���oP������ƾJđ������N��?�ݽx���(
�f����j��X��l�H�i�O�몏�Q���c�����?7�?�=���W�4��S�L��b�=�_��Z��������R�������������:w+�e-�5�9��>���������s���2�7���Y=!�7?��Y���) ����=歺=��^���BԔ�#������.i?��<?�žD'��e����=��>���>���>��C��>��q�>I�$?N�?����`������b6=�ع?�r�?	1B?��߽��6��T�X��U� ?���>��>`���8慾]����?HM)?
H�>���6���+90�6��>��o?*`l�:q>��>�W>Og�c\�c�=��׾J�
��p�>���i0�=Zq9�������>�(�>�5K>b���6ܾ���>�3ݾ����E;�^�+�F-�sTM��?`��SÐ<'�>�}=_�"�Fs�����Z�ɽ�M?���?a�@?��E?�z��"��l!��=˰.>N*j>v����u�1��=?��>t-��{m�ύ�@�/?Yt�?�?�_?էN�\�ʿ�P���믾贾�<>��=Z�o>D�����='��=�~��,=O�>$��>�K>�3X>��9><�O>!PC>�b���(��+��WĔ��Z>����A��i6����b��5[�Z���)ﱾ����Ͻ�]�������7�MY^�>bپiO2���?X��>Y��>���>X@=h�b<�3�b�J�\h��� � ž�!�Ⱦ��������U��ƣ�K{�<�x
���?��2�(T��$�>O��:sX>6�6>��5>���>�h>"��>n>��>�N>��e>QoK>6<��>�z�=ƶ���g����X��������>ꗯ����~�D��B �;���f��>��/?3K�>�Rﾄ����o+����>RZ���*��p��!{��E�>��>)���n>>�/�=�]���ҽ�!O>�Z?�G�=`�:�쾾�����>ee�> iھe��=q�\>��&?	x?'�.?pa�=K�>H+�>�آ>'t >��r>L�4>��t>��?�D4?K?1?���>��=�]���=��=�7��t���G��]ļG���d�<�&O�.�=�u}=��Ÿϲa=ƃ�=K'�<����l=P� ?��4?�D�>;_�>� ���B�E�O��.�kd�=�4m����>�>�?&?���>V�d>��	�E�ѾEFϾ�$�>�{A>��_�s�r����㠃>\u~>�:C?\�6?մ���k�po�<���=Y��>��?��?�N�>^>�2�Y) ��̿�ɾ,���E�ąS>+�P=.�)>��*=�N�=�V �q��+>n�<�׎=lW+>n�>�7T>���=vy�>v#�=M\�=Z�>MM�;��I=�ւ=)�<��:����i�tF�,:�
A�gzݽ�<h�o�}�
�it���?��?k���b�=�m��R	�o+��e�>(u�>���>L�>��=�?��]R��P>�r�[����>�Y?�
�>w>b�	�>�����<�ܲ>�8�>Hf8>U���`H��
�O�rΖ��x�>�Z?-g�>��a��Yf�J\��,���{>Ð4=�M9�瞤?x	7?�#���D������Cd��P�<mt���=��󇫾�/�&�>�0�����;��� p̻��?�N�?�꘾�%;�� �_{����~���ž#�"���ν�?�k�> ��V雾���ơ��n���	;>���>#�=��? ��>TY�>�o�?��?�V?�Z���?~��>h/?�I?���>�~>?P�=y9=������'>u!���W��2 ����=aw>ۛ�>!�=�O�>iq�>J��=5��=��0��q��v����w�<��u=;_>��2>9O=Lw>y�?Ud?Z뫾�Y+�����T��7��I,�;W�4>�[���=��@=��?�C@?I�?�Te>[  ��^����>�?�Dg?���>�����x>���� %��k?=�&�>L�>-��4_����HI�j��>���=�;&�e3f>��?w��>ܛ)?���6�J�����H'�G�<�y>�@�>��?V�+�7Už�J�B���b"o���0��ݾ���>��>�S��%F>�ƨ>�G"�F���s��=���B�p>ڪ�>��>B!�>���>W8�=D�G�\�޽B󚾗�L?(�b�Z���޽��ɾ`�������l�=�����\����$���d�����#��x ?:K�?���?��?n�(�|���|>��A�:k>��>���,��*��L�/>l�;>e<پ��P�"���&�>���>-�S�Ӿ�"�.(���ۮ�ko��j>' ��S���<�%��L��>�;&�{r<(�Ҿ����Th���w���yz��88���M�����ӷ����?��f?t��>�9�u�!�2�о�����L>���$���àp������|�W���)|�C�ھ�t����{g���>�;��c���`�����&��J-�=$�?�d������)�9�p��(q>��t>+�����o�C�������w?0�0?^�澋,¾h6��`��2?�	�>��>HS0�Zq˽k��>l�'?�94?Ջ����\o���l����?�
�?��a?�!���wW�Q�7�n;��r�?��'>���<�aU>N�."̾ �2>y^|?�|A?�׳=�`�}B�-�L?s=�?Y�����R>��]>�j=��+������ͼ�a�:������9�	��g������"W�=�8�>���>i���P�>&�Ծ_$�3�1���M��)N������\�>�	(�t���@�>�Qνu9��M���{�h�A8F?v�?�+`?��:?�_����� k��{=��=Z�f>)�'<�<����/<͑�>'���S�z��Ӿ	=9?S��? @v X?�̅��e߿����Ɏ�B���<�F=��=``���<��>��<�}ں��=lb�>��\>�wU>G�+>:��>��>���c)�?������0�����U�1�T�ۼ"�*��ռ��ceh��оդ�����U�����N������ʼ�9Ͼo�0���?���>M�>S��>���=�k����E�ɽ`ؾ�]���|����;�������%ig�E���sc�i�����>��c=��>��>2ﱽ�
�=��>�[�<�4�>C�&>��=a"D>��>M�8>�m%=-�>y��=%�>�t�=ӈ��t�д+�r�Z�u����=!?&hY��!���.4�o���y��9��>��?C�>��t��q�VY�>�����
~��4��3żuU�>��>�Q�<�1�=���7�,���"�m>���>#>�����������z�=���>�㹾�`�=i�^>�@?�g?yS9?��=��>k�j>�ڃ>�>���>d�q>f�n>�?�&?�2?���>M��=�tB��b ="9=}*K�X1���U����޻Kq�=�F�9sR�<�ƻ.A/��y=]7=4���k�;�N�
?��G?L>\��>�/L��Z5��?��HP�IA>.��=T?
�>9��>?�>wj>���;#�=�K���.�>���>�_�~��a�=b��>�9�>�?ԞL?��h��]��I��>x�>� ?�� ?և>];->x�)=�����տ���61��Z���
��0�Vh����ɽ
#�=y�!�W��;��<N
`>�ۀ>:jb>8>�->�IH>�6�>i�>��>d_�=��=�2w=��Ľ7�>�����Lq=�j��D@�Nv��B�M���#���7�󜂽4v� �?${?I
��I��=bHP�x(�X�����>%H�>���>�e> �=\,���P��-:�X�q�|�?�_?�޲>�vx���=!E�=�̩=a��>��>\���n�=ti<��=z�*�M~�>�)U?��>w���*�|�pɐ�Ko6�)x�>�Y��9��fc�?s.?>E �%���4p%���"�~l9�c��=���<7d��BGݾ��N���3�(��1,�aH���Jg>Z	?W�?qfվ`��=DD7��7���a����%�_��r0�|��>Y��|�����4���ImǾ[l�=W�[>G/�>���=]�K>���>T?��?_�>��8?�{�>��B??�F>�!w>�&?zRG?n�>���~��|.(<3�>}h>B�b�,I����$��,�<g��E��:&^�<t}:=��"<J��<#qC=0��<9���ӽ=DL=k�<�+�=��=5?�<��?�+!?�̾��ɽ��a<�r⼧��Y���t�>`��=,��^ě�F �<`f4?X�x?D� ?_�>�0��7���:ѾA})=l�?&�#?�l�>�Y�=��>>1������ �=M݁>�ὼ>�������k�����>׎�>��n�/ٍ>�j?D�?5�E?�鑽m�L��=�'������cS>%�>JI�>o��=�Q��Y)>��h���&N���+�3|��J�u�=��3<��M�wE�=�<>�$�=b������Z�==�>Fj> ŋ>�e�>�k�>.�=!����*��h�ɾB�T?�M"�zwE�V~��g$�v���o|��\�о�Ѿ�g��Ty���4������9� �9�K?+��?��?�?��j�3��>�i��4>v��>a|��s�'>}�T�ʑ_>��>9#��+�>�(>��>즴=�rȽ�ǒ�����UĽoɿ�ߓ�8��>��
�Cg�� k># ���>w��ĕ�>���kd��T���J���)�Eܽ ��MᖾC�۾F��?�GB?��>�Ź==�(�-�z˕��ּ�ū�4�=��y��i��%������_���U����'����W���ۛ>j�W��B���,}�>o(�Έ��#@>:�.?K�ž�j�������h=T�%>@J�<�[�#���ƥ���
�+UW?��9?���ܳ��h\㽔&>��?�K�>�%>�1��6���ߑ>��3?�A-?�.�鎿s��E���G�?�
�?��#?��j>�\@��qd�j��=7�?�B?���>�6׼�����>��|?��6?���>Z��`ot����ð�>�Z?�����>7 ?ɥ>�qX;.&.�X�R>�������ȼn&�<�\���)�K���c>���>��>���y<t����>�3ݾ����E;�^�+�F-�sTM��?`��SÐ<'�>�}=_�"�Fs�����Z�ɽ�M?���?a�@?��E?�z��"��l!��=˰.>N*j>v����u�1��=?��>t-��{m�ύ�@�/?Yt�?�?�_?էN�\�ʿ�P���믾贾�<>��=Z�o>D�����='��=�~��,=O�>$��>�K>�3X>��9><�O>!PC>�b���(��+��WĔ��Z>����A��i6����b��5[�Z���)ﱾ����Ͻ�]�������7�MY^�>bپiO2���?X��>Y��>���>X@=h�b<�3�b�J�\h��� � ž�!�Ⱦ��������U��ƣ�K{�<�x
���?��2�(T��$�>O��:sX>6�6>��5>���>�h>"��>n>��>�N>��e>QoK>6<��>�z�=ƶ���g����X��������>ꗯ����~�D��B �;���f��>��/?3K�>�Rﾄ����o+����>RZ���*��p��!{��E�>��>)���n>>�/�=�]���ҽ�!O>�Z?�G�=`�:�쾾�����>ee�> iھe��=q�\>��&?	x?'�.?pa�=K�>H+�>�آ>'t >��r>L�4>��t>��?�D4?K?1?���>��=�]���=��=�7��t���G��]ļG���d�<�&O�.�=�u}=��Ÿϲa=ƃ�=K'�<����l=P� ?��4?�D�>;_�>� ���B�E�O��.�kd�=�4m����>�>�?&?���>V�d>��	�E�ѾEFϾ�$�>�{A>��_�s�r����㠃>\u~>�:C?\�6?մ���k�po�<���=Y��>��?��?�N�>^>�2�Y) ��̿�ɾ,���E�ąS>+�P=.�)>��*=�N�=�V �q��+>n�<�׎=lW+>n�>�7T>���=vy�>v#�=M\�=Z�>MM�;��I=�ւ=)�<��:����i�tF�,:�
A�gzݽ�<h�o�}�
�it���?��?k���b�=�m��R	�o+��e�>(u�>���>L�>��=�?��]R��P>�r�[����>�Y?�
�>w>b�	�>�����<�ܲ>�8�>Hf8>U���`H��
�O�rΖ��x�>�Z?-g�>��a��Yf�J\��,���{>Ð4=�M9�瞤?x	7?�#���D������Cd��P�<mt���=��󇫾�/�&�>�0�����;��� p̻��?�N�?�꘾�%;�� �_{����~���ž#�"���ν�?�k�> ��V雾���ơ��n���	;>���>#�=��? ��>TY�>�o�?��?�V?�Z���?~��>h/?�I?���>�~>?P�=y9=������'>u!���W��2 ����=aw>ۛ�>!�=�O�>iq�>J��=5��=��0��q��v����w�<��u=;_>��2>9O=Lw>y�?Ud?Z뫾�Y+�����T��7��I,�;W�4>�[���=��@=��?�C@?I�?�Te>[  ��^����>�?�Dg?���>�����x>���� %��k?=�&�>L�>-��4_����HI�j��>���=�;&�e3f>��?w��>ܛ)?���6�J�����H'�G�<�y>�@�>��?V�+�7Už�J�B���b"o���0��ݾ���>��>�S��%F>�ƨ>�G"�F���s��=���B�p>ڪ�>��>B!�>���>W8�=D�G�\�޽B󚾗�L?(�b�Z���޽��ɾ`�������l�=�����\����$���d�����#��x ?:K�?���?��?n�(�|���|>��A�:k>��>���,��*��L�/>l�;>e<پ��P�"���&�>���>-�S�Ӿ�"�.(���ۮ�ko��j>' ��S���<�%��L��>�;&�{r<(�Ҿ����Th���w���yz��88���M�����ӷ����?��f?t��>�9�u�!�2�о�����L>���$���àp������|�W���)|�C�ھ�t����{g���>�;��c���`�����&��J-�=$�?�d������)�9�p��(q>��t>+�����o�C�������w?0�0?^�澋,¾h6��`��2?�	�>��>HS0�Zq˽k��>l�'?�94?Ջ����\o���l����?�
�?��a?�!���wW�Q�7�n;��r�?��'>���<�aU>N�."̾ �2>y^|?�|A?�׳=�`�}B�-�L?s=�?Y�����R>��]>�j=��+������ͼ�a�:������9�	��g������"W�=�8�>���>i���6��>��Ծ�	4�4,��U"��3n�[ӓ��
�>J����=�o>C�a=�-<�v܎�/������m W?t߶?��N?�4?c����E�r�<��@>Q^N>���>��$=u�b����=D�>���.Ik��k���t.?%
�?�>�?Ѯt?&~c��ҿ�����!��|NҾGZ�<�]��@?>&��oX>c+>��=��ռ���=ǸO>��4>$!>]F>�4d>�ϖ>*���4&��U��d��=>&��������G�,���6�������侂�˾����P���7K�E�z�/�J[;R�����>j�?1�>�ڽ>O�2>4�Y>"�1�[���д�.槾$��־����'׾#6��¦���]���Ͼ߾[�B�ؾrs?C1�<T>���>."a��ѽ=���>�m>|d�>��">�,�=/�D>�>�W�=t��=��d>���=m��>wz>����c���K��v������`+�>��b��j �{gu���"�!e��T?��X?���>w6��l����0�e?�>���=�����N���ʽ4��>fo�>_=�=H�h>�WŽ��<����4W>)?���=���!o���q�;1�>�s�>�����&�=�SG>�;?��?�Q=?U��=�j�>��H>���>�>>ɫd>�]>7�=>f'�>F�)?��#?*��>*"�=�r���)�=��=�rY�������d=?����V�%�ʽ��<�b=/ =u��=��	>�+�h�~��/8=��?�F?ܥ�=0�>���t ��SZ��u��by�=��Խ���>"��>}� ?>x�>W��>;�=�r׽�5Ⱦ��˾�$�>掇>�q��Q���/=^L?�c�>��?�Fi?�<
���0��z�>���>�<?�?6�d>�C>z��=I���ʿ���=Ka������5���=+nu>v�9��r<⓾����n*�=���=�z�=��!<���=l�>��>�0�>h��<5�>��=Z@=ݏ\>[��j>M���xZ�<����<�:�=/M�<�2=���ռl��� =��:��?��(?�8ͽ�Wx�H�;.�ڰ��^��>�p>��>���>�E>�����Z���;�nXZ��]�>`cS?E�>]�]:r=A��=Ӹ�=m�U>3Y>��>�A>酊���V��L�K�>�m;?�v�>N/��r3i��Ӆ�B���J>�=yf���?tF?gi0��^���!�Db����mH�>߱�;���U���&�ہL������.����;��?S{�?����o=v�㚓��������&�������?�s�>�XY�xq�����Z����=J��>��? ��=n�z>M>%?V�?%8z?j=?\�R?w��>O�M?_/�8?%=?v�?>�#�=�7��}T�>xj>6�>�,½5����~=`1�=Uf�������=�Җ=<�=5R�="^�?��7)z���<�`=�#}=f��=v��=.7>e_.?�_4?������sH����j�s��8����>���~�۾�uľ��>� w?��g?+�8?�`r=��&���A�=�>p�?�?$?S_����>j��wٝ��W�>��?�s=f/��G(��/߾�f��?��><e
��4�>�~?�?�U6?��o�j�Y�v���	���a��w�=�k�>�5�>AM=�`۾t4?���i��(h��Mr�4��a���8=�h�=��=?+�>A+h>2�>-f>G)">����؇O>C�U=���>0W�>.�>>CX=GT���)���.��O?�`Z�G$��e5��оL����b��$V�P����;�I���d��[���')��?���?me�?��Z?�Å��%�s.>�輙*�>��>�揾���J؏�?t�������ʾC?>��1>��5= :�>ѡ��;���v������'����1z��?~>����p�).=>��Ҵ>7������>�X������)Y�?�V���$���J�:ʯ�>q_������?�c?��g>��=�4���5pƾ=��+�r��i������g����Ͼ.̫��9���hվ���͚,��7%��b�>��K�޺���{�'+�鋛���>��#?�����þSO#�D}=& <>gH�=Bb־߅���ǚ�{��d<[?%�6?�6�����8}>֟?�/�>
�,>�ن������>�13?��,?����l����O��Cώ�[]�?�e�?aH8?�m���>��6�ȱ:5&?�
?P��>�ƶ�)���9�v�?W�<?���>-��X���&����>ҟA?��V�u�=r��>
߭>%��q�g��:�=�E��Ԛ;��>�/������N�	K2�,k>g!�>��C>}nX������P�>&�Ծ_$�3�1���M��)N������\�>�	(�t���@�>�Qνu9��M���{�h�A8F?v�?�+`?��:?�_����� k��{=��=Z�f>)�'<�<����/<͑�>'���S�z��Ӿ	=9?S��? @v X?�̅��e߿����Ɏ�B���<�F=��=``���<��>��<�}ں��=lb�>��\>�wU>G�+>:��>��>���c)�?������0�����U�1�T�ۼ"�*��ռ��ceh��оդ�����U�����N������ʼ�9Ͼo�0���?���>M�>S��>���=�k����E�ɽ`ؾ�]���|����;�������%ig�E���sc�i�����>��c=��>��>2ﱽ�
�=��>�[�<�4�>C�&>��=a"D>��>M�8>�m%=-�>y��=%�>�t�=ӈ��t�д+�r�Z�u����=!?&hY��!���.4�o���y��9��>��?C�>��t��q�VY�>�����
~��4��3żuU�>��>�Q�<�1�=���7�,���"�m>���>#>�����������z�=���>�㹾�`�=i�^>�@?�g?yS9?��=��>k�j>�ڃ>�>���>d�q>f�n>�?�&?�2?���>M��=�tB��b ="9=}*K�X1���U����޻Kq�=�F�9sR�<�ƻ.A/��y=]7=4���k�;�N�
?��G?L>\��>�/L��Z5��?��HP�IA>.��=T?
�>9��>?�>wj>���;#�=�K���.�>���>�_�~��a�=b��>�9�>�?ԞL?��h��]��I��>x�>� ?�� ?և>];->x�)=�����տ���61��Z���
��0�Vh����ɽ
#�=y�!�W��;��<N
`>�ۀ>:jb>8>�->�IH>�6�>i�>��>d_�=��=�2w=��Ľ7�>�����Lq=�j��D@�Nv��B�M���#���7�󜂽4v� �?${?I
��I��=bHP�x(�X�����>%H�>���>�e> �=\,���P��-:�X�q�|�?�_?�޲>�vx���=!E�=�̩=a��>��>\���n�=ti<��=z�*�M~�>�)U?��>w���*�|�pɐ�Ko6�)x�>�Y��9��fc�?s.?>E �%���4p%���"�~l9�c��=���<7d��BGݾ��N���3�(��1,�aH���Jg>Z	?W�?qfվ`��=DD7��7���a����%�_��r0�|��>Y��|�����4���ImǾ[l�=W�[>G/�>���=]�K>���>T?��?_�>��8?�{�>��B??�F>�!w>�&?zRG?n�>���~��|.(<3�>}h>B�b�,I����$��,�<g��E��:&^�<t}:=��"<J��<#qC=0��<9���ӽ=DL=k�<�+�=��=5?�<��?�+!?�̾��ɽ��a<�r⼧��Y���t�>`��=,��^ě�F �<`f4?X�x?D� ?_�>�0��7���:ѾA})=l�?&�#?�l�>�Y�=��>>1������ �=M݁>�ὼ>�������k�����>׎�>��n�/ٍ>�j?D�?5�E?�鑽m�L��=�'������cS>%�>JI�>o��=�Q��Y)>��h���&N���+�3|��J�u�=��3<��M�wE�=�<>�$�=b������Z�==�>Fj> ŋ>�e�>�k�>.�=!����*��h�ɾB�T?�M"�zwE�V~��g$�v���o|��\�о�Ѿ�g��Ty���4������9� �9�K?+��?��?�?��j�3��>�i��4>v��>a|��s�'>}�T�ʑ_>��>9#��+�>�(>��>즴=�rȽ�ǒ�����UĽoɿ�ߓ�8��>��
�Cg�� k># ���>w��ĕ�>���kd��T���J���)�Eܽ ��MᖾC�۾F��?�GB?��>�Ź==�(�-�z˕��ּ�ū�4�=��y��i��%������_���U����'����W���ۛ>j�W��B���,}�>o(�Έ��#@>:�.?K�ž�j�������h=T�%>@J�<�[�#���ƥ���
�+UW?��9?���ܳ��h\㽔&>��?�K�>�%>�1��6���ߑ>��3?�A-?�.�鎿s��E���G�?�
�?��#?��j>�\@��qd�j��=7�?�B?���>�6׼�����>��|?��6?���>Z��`ot����ð�>�Z?�����>7 ?ɥ>�qX;.&.�X�R>�������ȼn&�<�\���)�K���c>���>��>���y<t���>wȾ��M���#���`���nG�<��?U��2],=hD�>�m�=0D��i��s�ꢌ�N�6?B`�?�3P?�%?�|�Z�c壾�T>j�=I�?���>�Lսh�?��&?��"������N��99�>���?$y�?�St?��]�Gӿ�
��2���������=�%�=n�>>� ߽�ǭ=S�K=����B=���>8��>�o>�:x>��T>�<>�.>-���E�#�mʤ�ْ�\B�����vg��{	��y�f��_ȴ�P�T�������nѓ�׋G�����Q>�g��@T�=�v?;G�>���>\�^>&$>����oJ�?Wo����^~�6#��e������l���6��Qd�JL��"#y��[��?��=VO�=� �>���ԯ�=$�>��]=Y�>�',>�w>j�D>�d>�D>R�>qp@>f��=�T�>>�=/��3o��Ă.�{D�1�!�N�A?��c����n9�G"��S]��o�>�e?�B>3+��v��Vz��<�>"#�7�[��!���<yq�>=�>�{�=�蹼���є��@� ��թ=H��>�>:>]��<���۝(�Q�;��>��վ �=L�v>{�(?M5w?h!7?�U�=�M�>��`>��>�A�=/pQ>R>I*�>1g?]�8?4�0?ί�>R��=�{a��4=��0=@@��R�9���e���)�W�<*!2��y[=@-�=hH<f_Z=��>=^t̼�s;G��<�!�> 9?Uk�>4��>h5��=���L�vT��	>��+����>�5�>q�?��>���>�>�\����Ǿ�9߾���>��K>^�i�x�*�뼜}~>�vj>�L??/?Sm�<n�Ƞ	=W��=I'�>��?��(?���>]!>\�ͽ{O
�W�ȿ3��D��V-�~K��&���j��C�	��{���%�
ї����=���>ߌ�>��$>J�>�r>#h�>�F ?V�=ү�=��\>-y��=��:��>�3�K\q=�dB�(��	4�6^ͽ��o=���;0"�8�l=!�g�?�3?5��>��]��/��Xw�C����	��~>�Ү=�L?>�=�>���=��'�!�F��W-��7���>nwY?�a ?��S��/�>�+���=X�>�f�>�F������q����'�m�=x"?o�'?ϟ�>�⽍��-���d1����>���<`k����?��?�9�f|����y��l꾂� ��5��.0����?�+����(��V���W���d��Ĝ;?-M�?��n���ľe�����o�&����Gg=�_�D/�>x߈> �e�od���2�B.ƾ[L��fqI>l=?�茾��?��?ds�>�C�?q�)?#�;?i�3�oP�> � ��h�>��>�z?�{�>�v?fپ=VǨ<
u�Լ�=[혾0��8e��屽����䓼�D�>3=���� *�	�P����<k.k=����α�=����@Z
=�<�=��a>_�>E�Z?i��lᠾ
ޔ>	������&Ń>2�<��U��žeڴ>�ʓ>s#?��D?�>�����֦G���H��b�=U5?!B?�l?O#>�S�=J���X���I1�=�V�><�)��Ţ���ɾI6��X8=Eڸ>
d�>�>�a�>`u{?`�6?�t?�W��,��gs����@�������7�>Tk�>�5�=:RȾ� 4��{��a��S1�����'M���a=�=�=���=.�1>ׄ�=}]>��<=����ڽS�˻��4<}�>�>��?��Q>=�1=~���z>�h�P?��r�A�n6�v��D�����>�G�>"��>�p?�⼽	2��ǘ���
�DQ����?��?�o?y�)���꽋�=�~�=mH=2�X=�ä��,�Z�A�v��=of�����y�,��4�=f�>s�>��A�a��!Yr���X=�c��;�x��i�>axH>n����)>�;d���Q�p�ξ��8�M�2j���=�����>qi�����{܀�l|���d�?~?���>�x>N�>�:���H���A��=�v��t����1������'��In�u6��(e�|/�Ԫ����>��Y�/?��a�|�
�(������p?>Z0/?G`ƾmѴ������g=/_%>M)�<k<�֮��������?eW?��9?J�2��9Ὧ�>��?�w�>��%>%��T"��-�>�74?A�-?�W�]��`6���G���j�?a��?�pI?�i�etD�F��[Kнgs�>� �>-��>1��xzʾ����ϩ4?J)B?"��>̔⾏˔�+N.��Qu>��M?����0s�>���>ϡ�=��\�\�������A�H����=5A�EX���L���;���>(��>ޘ,>�3��l�����>H�ԾJaI������o����Qɻ"�>�o���<�B>��<�_���n��������VJ?j8�?F
n?��(?��G�5�=�˾�}K>ښ>��P�>�?~v)��#�>��?or�)ށ��7<�h�?�?�E @���?,�e�iѿ�T��E4����V�R�>0,�=�8>?�n���^Ux����=1f�<H�A>I��>�9">�$>�I>�>�桻�f�^�%�����$Ⓙ%�F�v^'�������!�56	��}A���龜ץ��ʨ�͂��߈�N"��`/�p�-���e��D�=�D?m��>V��>�n>���=����n�_���y�������d޾��ܾt^ƾ#�u�%�Q�����u���������]/?8�<��=pD�>��'�b��=x�>X9=>�:C>M>��R> $>buH>�+&>HL+>�B�=3y�>X��=̅��Ձ�7V5�3mJ��(�E�@?b�_�f��'c8�Q�־^Z����>��?8	C>5)��5���x����>������W�&�н^rӼ��>9��>.z�=7�������q����Y��=��>�%>C߻;����
P���T=HS�>��;�b�<`=c>K�?/�a?��+?�
�=�"�>s�)>���>uO�=+��=~�J>�&f>R�?�<?J�:?�
�>DŤ=k�T�w~�<II�=1jH�G9W��G̽�CҺ2�����׼j�<�J�=�K���\�A�R�7=��Y����[=`@�><�8?�x�>0@�>�f9��>�NJM�m8��>�#�C�>�l�>��? �>W��>�4>�{c��þ�#�� �>��A>*V_���w��U�sxx>�rr>�]O?t�1?O�h��Pd�^�<s9�=�#�>��?�K)?(�>�i>vK��s��ud¿,������b�N�(>�昽#F��@�����`�&r<�ш��W>�ħ>@��>�R�=��:���=k?>�[�>�wU>l�=L�9>���ֆ�=�-�U��2V>�i�=a���s�;�0����g���a������_o�<%FB=��5?�x�>!����xh7����TC���L�>7��>
=�>h�>?F�t>�C8�K��ck��"�p�>�vR?� ?�{н���>��νo?��4��>ٞ�>����?����������s��uW:?�E?X��>�N������l:��`��w�>��7=�ry��?{Δ?x�N��N<o�7�j�y�o������2y�h��w��"D�_�@��U ��&�R��mj���z*?�s�?��ʾj�/��K������80�a{��5C��n�=�1�>���=�7����Fi=�i̾�UP��Ha>��?}�&�w�A?�n?��>覅?=�4?���>V;�<j3�>�0�wF�>0��>�D�>��?��9?�����~^=�@�=�[���3���ƾ�
K=�<�.��4�:>�+�>�
< S����<��Z=N�]��O�<�>����=��~�s:.=���=o�3>�;?$�L?�JK�5Hj�I�*>��IJ���=36�=��ؽ�9���u> 7>(B?]: ?
��>P���U���+�$�w�Z� >�4?��A?�L ?5�ﻪ�=ν��������>�~�>�wͽoz���8ʾ�%��:9=s �>�(�>K�=�Fr>�}?��:?Qe?�`��+���x�J!+�i�$�fμ�S�>��>��=�Ҿ�9��w��b� �2�c��*xJ��\=O��=�h>فK>d��=�b	>���<�h��(�ݽ�?���[ݼ���>�w�>�t?a�X> j=����χ��Q?ˊ
��<��N�}4���%z7?�^7?�"�>ˉ?Ŵ���ɫ��Z�������>��?��?|�U?Ծ>��\��
>�M>�8�=��=�\^;S'�<��`<f�u>c>�^J�֖0�p4f>���>�܀>o��$��n�վd�����L�&�=���d�Ҿ��+���꾦Ԝ��,�>p½�y�� ���L����r������vվ����>����?/�{?���>��>Y z�iȾKq���*��䗾�~�V�Ӿ�{W��@j�����k�������.�f�=�E�!��˛>�yY��@����|�n�(�����^?>C./?�Mƾմ�m��9h=@\%>n�<GN� ���A����!�/iW?��9?�5�{.���:��>�?-^�>0�%>�+���^��>154?H�-?K}����d;��5����d�?6��?>-H?����V.^�$ �	ټ��>Li>�R�>�IH�e�k���+&?�C?���>������tw6��S9>~@<?᧌�M��>e�>q
>.�=��FX��9�b��)T�;>5X��*[��V��� (�Eq�>�k�>
q6>_3������f?�{��&sV�!��2��E��'4����>@���-�=If0>6A.��i��c�����Bj�;_V?".�?	PS?Ϸ"?�h�����m��.>ۼK=��>{�>�����>��%?�:����z������>;�?e��?�?��b���̿�'���u�e[����?=E�F���>>U���BJ=x�>s%8>��r>���>#�>�S#>'A>XQ?>`�2=�����$#�
9����˰D��Z���8�A�����)\��mž�xN�?�����Խ(�齉砽Ą�v==�E����Z	>�%? ��>d�Z>SU@>�+y>@���Q���m��ʪ�OJ�"����]Ҿ���w���q���������U=C���?S1b���\����>r=��? �;r��=��>��=���>�>�%>��b>�ف>�
�=Y�>��=R�X>��=�l�~	z�ơ/�$�$���<��1?�\�]���@�/�z{Ҿ�.w��j�>�7?m>߇$���&ry�1�>R��JB�T��oJ����>l�>>�>^P(�Çh���p��"A��B}=[��>y$>Z%w<�Z���"�[�=��>U��Ȃ0>	,>��%?�k?�<9?�,�=�{�>b�>I�>e�>�[>�),>��>�p?@Y*?�i'?��?���=���B)�=���ϊB�S�<���i�v^4�U�=N���>h)�=��<M��=X��=�h�{,�;�"=y`�>i�8?rJ�>2��>�~9�<g>��3M�*����>?���x�>b=�>��?�\�>���>� 4>��c�͝þ6侙��>�A>�3_�v�w��]�Y�x>�mr>knO?��1?R�f��@d��%�<��=>�?�u)?�1�>λ>2����N�j`���n�#v�^��;�� ��Z���e �F}���>�N�=��Z>�ف><�>���> �\>��`=z��gZ���>�>�4=�)>h��<��S<�]�=ޕ<�9���<8d���c}�X�<���<�L�;�y�=m�;��i����G?�f�>b����O��ϥE���9�����H4?U�?�!>_P ?�>>�.7�BeQ��V�{�����;?�W?�0?!&���>f�2��ժ��/�>.�>�p�����8�q=�`��1̎�TO?��)?�ݰ>5�	oo��y}�/r.�H߮>�W[=�"��m��?,r�?��f���}<�0���b�	;2��z��d����H��cn�Z���*0��6ľQi+��z߾>��9�3?>�?�$��z������,:���Ji�*ڃ�4�T=I�+=iH>��>��Ѿ ��xw!�D������ԃ�>���>q���ZG?��?�|>��?�k9?��,?�fI>�?.�����m>�#�>���>{��>7o/?�����c>�8���Z�'>x8f����F=zn�A '�H/��m��>�p�<�=������>':��O�e�~�˽���"h���=}-!>�C=>�?Z]?i�S�y7g�D�O>k�)>B����f'>S-'>A����	�� �=s7�>9�6?��R?j�>kq���N��{4��m&�l�>y3-?w�N?B-5?��t��8�;�5辫������=���>����GȾ ��#�S��;�<h>��>r�X>��f>G�~?�OB?��!?yF����.�6w��K+�,���jdL��2�>��>���="k۾U�6��Fs���`��k1���9��F���<���=ޚ>F,@>��=>�>E�=�Y�׽��/<�C���v�>���>VE?��\>(U�=�_������W? h��� �m҇�R��W䯾��9>�}�>�jV�HM?�C>ȅ�׊���L��=�O�?���?a_�?(ې�=���"�=�\{>h�<>j9�=1�m��CB<%�<>r5�>EЉ=c�t<�<��p(>9>tAC>��'�7K���`��簼�	����_��<H��i��а�4����Žq�%��澾K@�n��ڪ���J�j`���q�T�+�����*������?.�o?�>��o>p7_�� ���*辅�2>����&�¾�Ⱦ����g���$Ҿ����d ��$��f�⾲;�>�X�J��9�|��P(�Y����E=>x�.?vľ)i��]���s=c�&>��<���<������{�G�W?uO9?��-�������>�?���>�" >ҟ�����e�>�3?a_/?gٳ�ō��ދ��B��m��?")�?	�R?~νSY�;�&���ĽW�?H(�>��>�C�8D�����ھ}t?�W?.?��LĔ��c2���@>�@?�Sa�7 �>Aղ>�F�=��K@�<�O�!�d�!_<S>1퓾d�v�5�<f�?>�1�>�>�>�EW>��]�V�$���?/̨��A���)��3!�7�߾���=�(?����<��9��>�'D>4�5�s���(���v��|H?:Ŧ?J]?��?d�+w���!&���9�2Ч�)��>���>X��7#?9�;?A,��Uf��ju���>�1�?��?��q?ii����˿�M2��I܁�T�j>T>�D>�z��!}�;B*�>K'6<�*��p|9>DҞ>٬>|�>�=�=��K=�G*>]3���q"��L��Ȇ����&���O�%�$Ǿ�<�'{���ܾ�Rh����徽٩�<&G=췛�����N������&=� 3?�*?<��<'�>����ͷ�"I������U��k�kd־վ����<�M������r����ۤ=L�9?B�N>�`�}�	?v�@���=/��>���``D>;�R>��:���>�<W>�(>�#�=^q}>aѻnV�>��->����R������x�M��+��N�I?�p������jP���l��b���5?K5?��y>6}B�����r����؇>U�=�猾�f{���
=Pg�>�Ƥ>�I �
2�;A,��ܾ�Zd��2S>��>�s>wVd>i���i������>�1���Fh>ZK>��$?��?�X?��<͏>��>�=�>g�>���>�X�>�M�>k�?©F?�=?s��>vS!>g p��O�=w�}=H龽B�=&���5<0F��MB<1�����=��=�ͤ=~�=z�={#��X����<�V?��1?F2�>}b�>�,���A��A�<6:��j=&׶����>�E?� �>�?�>���>�h�<�諒��ؾ�뮾k��>�b#>�Os��|���3���>��>m�@?��
?�4���҂�"r>���>{�?��'?h�:?F�)>@�=�������Eǿ�\�����m|H>��5>?s7�B�k����>>+����/۽ѻ���j�=E��>��>�wl>��t0>wS�>:�M>�>'p�=�����F�IKX��$+>��2<��T�(*e�q�H�5��=4��d
���"��l�=��>��<��:?co�>���<�O*����m6S��?���1?��>fi?ˠ?H�=�	�6�R�`��K����?��z?DL?��}�>Ռ`��̏�ϥ+?d��>��(��AV��\X=�BϾ�+̾�?��>w�r>pɡ>��h�=�A��31���?Fn�=ږ��{�?�[�??!U��H��B��S�����
{)������̾����S-�<'�����@�[�돾�����(?d�?1'���-���Ǿͤ���:����i��E<h��>Z��>6Mɼ<����f��R���T5�L�>��>1B���?Z[?�"�>(�k??n?7PE?N�1��r�>��A<��>G��>Ϳ5?�f�>��?zhe=j�>���=A�L�����%���hn=A��=dy�=�J	>��">.�����UoX>���=��{�^gȽ$�Ľ~C�����-��=�{�=�x>5&?φh?�g"�&���_>�[�����7nY>)�;=!�n��R�W>�|�=�C?��L?$�?໧<����8�|�"��,�=ʥ?ץa?�>��=��d>�N޾JOս��=֑�>�u1=�9.�W��(��?1��s�>xY�>$�s>��q> j}?4RA?� ?�'�t\0���x��'&�Vx����\��1�>T.�>�{[=�����4���t�"�\��+/�[�ü�W@�
��<_��=�>��4>�=�=�+>��3=/���Y������<�g�;��>���>
?y�W>��h=s����2�M?B����d�қ�QLݾ����3>�>����ľ?��)�b�|�=Σ�y�/�27�>C��?��?��r?��G��4�f�j>��q>=�K>���=̱+��3ӽNv��̠/>�*F>nz��n��Q�Ļ� x>�p�>E���0ʾ��ľ#�˽>�����J�2��!7���x���B��?c����Q�$���@ݽ�˾���������^�����&_��皾k ���mt��ē?J�?
#�>\7�=ES�V��q{ؾ��=Cr?��p��p��ZP��"���������� ���N���1�A����>j�I�o���t��B-���v�8>�6-?
�ʾ�z��c����=�&>�Z������凊�J��|����V?��9?H.ݾ6��Q���+$>��>э�>}&k>���i�'��>�y9?:i ?m@D�i���Y����
=�޽?㙼?�L?<v8��=�i1�|/��a�>�R?~��><�s���&н��?�$%?Ә�>������b �]��>\?$�6�/wJ>E��>�I>�Ni�`t�,n�G��D�/�ur
>c2��7uh���ƾ�i��0�=�̿>�"�>��_��҈�yV�>پ��J��辍7,��0þl�$=���>~g���>Vݜ>�¼v�@��`���ʈ��T�<��A?=�?��V?�'?��aJ���Y�U�>Ҥ�<�K?�N
?�����m!?��<?M�!�Rx������?�7�?�� @Bk�?HS��̿\?�������j����=?�=�F>l��O�'>i=�=�U'��O/�=>�$�>�Rj>�<�>��U>�4>`�$>%d����&��Y��8$���I���#�?���L��޾l�f��;���ǾgL��~7��\�n7���4.�]����ŉ����>�E?
9�>ڍ�>A>��#>�慾��_q����p���a���zXʾ�{�a�+��_b�8e��V0��a� �D?��S<1�=˭�>H��W�>7b�> �}=P�!>�MC>S�>|EJ>��3>
�J>�%>Q�R>�z�=���>�@�=X��0p����1��7������=?�hL��P���m?��Tɾ��_��>0�?W�8>�/.�0���#{��!�>���;d_R�)p��9;	g�>t��>�'�=��w�ļ��@�d����:�=N�>GoJ>�=��y��u��<�k�>�Ӿ�V�="r>)6)?L�v?�F6?�y�='�>`c>T��>Ȱ�=��K>s�O>�Ћ>��?��8?hZ0?/��>|�=6+f�ͺ=��&=�8@��V�?��������9-�r�<[Q3�IR=�'r=�3�;F�c=ůF=���<�;�- =E��>��8?�<�>��>Nl7��><�Y�M���e&>$k �!e�>�a�>��?�#�><��>�(>������ƾY
���>�EM>,^�Q�y���*A~>ҡg>H|M?0�-? V���i�R�<�L�=�Ų>��?��*?YM�>�><�Ƚ1��V����8���D��ߍ=�`�=�5X>�f����b>��� }ƾJ�=U�>Zq>�qp=,F�=z>5�:>�_�=���>�:>i��=7��=��H��[3>����a�W`=�>I=E��.����uP=�a̽�6`��i����&�����^ܷ��pA?��>���o
~>e�:���6�t�����>:O;>���>�Y�>$��=X����7�4�#�D&˾8��>�'9?7KB?�"����>g�b���ۼf�8>g��>,�>���<�X>pï�t�n���D?�j?im�>򤢾�`�n��B?�p��>>��=ʿ���	�?�p�?a
\��戽�E��r�q�D�ۈr���i��J��o%����Y0�3/���,�Bsܾ�옾X�:?���?@����g�=�x��Aa����M������u
>d���>NS�=�Ǿ���q(��?ǾGe��&=Z�?D0C�*�+?M��>n��=�o?ŝ$?��1?d,�5�>tPX>��?m�>6��>��>��P?��=��8=0�����=��E�!ھ����B���L��+�=T>^n��ޚ(= =ٍ=2|Y���Z=�4���ī<{ϓ��*�<u*>��=9�?�^?���|}��h�4>`�:KH��#��>7(�=sMe<pR侞~I>��U>ן>?�N<?b[�>���[�����&+��a'>	1'?��L?��?a2D��\H>;��?ơ�_��=���></(�qE��0E���$�(��=z�>�ڹ>%�s>
Bh>��~?�A?�!?���%�.�$.w�@/+���cV����>a��>���=�^ھ��6�Ƒs�a��1�f"7���G�A�=f�=Ц>b,B>�ڽ=~!>��=}���Uؽ��<�ě�X�>�f�>��?xq]>���=Ԫ�[����b?�_�R&�U�!�ud�~���ƥ=��>_���-?ޙ�>[���E^���g�H���k;�?c/�?��?.�\����>G�>,`�=��^>��襓�	�y���K=��������߽��<D�>N`>�Ҏ�_A�����~�J����[���=3�t���վ
��R���z��������A���H�=��<��7作I�����}!���}Ծ!�?o�r?� ?P�>��z��N��"g��P�=����f�f�-����ˤ�?f�������7��?��E/�F�>,YY�n5����|���(�?=����?>x@/?��ž�ߴ�K��G�j=ʷ%>d�<8�ﾟ���Q����m��W?Y�9?-�뾸!������>�?4�>-%>����`���`�>6H4?��-?c���^7��B����;�?���?q�L?C-���QD�O|�	��J<�>mw�>6��>�=��־[���9�%?�,P?�� ?ǥ �6����H��F]>�Z?g����D�>�Ϛ>��Z�K��=���<���Gu�����V>c񌾷�L��C\�M�=ϥ�>�-�>2>>8����y�>�̾��ؾ�8G�I���A�����r��>�m���j>7@��&=��'�i���P����8�/*?o��?�iE?s(e?
�R���|w�-_ >[�L>�	�>D�7>�)����+>��>T"]�	1��н��9?��?V��?��V?q���Ϳ=斿1ﺾ�{��b�> �=�[><����2�=7�=��<�6,�:�=�Q�>6�z>qr>�5a>wz6>��#> ����&�\ب� ���2�֑�\�%��������MV����������qh���&4�Zߛ���_�#hC�����J=��Qg>�{?���>8m�>�8>���=<x��J����l�7����9H�O����M颾�{� ]l�KkF����~�
��?���	>���>��x�?)=>ǂ�>���=&�>S�X>�>��a>��5>��s>�/>,2>�K�=���>S��݊��X���������=�<?<�ľ� ��V��	�{�P�� ;�>x��>5Ȇ>I�¾�Y���y�r��>�ޗ�Zߥ��@����=\��>�;�>�F>�;O>E��QI�q�B���κ_��>ma>�y��T��[�_=�?�=���>��վ�]=�2>�?,?��~?��,?(ܭ=$n�>ul>:�>_P'=�}9>X�x>	f�>��?~54?�d(?��?�=�wZ��Ѓ<9M�<��I�p�������c�Y������������=�h?�p��Ň=~f�=���vz׼O	�;d�5?���0<K>%��=�a��E����7T��5V��8�����S�]?ݵk?�Ep?�)?ߚ=Fޖ>�E�>�۾��k�a��>�mg=tJ{�(V����=N�S>f0�>��?��>I���u>X�{>�R�>�fq>aA0>S��>O^�>�
��m1�����,�ӯ:�<��>�|�":����<觯����>5;,?�%>��];�0�П+=���>*{`=s�����>|Y�<3k�>�� >�+=<��=����>*F����:J�>:��!ڂ��3&���	��	ǻ2�#��՗�O��/> f��w0
?�6=?@�O=_�=>�G�%r������)�>�}v=��> A>H�+�
�!��Hs��RZ��k*�T��>Ё?X?�ی�m>� >��>!�x=Pԫ>�<�Y����$�=�TF�Λ�<�n�>��%?��l>Ew�P��U����g��>�=�61�b��?�.?@�-�w��=:J�Te�"�� =;�q�>�q�~��f���&��$,���<���ս�3>]#"?�T�?�D�S�=ǝϾ�R��Y{���h����Y<���>��>i���0���.�¯����,U���>��O���?`�S?	�G?�N�?Ӣ�>�b?fs�=�>�>�E >y�>��>,�>7�p>{�R>�5>�9�[���7&=,o;���˾ �E
��g��>�>�%�>��>8�0<���=ᐩ=�����ɽ�a<x�l=���=��>�f9>�?>1�?(��>�4T��k��U���ay��O�9�>�=a���N�:|�(>�*�>�Y?2�?}�	?,��>��ߵ��龽�>�?��.?�>}x=_wq>3�¾p�A��+ �)D?>L��<X�F�8�ھu��޼�[M�>A��>��=F��=Y:�?�[_?�fK? ��X���3'�>�G�Q�=h=� ���T<��
�Ku6���T�����`ڀ�b�X��Op>������>���I>�}���w(=�����Ǥ=�>�,�=
��=O��>y�>;`�>�Ǎ>P^=�6羔� �w?S?��P�0�!*��j�D�>,��=�_�>T���ʑ>�˟���h������?1M�?Eӽ?��K?O�+=>�ڹ�>��>�x?��>����>��$�D�v�q�ȽM�2�7�2���؝t��.����H��I������#�����,/?���+��N��9Nž�����޷;����2� �@����,�U���	K�b�y=�]� ����qI�h�����?l�?P�?}���EY8��5��,�e� ��i��þxþ��l���������b�,���8������|���>>da�<������2%�/��9�F>��2?ʏɾ�;����e��=O<>�-=Y�,~��}����ШP?"�7?y �ݥ��|Xý��,>\�?I^�>=>�.��Ǎν �>��)?��(?��ʲ���q��"'���?���?z]?T퀾00j�4zL�ႏ>GXf?1�?�{q?�Ͻ:�����ž��=CS?n�_?x����K��񾡍%?��S?1�R���>k��>��>�-�=�
�&n��䡳��Ԁ>9n	?�����)-���&�nW���>?/�>�d̼�m���i>�
�>�r�q�N��H����3�����<c�?��B>]jj>H>`�(�K댿P���X����L?S�?�S?�O8?�Y��Y[�����=|�>|��>���=�F���>RD�>���q�D�L�?�3�?���?M�Y?J�m���Կ�����ǩ����y��=�_5=F/>���>>��=T�l�f,��o]>錒>J�>�>^V>$�3>��>�[���-#������&��{��������-����������ɡ�,��&��������=۽N>+��f���tҼC�!���>t2?Gs�>�>,>�G�>U	<�EM��!���U����о�K�����/��	��]���$i:x�S=�ǾŎ*>#��z/?;��S��3X�>������>M��>=$�>?e�=��->Y�,>m�I>��'>O�>��>4?�>Q�D>���>D���)���~}���f޽��J�A?�ed��&�r���!�}���ߌ5>���>)��>���=����\����>Ƽ <n���%81�*��=���>o��>��>�Q�<�N<��Ǿ�_�ƍ>�0�>͚�<r���3T�'7<��!�n�>c9��J+>�ǖ>}7?�~?��D?��<W2�>��>Cb�>�y�=9>�X+>0��>^�?bA?�A?C��>c�=�S��|�<:ح<�,J���i���`�x=$P��+��H���� k=�w�=�:D���ϼ��`=Q����X =kg�=�?�^^>�,A>'������}:��X`��#����>y�>(�4?�4A?g��>�Њ>��>/t�><W;��.������l>_/c<��y�C�T�|�> ��>�F�>�J$?��>+_z�_�;�/�>�ڥ>&
>�Mk>Ct?鞿>o�/�^T��m� y���7�%Q��5��=�֑��#�=b<�>�&�>�f��j���=�6�=���$>��<�"(��8����=i��>毢=�>{�ڤ8>�
H�����)<,���5e<�Z=�B�@�G��=��ּp�ݽ]t�=䛽=�ؽlm�-���#�?�B�>:h+>����޾�W �pV���$�>n4�>af,?^�?w`=�0��%*��f/�ǞǾ�>�"U?aI?;�<��/�=
>��=��u>��M>1y�=�&�=r7�=�� ;��@:;s>c��>��>�ƽ0�Y��~�3���eV�>���=jʏ�tޠ?ʋ2?�#�����'���=����:�<Y�l�􋙾Q(��TR�y|C��i������0�c��<ą�>�Si?�]���_齼yپe0���k���·�9*>J>]S�>9��>�]=�)�D���J�˾g����&��$r>��/=k�>Qw?J�?\�_?��?��?����	?��=:��>u�>k�?�?V��>��{>��o>��<$�+�v	�i��qo<�Ȋ���=0>!>S�'>t�<��=�@=�(�<��6����iq<�eJ<��=*��=�v�=�>(�?�;?��e=�2A>, *>\�4>M�=(
��/��L�������8YӾ�����52?
w?j�'?>�>.�+�"ة���r$�>�f%?{~T?c4?�͋>��>|�es��C<į�>h�v��\쾵���_A��I==� �>;\>K(�l�>9Fp?>T?�T?N�b��K'�qj�/���\�=3%�=�i�>��>2� ��m��q3�®|�؈q�<�'�1�>Yc��:+<���=�.�=��>�3=�uR=��=�����콌�= ,=��>q�>J��>�Z>�q<�׾�#Ⱦm�:?hK��Z��p���k��g^_>��>� 2=c;��Tg>��)��Hr����K�l�>?��?�)�?H�?�H����
M>4�>[��:�����6]��Hܽ_h>��>�>��ƾ����f>�=��3=������,x���jϾ�Ͽ=Qܪ�<J!��i���O��q��*�¾����"����G��F�tվȄ+�/�p�r5k�=����½'����T����߾? �?7X�?�8:>L�S�?�"�.έ����0F��H	�v|��<m��U����I��??����� !��˾+����S�>��`�Đ�Yw~���+�����*>i�,?�@��-��s��L�=�\$>�ܪ<����C��B��d���V?�]7?��꾯l��,�ֽbB>U/	?���>��/>�팾���?��>��.?A�&?���}Ќ�������?.w�?S�M?BRͽ�p\�BhO�щ=\[?��)?�?F�ǽ����񫓾�C�>By�?L�O?]��_���=�o��&�>��>�i��(9>K�>;��>�CT��ݾ�<bծ��T��!�);���A��)�ȾS/>�A�>�y>�Y_�Qڬ=<��=�*�>�C�W2M�1�H�M2�ݫ���c<a�?1��>�e>�2>=�(��ތ��n��bt�C<L?S�?��R?�w9?
|���C�2���	��=SL�>�>�Ъ=���R8�>���>�6���p�6���?t*�?���?k[?��l�9GӿF��y���/��P��=K$�=��>> �޽uǭ=k�K=^��\Q=���>Տ�>�o>�;x>D�T>S�<>��.>�����#�ʤ��ؒ�"[B�� ����xg�I|	��y�����ȴ�-�E�������Г�P�G�E���X>�읾hl4>o�#?�{>�<�=��@>�����]/�����9Ϫ�^��;9 �$��� �������҂�Nt���G!��N>x�&�6�?����D�>ff�> ���AI>0.>[0=�+">��>Zm>=An>{��>�ϛ>�	�>�>/7��u��>oe=��"v���4�q�L�a��;��D?s�e��l��)F/�<"ξ�z��]p�>�?:~M>��"�񵏿�{�1�>�,�kt��򽊫&�y��>��>��=�՘<p�x�c��"�콫ҥ=>�>i�>;�A��|�����=7X�>n&ӾfJ�=��i>�)?ww?.o2?pV�=/��>	�`>��>RZ�=��E>�9Q>�
�>��?�7?��0?�	�>ir�=�bW�O�=˴R=��;�x�t�v��5\ż�P<���<A=����f=;/\=��"��c<=�Ld=K�>�7V�:B��<Ɯ?	 �=W��>��o>��j��5��P��*ڼ�ܾP*��,?��]?*�`?K)?�	w>P��=���>]��\�\�sk>�=$�����$��Z�<�+=? H>�;?)3�>M2��´G�>�ϔ>f��>㇑>�L�>�=m>���=�}������^ӿ�9�~ ����Pe>+�m=f��<��>�9<��k�f=�{�>LD|>���>璧=h��=fz">���>��)>b3�=��=��W��k��-�o�A�+�v�U�����y:�q�]�ׂ��0	�-%��μΐo<�~+��b����?9?ho�<�u��ܽ��4�U��{�>9��>���>�)[>%Sm��j�A�w�9J:�n�.?BAJ??�Ͼ���=�
>I�=;B>�&>�Gv��C>=��@�$�����>��?��}>��)�
�i���l��b�y��>ZC]�ϟ���Ǔ?�O?'p'�\�����"���w�H��m�=.��x�)*��+�	�Ϫ2�c�#���k���=�q?���?�؇����������=�������ʾ�z)>�=���>�^A>#�;��#���ݳ�������Z�����>��<<��>��?��#?*�T?L�?v ?�ݹ��l�>RO�=�b�>s��>b�?1?s4�>�x>c�k>�:/=��u��^	��S{�D��;��+�m��=��>��">x6E;Ì���=�w�<�{;���%��<P<,�$<�O=���=��=�}�=�J??h�Ҿ+Ӳ���>^z�>����h��B��>�u���\���DV��� �Y�>)�i?:�>?ݔJ>��x�MV��-��z�>�f�>��"?_l�>{�-�,�H>ҕ��^�¾;E��ۍ>"�=�[;D�1��Ᾰi�<S|�>q0e>߶����=��?t[?&?���c�"�h0徛'��F>�8�>l(�>�� <	�ν>,���X�����x��S�`�EZ�>��w���*��f�l����8>�T9>�.>�<>�9��CQ�6�=%->���>�k�>Y��>ƍ5>h���X����ؾ�C?wI�e}1�,l��$���qM>��>�<����Ȃ>�q<��2e��e���A�w�?ZX�?y��?�N?��s����2��>ݭ�>�=�>q*�����L+�=8^G=b<Y��;��@���� V��m.���ڨ�5r�� �m?��a�a��;Ϳߎr��]潯�T=i�[�!�ؾ'�*=۠�=��-�S���%d�N��Kh�}�������N��"���@���`�u�=0�?�xa?��>9y/>)�f�ј����6\	���¾5�潄i������/���:����־4#�p����Ⱦ�O���j�>\<]�2�����}�X%&���u���N>�3?��þ�*ľj���5�=n�>>e�"=���������ֽ��M?2`3?h�1�����}�>��?��><(>o?t��T���x>�+?yr'?��y���������e��w�?�p�?y�G?�Nb��7d�� C�YNX=�?R>�>T�$?��h<��?�仡���>�^?5�8?;��ŕW�@����6?�?̭��Ё>�s>\Ϛ<JX>�@
>�)ƽ*x��s=�>lo�>�r�>����ܼ�����>�>�>^0O=�g��v�=�?�>��u�N���H����X��}�<Uv?G���>��i>U0>�y(���ӓ���� �K[L?�?�?;hS?+�8?T���+��>墳ӳ�=뗧>3a�>}��=������>��>���-�q����?�?P��?!NZ?n`m���ӿP��i���௾���=<)=�|R>�J�x��=b�=ur�;��Ҽk]�=���>�tW>^�[>�E,>�P!>e�3>�o��[��M��9����KS��8,��y'������H�9�_�����XѾ��Ž(ƽ3黽!�S�&=��c��o���̶>E ,?]�>�-�>\��=�"�>Z��?���?�/�	#��?����Q˾&���T���璾$���,��]�徘�'<��=p�>Ö��50>��>9D}=��>������>�!A�@!�=��V>G=>z�="�(>��<>�p~>~[=�g�>���e!v��E��12"�����1�2�>q��$}�=�@�au�=��)������T�>���>������I*�\��>m� >�!��*�佞��>E�?)��>6/�>z�.��:�k3���\���!����=Pr=�1��.v���sG&>�s�>̾w{�<��6>�_1?�w?�;1?��>3�>Yt[>M�O>	� =�w/>=w>��>�?[�2?�64?ܧ�>�=�O&���J=���=�!P����R���<a-��1��띵��'�uD�<�4�;$�⼍?�=�f�=��j�>��;���<�>
?Bu>�\>-:>XZľ8�g���^�wԠ�ah�"�3>p�,?�w&?)F*?���>�[�>`ߟ>۪���\l �,��><�= �j�}n�E�N=:�>�e�>�=:?�"�>o��=���=/�>!Ϭ��%�|Ҽ>\.?HV>�����<����lӿ�$��!���e�*`�;��<���M�i��7g�-��������<��\>��>X�p>�E>��>�<3>�Q�>�HG>UЄ=��=�0�;)�;	�E�:�M=� ��AG<��P�3���/Ƽ��������I���>�-:�F0ټ�>؊5?_3�=��>䲠��g�*%�����=˫?W��<�SB>&���3�xGk��C�2���PO?�E}?[�?�RR�ds>O�$>l�_�O�s=�X&>!���]=�d�=��f��f>�-�>�>��>P�`��������I2���?�N�=|g��`��?�I?ܔ�ˠ��C;D���A������=*��������>�l�ھW��,Lھ\Hݾ4�1��K�@�?�5w?���m�<�Ǿ����b�l�����q���=(W"?��>��=�H�e����:'���콍��=�s.����>�-?��#?��N?�;�>��	?����?i��=���>!g�>���>(�? 3�>[�>��X=�W��zW��L��ĕ�}	R�V�=Z>9 5>@,�>��<��6���=�`=V����@<�<����$�="��=��=��=��?xT�>����񇱽r�	��9����8>ep=�iH����<;-�#<K��E�L��>�cJ?�+.?��L>��D�Վ�3Y߾X��>��'?x�Y?��	>`���s�=	����*�;�h�>�V�oV��q��D�!�,�V��>���>@_a=�@���w�?J�l?{�6?K�ɾa-Ҿ�_\������>����>I�	>��u�O����?������6~���Z�E>螙��5�;�
>*��=�U�> M��v�=[���@*���Z���=��G>���>z�>W_�>�q�>��9��ݾӄ#�{s4?�"�	�������!��sb;�/�>Ԉ=N�Խ���>�o��bv0����C�;�>Z��?���?�,}?J��)�=���>��>G�N>�mS�E�U��[:��\u>_ȍ���n���;�k��+�$=���<��6��F���`}�R콫^���B����=�VO��K����̾st��������ѽ���z�f�u���;6*�r�q�J�P#���W\�qA�����?v��>�7=���ZG����r'�Rz!>�o����9�	���=~F=���=�Jܼ��ͽI�����о�ͫ��t��}�>�f���~�*�"�-#Ի�a@>[�0?��̾����B�r��=�D)>�-��0J�Ԅ��N���j��.vU?v8?�����[Wҽ�->D9?���>�;>X������BS�>�
/?�-?_��]���j<��?+V�?�NQ?�뾾�ht��!'��?��Y?*?�9c?泌�3���]3��T��>��P?X�)?G�"��T��?���>U��>��%�>��>��>(�a>�Ar�Q]�I��nW�?�Z>�"5>|���;#�Ѥ��`�=L�>�>E�=�>�6���>�侞�1��:�Y�L=����l���>? �A7>NR+>He�=o�*��r��)�����??$\�?��J?PE?�.���˾� ��Ʀ�=}��>���>���=C�0�㏛>�ګ>8RϾ��W��׾�?��?���?�c?�j��Tҿd���e�ž��Ⱦ��>d�=P�1>]'����>�=�ϖ=��;O��=�Հ>%�U>�D[>�<>h̆>�>�����#�פ���o���;=�5�!��J/���]���������ܽ��F�!w¾ez��n�h�o�̽�������������B>7�?�2�>�q<i��=�����nT �������ֽ�}�j���<(Ӿ�ɾ�곾�٧��z���a>��8�?�1ռ���;W�?�����G�>I�:>�Q�=��TB_>]�x>7b�>#x>�\�>~λ>�U�>s��<Kͺ>~���������:�����=/ާ>�|D?t����cy��bS@�9���=>���>�>��yȑ��߄��G�>�%��$��N���}� ��?Yv�>fýD�=��P�]�����=�>��)�+���U�����?�o%�>���>.!վ+i�=%F>��&?{?�s=?��=ˁ�> �6>n�>�	�=}�V>��U>��>\?^v7?,�*?���>�ǫ=��P�z�<��#=��H��2�p�ֽ''�g���Ϩ;we~�b=]y=f�<�=8�>=��ʻ���<$aG=�3?�b�;�6�>@ �>&:��l�Dt@����=@���K>�4�>��#?�]?�)?��:>\:>���>�.Ha��*�>���=��w���`��B�>��>�L�>�rG?�1	?v�t�>C;�>"I>p~K=6ޮ>F$�>u�>���wW��nJ������5D�)#�WD�=�V���M<�z>��9y#��o>4���8�>v2>\�>�R�=�L�=��h>�!����>6�5>�u\=�\�>TM�=N�Q=��!>�_=��.�.]o�au���݁��C���n�;q^�n,��I$����\�(<�3?1&7?;��=�j'>�ɺ�9�¾Ү���/2>�3?�ֈ>��4>��!���o�{���I��:��}�>_�m?x?AI���=��->W�=�V]���=:��=�!C;��->-��<P�>�0�>�?>^�>,Y�i����H���#C����>���aŽ.�?��Q?��J���A�F�T���"���=����Zn�0^��B:��{����qH��˚����=fK?�m�?}_����=,���/,���x�I���Ɛ>���=YL?��>X�>E˽~���㾴�o�G%�<>��=�7�>WG?�x?Ͽa?�	?c?���?���=�a�>'F�>c[?��	??��>��{>��x>r�	=�K8�!�G׋�k�<��dܺ=��>�`)>���<f�=�L==�ا<V=�tp༰��<��s<c�=��=�$�=�$>��?�*?6�\�Ts�:#p!>><,����>�.�<�j>�l�=��ھۋ��ML8=��?��k?�;?��->� ��0�e���Hk>�?�?U�F>��]=Mv�}F�D�Ǿ OR�H�d>�
2�����a�7������5>��?���>��3E�=�(�?�?��@?���¸���9�)U�v��>���>���>R��=ظ�߾8�rM^�Eu�=���A7#��^�>��o�"� ��f�=��.�P��>��>"Ԗ=�q�=G�3�/�<�+�=�c�>�n�>
��>��>�<> �Լ���$:?p�
�	6��3�]O���D=n�.>=���Ͼ�> V>����J\��(���D���>C'�?�?�?uӉ?~���OG����>n�>#��>�qӽ*��2�H��Z��G>���>~Q���V��ͽ�����^�EW������[���������[�9����8$���!��,����q�v����Ө�C��5 ������໾���z|q��[$�Q~��A뾨���?�?:��?��>�|�<WoG�����X�3�G�gS龩���վ,M�/e��������ξ�	���7�@��󫾪��>��Z�,��x�}�b�'�-�R��;D>f+/?@ƾ�A���I��.{=�f'>z�<�s���}���x�`�U?5C9?�}뾎����d���>Ѡ?U�>C�">q6���i���S�>Ԡ3? 4-?���k���ۋ� ���6'�?h��?��M?�cL��dl��qX�ɼ>��\?�5!?s�1?h�=+s%���վ��?�[?�	2?x���U�<������%�>�?��m�|>�	\>b�?A%
>�����L�|���U>2��>m���-K$�Y���;�=$��>��>>��=���=�+X>(d�>��
�3�����>2��`�=-�b\�>���'> V�=�6�=�R)����)��_-���T?��?��%?�T?ׇ�����'4�8e�<��#>+��>��>wC��ҥ>o��>�	�{��)#��w?���?���?pw?<B�?Gӿ��������8��=F%�=��>>��޽�ɭ=Z�K=%ʘ�KY=��>���>o>3;x>k�T>Û<>��.>o�����#��ʤ�2ْ�\B�� ���	wg��{	��y�����ȴ���s�������2Г�s�G�P�� U>�����N�=\Y�>�J�>ߠ>�>;>�}�=�S��Z��­��Ru˾fU�����V	��E���:B��f��W�E����!A��e��J��>O����=��>v/��{�=��>8U�=�NC>@IN>�'>�X!>���:Z��=E;(>�{>�!�=|>��=�섿� ����8��^��#�<�'E?��L�4ɓ�,�3��߾�}��B��>�
?�W>Os&�+k���hw�a��>��`�E[��z���:%����>o
�>�=ؔi�A{�4|����H*�=�τ>Q>�Q�������&��a=R�>�x־��=�pz>�(?.rv?j�5?��= Z�>�^>���>א�=1]J>�M>���>��?�1:?�1?[�>�r�=��_�ϳ
=J�3=�?��(Z����m��!�!��R�<},��0J=�Ww=� <�K=o:=�R��*_�;R��<�"�>��8?���>?��>��9���>�6+M���Ā>;B�hr�>�>��?Y��>}A�>��5>�8_� %þ�N��$�>DA>�l_��x����){w>�%s>ّO?|�1?Yh��!c����<���=��>��?�L)?�>A�>� ��޳��	߿؊�C$�5d�<]n=� -=	�U��lk=��&=���ԍ��s
�=]�b>�ā>zj>��2>�>gV>���>��;>죊=2� >��<�/:�8����x=ι����<����i>�q���v��j!h�և;�Ә���������?w ?C���Tѷ�!w��]a�3۾j7�>�$>�@4?�y,?�,�=FL��c0�@ e�����yW�>F-b?��?(��z��>TwJ�%VY�Tk�>N&=>��d=�XU>�K=1����>W3?N�T?��?X9%��n��M��N&ľ�x�>��<�tS���?�d?������		0�uO�"���m<x��%V�?A���
(���=���a?��,Y�tf4=��?���?�a��+��=9f��|���瀿��K"=���=E�>�>�t��ǻ����m���^J���K>�?�>��x�{�>˒)?��?��{?9�>��?���<�?��7�;C�>�<?�3?.�?|��>'쥼L�T��M�3��=�|�V�����=��t=(^>J9�>|�}>�%��Q��<�S�=������%_k=�SK=�S弮��<��q=��<>vY�>�?z?I'n������۳�
���څd=T+3>���=0�]=�0��z��4��<�?�>�(9?H��>ph�=�������^�������+?��O?	E�>b:�>I	���>��U��NA���?>8HV>Z�z�Y�]��:i����>r� >7���R>6l?I;?/m?g����`/���m�8�'�N?g<q�S�&w�>���>�{�=��̾Pc.�D�q��#a���9��$�+Fg�n:����:>�$7>fkN>�I�=�U>�&=�m��"㽟�=C�T�L��>⺸>'� ?M>t�=l����ᾏtF?��~�����M���K�{v^>���>Z�.<��>�wV��ǋ�YS��Ư�n.#?���?0��?)5r?��W���F>nT��ٲ���= ���~M>Ⱦ�>��>�-0>���w�ݾ^B=d��>1��>�<�������� ���ǿ��k��^|>�Џ�����F�;I��až��N�0D��Kl�(��� c�}��v�CJ��3���������q�?�!M?��%>]Ib=J�Z�B岾����t=?��������쾾�͋��ž�P�����쉵��8����ž���c��>��Y�XA����|���(�꼏�}~?>B6/?�`ƾ2ʹ����1�g=�d%>/ű<�<�r���㯚����cW?�9?�O��*���ὖ�>��?pt�>�%>w(��r?�'�>(:4?��-?)6�;��:��̓��l�?o�?)z/?8 }=-X��!���c��>�\??&�{�wyݾwE�=A�)?��Z?!H�>҉�V���:L�dE�>��j?�����@>3�>�A>�r���H|��SS>�`�����=�!�<������%���?[>���>�`>b���$��q�>4�ݾ�
�_���HB�y���<lf����>��侈E�>'Q>;�u=�@�T����Q��ݒ���x_?�ʾ?��?:?�o����,�z���(>Q�[����>|!�>�ʾa�>�?�<*�Y���@���~�>���?d��?
i?�]��Ͽo옿ǽ���4�O>�=ڬ>';>h�>���B>9*�>5�=]�r=��->M3�>N�>4N>x�z>��>�7>yV��q,���Y1���H5�T6$� %
���c�����O�+���� ����̾͂�����.�%�j%���,�����1��`�6=2`:?�T?�o�><>�S>=����n�ݲ������O"�X�!���{�Ⱦ�^��ay����Kﹾr��=�������>���=ˍ��� 
?C>⽊,>���>���>��>�.�>k�d>z��>k.=���=���=��>�+�<#t�>l�C>娏�>��ZB0�,va���4='7^?f����׾�)�:���{�O6�>xy?N�=�1C�zJ�����$	�>w���U�{��,���^A>���>�݂�1��=�,��O���d��tD=��>�HN>��=+zR�TC���#���>LR׾�s�=�g>�{+?U=z?ǜ7?Ja~=d�>j�{>�{�>>��=��h>�Hm>�^�>I�?6?�+?3?���=v�Z�1P= �!=S<��T��B��\Ӽ�x����< 3�Z{7=��^=�[J;�w=��a=nI���ș;Г�<;�>49?Є�><l�>��8���>���L����lV>/�,���>�]�>
�?�z�>�[�>��/>�^t��Nþ��⾓��>1�@>�^���w�L��0�y>_rt>U�N?[�1?��o�$ d��b =>T�=�E�>�f?�$)?��>��>��\�l�߿U�?s9�V�H<ߑ��i����ľz
�u2!=rK�y�=ը�<���=��>��>���>o�<>A"�>�l�>-�,>�=��X>gi�=��<�����{5��q��Ƈ$����0����;?ӽ�����3�s�2��^&�<2W+?�%?mӾ��=�zȾ�A	�>�	�=P?r�F<)��>���>�ޝ����msE���>���¾���>�hY?�^�>n��t>fOx��݇�:�>*�b>`�޼���>j�<��M!h>��?vi?_�?�g��2��q;����+��9�>��P=��i�mB�?��~??�"�`\�=�DH�#V��[߾&j�=\V�	P����"Q���e��O��������<z$3?��?b]3��r�=B�U�R��� ����;e�=n�=>$��>6��>��¾c�-�E�Q�z��]���6�>��>A��<�)R>h�>�6>�nm?1�?�� ?�k�)R?&{�=yr�>��#?@9?RxG?f�?5�ϻoĽD���Ud>1 ���3��!�"���ɽ���=�`k>۰>�ݼ�o7>|@	>b��<�rP=�s����=X�O=�-�=���=v@>��	>ju
?�*R?wJ�\�<ﱯ�|fԾ}7�<f��>3}�=��k�1 3��7�=I*�>�P?�GA?�D�>T�N� \#�&1L� ���ŵ<��S?�:U?�D�>R�Լl�<�N%�����&6Z>Ҫ{>���0�����,ھ�A���ۧ>���>�K>�a>�? �@?��!?殴�^}5��c���?���Vp}�0$�>�ߦ>r��=��ʾ�H&��p��`��3�jϚ��:M�_&�;��=T>��\>�^�=s��=܂k���>��͔���<��l�Y�>��>���>W�O>l{�=ɏ��b��g?ᗕ����8�����.�*a;*��>��>� �� �>�V�W矿E���,�n����=���?�:�?���?h�<_f½X��>�m
<�Qx>���=���r<�=��ʼ3�ȼ��V����5N�& >-�J>x7�>�t<�gZ��_@о��=»��#�a����:-��������?��3�������hM����.�Ʉ��j&l���g�����=���y��a�� �|��ۋ?�#�?귞>Z"�=�|�F#���՛��7>��P�����߾{�ξ����|��4���3��D<�>U�Gě>�{Y��A��N�|���(�vݏ�Uk?>�8/?�dƾ`Ѵ�����g={e%>�±<=<�p������d�IdW?��9?�J�*���0ὴ�>��?�u�>��%>F&���f��$�>;4?-�-?�����59������]i�?��?��B?fm��_�k&���"�W��>A��>�Y?����b��᪕�,?�Y:?��>�ƾ�V��9�>���>��M?�i���>���>�;[>0����&|����=���� �m=[��=��ֽ�z���'E��߽�>`9�>�(>L����}��ͬ>�7�b��[#���-�L?->O>½PՇ>;�v��>�Dm=�ҙ=Q(#�z���`"��4����6L?~�?~=?zwa?2������Zwս��r���>��j>�V!��,�( �>��9>�,�����	�ze?�h�?��?^?a?۬Z��jѿқ��ɢ��Ѹ���=x�=S}K>?�"����=�+�wt�=DA$=�I>�c�>Ea>�.c>.�A>�ZT>ƆL>�z��q�*�p��JG���C���#�8#��"��O�(�wΨ�L��r��7��Ϙ�����̋��8-�,���u$��A�B�V=�&?H�?/��>���>��F>������оԄ���k�C&��2�����;��<���#��VM��������~=<���?�=>s$>� ?��̽�&>v^>f�S>�x>kQ/>>>n�*>��>�,>H>+�p>�>���>�^<�i�������A-�7����\���.?�-#��4��0�\�������Z?B�A?���>���<����a��>/�=�i������AQ>.��= �0><'^=��>��5=��Ͼ˺�= �)>#}�>M�=��*�� ����z�$��>�S�>��־9�=�dw>p�(?ױv?�.6?�֜=�)�>��a>q�>U��=��L>yP>`g�>��?٦9?�g1?���>�7�=�7a��L=)�8=F�>��U�aM��0���.*���<p:/��H=7;t=N�<7�]=��B=٩���G�;�3=t��>��6?���>���>ȇD��m;�1iE��_�.P�=Lٍ�x��>��>?��>���>��>U�@>�S�;�X�������>vB>L`�3�u����nud>�P�>�_?�Z&?��z�&���H=��=�eq>Kj�>�H?�T�>5U>�DǼ"v��E�� �5~2��1��a��L=�Uo�1x�����޽�R���>�0>�C{>�SX>~�F>C�9>|�8>���>+�/>R=�i�=w�;;=2b4=���=�=��;�h^�0�K=��]���̽t��3L��\���b���g�����?�? ґ���%��c��:�M���3�$?`�!�F/G?�E(?`>�)̾�^^���L�pg�� A?tϒ?��?5h�64>I�;R�]��s�>"t}>�' >�a�<I*=�jϊ�s=�k#?L�_?��>���~�bߛ�����'�e>�]=�8&�>�?�a?�u���H��!��H��H��#t=��DW�!�����"��:�#���" ��&g�s��=<N�>ڂ�?�"~�U�=mW׾�A��ce��0����:=dė=���>H�#>�IU����#�;߹���,��^S=�j�>�I��9[*>yK ?O��>��?��>�C?|P�� h?uϼ���>�:?w` ?��=i`�<�v⽣���aA�nK>gO��-�X�&��5�r��=`!x>�9�=a���R3Z>a�=����[��M�V�c�=E@!=�.>��=�;>_�O>�?S%$?�.�����<�ԋ�����b�F��(?������d�7�ʾ|�����x_.?)uP?�R?��>���`�����_3X>�?��_?��x>�p/=�|>f���l��C�=�p?2|������!�Ѿ�_��*q�>�=�>�m^�bz/>�ڃ?�v3?Y�?x�b�M>�G�O����޸<��置��>�
�>�/�=���+�/�� p���e�>�:��x{�r�w��咽��]>Z�>͈i>�ӳ=>�?>&��;��R�.�ٽR��=�B���|�>�>0�>���=��=�c��	���ݖL?w_���޾�^��=:���->kM�����;�� ��?�����#������������>�	�?�p�?/+??�X���<���>��m�GM�j<6>|���.��|>:�4>��Z<�K�+_׾������>��>q̲<t���g���>�=J���cTX�3"��۞�A��:2��L=��&���V(�3���H�оEsE���R�x)�����[�����$��ȍ���?{Ks?a��=��!�N�R��o� ��~�=/��7n�qʾ!/�$���f�̾�N����پ������5�
����>لY�.A��<�|���(�6я�s�?>}6/?�aƾ�ϴ����g=Z%>3��<g8�D���!�����bW?��9?_P쾯*��%ὀ�>G�?gt�>e�%>M+���#�)�>�84?��-?�켇��:�����gm�?N�?�1?�K�=�jC�����н���>�?pI$?b������@J���U?�L?ap�>� ��G�T�O�a)?�I&?���|�>��>
�a>������3��W�=�r��NȆ>x�<��q�0:�P�1���$�5�O>|��>��k>=���N̺>�SﾵuA���>����=ٽԱ�<$b�>,>���>O�Y>�0>�'��w��ί��V�r�J?�Ѯ?��O?��@?ڐ �+��5A���
=;�>|��>_�w=��R��>{��>�+ݾ7"h�Q����u?��?�q�?dw^?[�d��M�D���驃�RE���]����=fy3>[�K�n�Ļ9->��a>�I8>�>��>J�">z>4�+>��F=�N�=��|���'�[\��A)��tQ�"�#�m��t�|�V��ad��5
�Hy������-�7����q8�B�7�����-������G>�Q>?&�?؀?�̟>��,>�������	Y�r}���[�����F����T���)���Ͼ;@˾��>�8��?�>���=��4�?���j`<=���=OF>�*�=��s>��> �>���>���>;5�>�=�>�6Q>>��=�z�������F6��fO�6wA<hj@?�eM�<���c3��e�h���C�|>��?d�Q>t�%�� ��q�s�G�>�a%�Y�P�k`����r��>�w�>!H�=ͬ�<t�)�N�n���	��Ǒ={�s>m>;�M�ר��K;���`=���>:�ؾ��=BV�>nq(?��u?h<1?�h�=��>~Id>�ݎ>f(�=��Q>K�Y>�1�>X�?U8?-#1?�X�>��=�2[�=��<D�0=2�?���^�﫩�]����!�^�=� 1����<�DV=��&<�V=��o=�������,=a�?��>�3>���>��D����^��>���]���f=N��=��=ޝ?��2?]@?�
�>�����a�qAz<ŷ>��>�#}�|ޑ��bS�J�3�A�?U�Q?��9?���@þa{�������/>�"�>�\#?�Л>ֵ���§�#��mӿ�$�A�!���P���;Z�<��M��ʤ7�-�A���j��<�\>>�>��p>�E>��>�<3>�R�>�HG>�ф=1�=�;�;�;%�E�1�M=.
��CG<��P�����$Ƽ럗����J�I���>�S:�38ټ�?��4?�N����Ѿ��ӽ<�!���?\(�>%��>�?YA%>[C�Ƚc��P���н�L�>�PU?<�n>�;e�q+6>�Z�=^��;U?J��>H�R�q�o����@��0?�>� ?	\�>�����a��t󔿹�g�L>a�=�l���ə?b�|?Up����0>��N�q����j�<o���
�3�q�ȸԾoMϾW/��]����(v1>�'*?T�?̓�{������ ���r�����CF=/�Z�cP >}�=V>���=�;ؽ�i �	¾9��=7� ?�Ó���?t?���>O�?��?I�?+V^>�:?�N�>��>�e�>��=-�����<�D>1f�>�'�����{����V����=5�<���=$:>&XI>�����}0>u���,켝rS��c��}<h2[���L�X�>�	U>�[>ת
?=[ ?�^彞!C��	����*�w<E� >?_B>n�@�YO[���;y�N>G��>x�'?�>qe,=�پH]�E������=�?Q�6?���>��9;��=|�	by��<�=�+_>�����q��P�Ƨ����ҽ �>��d>���=|d>8�?{�%?� ?�E�H�$���5�l������=���=�H�>4�>���ԥ��S�*�O�X J�UQ����|�]�c�=�c�> ĥ>�s>sj=�ߟ=l�����D�ʖ= �F�3+�> �>�(�>�{H>���=Bؾ��澐YJ?��(�[LJ������(�Lל�/��>�_�>�KY>��?��Q��2��㛿6�)�� �>�?��?�?�h���ý<��>�\>1��=�(�=��W����=wH>���>��R>�C�=�������a���`������u��mC��\��Y`��	XQ�[��Ͼ;�����;�,��_}ǽ�Z���^߽��ݾw�Y��w�g��t�?q?����*|���饾�o�?�g�?ܓ�=�H��L1��%����8�=�g���w�(�����)�Mc��+�ľl崾
����*�a�*�8W
�L/�>����!��a���4�����8�����>pvݾbj�r�F�Ȱ���>��>�5&�Ǝq�1���ǯO=@u?L�$?(�������^��<:Q�>�B?Ň�>Oϥ�h�����>��/?�a:?���Uކ�g"�c��?~�?�D?`r���&�˵n��a�]�>�Tu>�̗>c���P�J�Pp�t�C?��}?��?{�����о2��R?��X?o��7r>��?���>=�>�+��G�.�ξ%����>b��=�>�<�7��s�����<,�G>X^�>����L̾���>�����]�W!�/��$�0={���y�>D#Ⱦ�%>Dh#>�<>6�(�(��/������:U?  �?J�4?J�R?��
�� �,��L�����>���>�)m�&ZT�7-�>I��>IP���i�A�۾�.?��?��?��Y?�U��пg����s��& �@S>�ԗ=�:>QU��0@>��/>,�F>%�O=��>�D>Ѥ�=�~>b�k>�!>�6(>W]~�_h#����	˞� �7���)�(���o��1;�:km��,������>�����齖��A�f�j.��~���� 5�����a>��K?�?z�?
��>o:>u�4��^6��Dֽ�&6�y���ԓ����-&��ě��)�������G�>�˻�I]?-/>EU;�v?DZ ��/>\3�>��z=ĵ�<��>"��=(�s>��>���=�!>TT>+YҺ��~>�ԋ=
���π�5�:�x2Q�5�=<n�C?��Y����Z�4�!�ᾲ������>G<	?��X>ߪ&�
����u����>��8�5$f���ӽ�W!����>"��>0g�=�jϺ������q���=䯀>�	>�!�������1X�=�	�>�־��=�gw>@�(?u�v?FG6?֝=r��>T�a>޺�>D��=��L>�Q>jψ>7�?�9?k�1?c^�>�B�=�^`���=&:=��>���W�?���$��p-&��!�<�S1���F=�yq=r�<`=p�C=KBż��;���<S�	?��>���>]9�> �q�L�4���a�<����ܽ����5ʑ>�	?�?/#?1?x��\E���uӽ`=n��>İ�>��H�lhk�I��=�:�>l\�>c?��[?�Y=F Ӿ#��8�E>v��>��>J�?��>�=_��=Dy�F�տ^��S�T�K+�8����v=\]|��@t=��%>��a=�g��X��<���=��>�N�>���>1xg= �>���>�/>��5>��3>{06� +y<�oQ��7)=�ܽٓT<]4����)������R���X\�ڳ�a���j$��/0���?�m2?��սǤ.<!P{�_��-ɽs�?�v�>���>�8�>��̼3�!�z$`�p�>�io���>v(5?+˫>i�l��)>�C=>5�=�U�>\�>�4<��Ľm�Ͻo��0a�Mp�>�?j�M>Ŗ~�)�[�Q��(�u!}>J )={�%�d��?�d?���~��]K%�H�E����N�N=cB�y�U������ ���7���@7��n�Rh�=�q?�1�?8~�:��=$�羯N��wu��Xɾ>�<�ο=�v�>��>�a<��I��R� �赪��q�ǥB=<y�>Iq�;��?��?�?�j??��?V��=�?▂=b�?5]>iq�>l��>R�>��O>cҠ=JM���v��k	��U��j�:O؋�#�%=f��=  �=?$��8,>幑��(�=����.�"=�D�=�f�=�8T=��=�_>��!>�*?��$?-d,�!ʰ�L:��n�+�1��=ݗI>?gh>�&`���r������'>1~�>�y.?̤�>f-�=� Ծ�+Ͼ�L����=��?)q+?���>�&t���U=FS޾�r����=���>�k(��d���3�@Q��m�߽{��>�Qo>��=x_O>�)�?�'?,:?��<���9�)���fU=̗>[b�>sv�=���A��6W������L�F�CXm��/�*�>�a>�F�>@�N>��=�������%B½��=�_�<�Z�>��>u8�>�>��=p3���U�3D?ԧe���@�6�9A�[��<Q5d>ޱo>��<�(0?d��겆��E������?xX�?�C�?t�?�ǂ��ޓ;�>�g��+�<�.�=��ξb�;�v۽�M���=�"9�e�V���ƽc��=Y4i>B�<�˥�SKp��4���I��B^N�Sk�����_�v���Ǿ󔭾b6%�`(��@��vѾ>�P����x�8�Qe'��@-���}��G��u9��� �?�n�?�k+>VnV=��b����ξU�=eA����?�8k����e>���ӹ���� �����"��/���I��>\6?�I��������'��j�<-=>�>sX��5�����O�T�����>� y>����O��]��ܝ�=Ö{?��?x�~��!����O�>&��>̺�>��j>Ȩ_�ʞ���Z�>U�d?YK_?�.�={ʋ�����{Ƹ�6��?�O�?�I?�梾�HM��x侠���d.�v�=_J�=y��fZ,���,�c�1?O��?�J??G*f�f�r�=9����L?��Y?����h̤=�P>/�>�K����6=Fi���o�g�Q>��=׵a������b���.u=�5�>R��>�M���_����>7���N��H�0��%�����<�~?���I0>.i>�A>P�(�7���ω��A���L?��?I�S?�h8?Od�������=�=&��>�>��=���$О>���>\X辱vr���q�?�J�?���?WZ?��m��Aο�$��*�ʾ����=V�>Sք>�<{�>�F��va���=Z������>�|�>��:>��=@Y
>��>����,����"����\$���S��(Y¾� ��3�E�� ����$ľ\Ə�5��~f�E����w_�-�<ꯄ�a�7>���>)�?��>py�=���=�P����9'ᾷ���w���9 �s׾�M���%s��I��B��D�F�@�о^�?wH�=:�>`�?��=|�Y>��>��Y�`�%>��#>�oe>&�=q$F>%�>�|E>�,�=�d�=Uz{>�ч=�(��o���p:�X�Q��D�;��C?��]��l����3�2]߾ڨ��\�><�?ӧS>B�'�ⷔ���x����>_�G���b�+0˽"q��[�>\��>�{�=l[λ����w��$�
*�=a��>D4>\�h�<���Y��|�=�-'?��Ⱦ>U��Q�5=N?D�p?C�S?*�5>K�>��0<��?��>��">4� ?�D�>�.?��R?�C?�n$?��=���j����<ТG�dۼy\��P����
=�@ȼe�n��E)��@�;&]=�q9>	ָ=F;<�Ev�w�=I*�>{9?.?�?5*=���267���=�ϧ>��
�F��>��>��[?Vn>f�r>�yz>��=����ФP�h��>���=h�*�~�M�U���->��M>_M~?�@I?:�j>�7�=��g9$O�-��>{?2l?d��>���>fB>>�O��п��<�T�>�s��K��=Oƌ=�����<@��=��O�ː������r>~W�>��>n�O>��/>z�}>?G�>x�=�5=e�>ߧ3�<�<X(U;�Ž�,��?�>������W�$7���� �@=�	�=��>�q>�e�=>6?\�??�=͘j=�kW�Z��v8��
e-?8�'?�V�>��#?�y>H.$��Wb���̾�S����>��}?���>�a���<>�0������>C%�>rq>�[d�᧾�J��gQs=���>֭�>;�> �����:��64��Ҿ��>s�ٽ��ν�=�?��C?#A3�:���W�*�K0�t9c��N7<���r`���ؾq�P���e�. ���-����D�	>+&�>���?59@>}�m��:h��촿Qi��X��k�{>mD�����>���>B���ylپ�F���N�^����`'�=@j?>���>���>��
?�[?(�#?�?�2���1�>E
�&�?O�>� ?.�?]&�>Wג>'3�>$P>�ӎ=��'=r�O{�;�鼼�=>�5�>X�}>~J�� �;_f�<i��L�d�=��=�+;�<x����y;���=��?��#?�潽�'��Լ�+��X�<�<#>]9n>�K��5Q�n�` L>��>2Z0?� �>'T�=��Ͼ�.����k+�=�F?��/?�(�>�/[�r��=m��C�v���t=f�W>���5�������쪾���K߁>[��>XW>A��=�@�?	��?�3>tWᾴ�n��v��YJh���'@Z>��
��t��PS�=�Y��Bi��×�����99b�d²���\�151�GR����q>Z�O>�5x>�dp>XQ�<��>۳���<>>�M�=��>�~�>6��>���>��>L\໚i*���I?
u��0���o���ϾY����> �@>_����?�	���}��ϥ�@q=�5�>*D�?9��?�Id?�D�O%�RI\>xnU>�>�*<t�?�+�v���Ӽ5>[��=�"y�Cw���g:cXY>�{>E�˽�g˾m�⾮02��D���9���ȍ���c�Z�	�ǡs���⽊]����Oڣ=ކ0�qOH���v���G�eT=$.#<��e�Ā[��o[�?ԏ?J�Z?���>��> �@���3�}о8B�>c3&�U�8����糾��&�<�Ⱦ���t�+CL�&�;�U������>&�Y� A��R�|���(�����-�?>�4/?�`ƾaδ�\��?�g=�^%>~��<�:�����ͯ�����bW?��9?5R쾒*��x�ľ>e�?u�>�%>*���4��%�>�84?��-?�@켹���9��7����l�?� �?�??�P�8�A�^���?�KF?޾?G��>K�����̾���?��9?�8�>1��>7������'�>B�[?�
N�e-b>�}�>��>��~���]&&�����-���9>��� �q�g�P�=� �=���>(�x>�]����Ş�>0e��R���I�c���3 ��<1?�g���	>�Hc>�U>�%�mm���w������4sM?���?SP?(7?I���`|�*��7uv=D�><��>���=�)��f�>��>t���eq�i����?Y��?�5�?1Z?�`j�Ϳd蕿����īž���=��=S>ϓ����=�����������#>��>;�>$n�>�B>�jw>bP->�?����&������ܜ���G�����
�PQ���!���^�������z`���r�An�tS^������l+���ԙ���>���>5��>h&�>�g>{ ��ю��{��3���������?�о��$��E	�cǊ��"�sj���;7t۾G �>ex�;��ݽ���> :<���<u�>�=�<�ӽc3>�t�=�|)>X>(J>:c>�#>��>�Pl>I��=��r��@q�nC�!����\B>bH?�R��>����^A��Sھ�����ͽ>RB?É>mm��7p�OME��H�>dT��Ն�A!����>�&pd>�z�>V�>�[����G��u���.��n,>e��>a�E=b��?���.��$�=�s�7��}���j>:�?�ho?�54?�u�>�و>�&�>r���jM�~fM>��>��Z>zr�>�T?���>��U>8>֝r�*��1Է��N&�0�0����
���nO$��h)�v���>H`�<͌���s��=x�=��=!�=q�&?��'?���>L�>׺����L��W���6Խ�+����>�m�>E2?,V)>X�F>J����"=���)����>����o��8�+��;�o>疘>+M?�0?Cvt�)h�,��>��|>�د>�]�>��0?�F�>%g>v/�����i���!?G�\Zg��Eh=�T=�&��8�ǽ(J⾔c����۽2׾􋐽���>\��>HU>�>]�d>�o�>ޗ�>i
�=�>��R>�U�=L�3>��Ҽ��<ZiC����=o��tM��B=�̳�uǈ���J�����=��<�;?}$w?��?&��j$���HB�i��@>�sU?z#??�7,?P��>�q���p�/�}��ƾ*��>2o?�V%?G������i=�>I^�>p�>�-�=��$� aR=ɟ��L.	>D>�:�>`��>h�=���C��j=�@ാ�>�>o'�>Π+>��?v|c?Gj*�P>׾�=#�P�L�'n4����y������4����3���1�S`������d��#ϒ=�>։�?���>�)P��&��I̟�p◿�˯������l>�m=?2������P�6� �]t2�?;�O���T�=K0=0�>;�?��?h�{?;K+?��?�8�>������>�Z�>�Z�>�	?�4?��<>s<e>4%�<-K}<�� �K8��Uٕ<og��n=�=��=�� >.�;��~���2<V��<�	�-J0���=���=HC=E52>9�9>�*>a�?�L?J����Ԭ�*����j ��g=i�>�F;>N�B��~r�ۀ3>& O>���>��>ʭ�>W�>>�G����T�Ѿ8VJ>x�#?�B&?���>�
+�����ϾD�<�=j�=j>.�����ϒ���=F�m>�k>�>#?6�R?)�F?�(H?�
�=�B�K:��p�;�o����zT?��>`4q>(����0��0��Ñ�I�M��ch����S���/�B����=-�>�Q�>���>�Ni>��ӽ�Y�)w2�Vf�$!I>�Z�>��?�<>l�=P�H�~ݾv�3?�17�W��*�y���˽��>��>�QX�f
?���{I~�ࡿ@�Ͼ+�?�V�?�[�?[�c?�Vq����� �O>�E>Vm��w'��o���g�=�0=���=��<Q[��he�o�p��8�>K��>��Ƚ0澽�����Z�g����`X�_�2�־��e�ب:������<,�t��|ü횼�M�t��툾 �;�ù�%�x�d�ц������?r�h?ё4=:w�=��v�7,���b�>�XM�N�m=����a����������a��8=þq���B�P�8����>AZ��ۑ��W{��S)�+ꎼ�@>.�-?҆ž�y��H���x=��$>�0�<�q�꼊��B��k�y�V?T:?j"��Q��]�޽/�>�q?E��>��%>d���PG�+��>�4?u�-?)�Լ����ҋ��ƅ�ӻ?՝�?54?;Y)�$�Y����K�k��>4X
?���>��Y�[���H��W? �9?Q��>�f�h�e�+����>�^1?M-.���q>P�>l�W>�9�;#ʾ]e��=��b�����A>9s�=��W��<��]��q��=?��>�T�>.�������>2:�X�N�c�H��������Ə<v�?���?">�i>�D>Ϻ(�����͉��,���L?:��?��S?�h8?�_�����ӎ��2��=u��>Ԭ>��=�����>���>g�|r����?�I�?���?�QZ?��m���ȿ9Ց��$��LϾ�P1�=*�=��Y>�yn��=�7�<Ul
;�+��Z�>mЇ>�fE>k\>�>6>ʈX>�>����j#�����L����OF�.��;F����97���׾8Z�CKȾ��ľ�2�V���֐>��K����x�o������B>�b?.Y�>��>�\>v�l=����+y���;����g	����z��~����[�_����ƾ�w;󏻽NZ��s��>�Z�<�V>	��>�/�=J�u>;_�>�*���B�˾�=��F>6J�=�)>YV>e��>��]>�y3�|�{>�F�=������|:��9P����;��C?�L\�t��p�3�"�߾<?����>��?A�T>�'�(Y��ҏx��t�>/I��`b��˽}p#�P��>!{�>��=S�ʻ(����x�|��?%�=A�>�
>*�z������m�<�=<�"?�������o-^>�;&?z3F?�?���=d2�>~ɼ>���a�pü�n;�=���>�3?�s&?��>֠�>�5=��"�e�����=�s�����?Y�p��	�����=�_������*Լй��V�@=�Ȁ;�y���s���Q=.��>rjU?{��>/�>��'��,�
O�p�����>G�'=�k�>Fڧ>�b?��>s��>��4>p�=�o���g�(��>�}[>�J[����������v>λ�>�J?WJ?V���~E�7	=dPU���?.
�>V&�>,�>K�>��P>��mӿ�$�J�!��)O���;�<�h�M�(2�7A�-�X���L��<�\>�>ۅp>�E>ů>�<3>�R�>�HG>�ф=��=�<�;��;��E�A�M=:
��FG<�P�����%ƼJ���A���I���>�d:��7ټ�@�>��W?�3@=���;B���־F���VQ�>��?�-�>T��>s�="���3�"	N�����&?��r?a��>oͽAE#�<�=�s�ɽ���>ܚ�>5��>�
.>��ӾX�ݾ���=<D�>'�$?r�>��㽓�E���n��Y� ]�>��2�!�Ѽ55�?g�??��$��K输A)�1�Z�3N��]�!XԽ����{���:��J{���@���8���Ѿ�y=��>	d�?��X>�}1>��;��K��� ��Aq�K-0>�*O>r��>{�S>�?4�
����V ������g�7uv�p.�>;�2>��>_�
?xjB?��?u��>�8(�n�?�ۡ>�6U>�B�<Mz�>4�#?��'?+��>���>m>���=b��6-9���罐�L��"ɼ���P
>�=3��=�����)�<D�<�D�=�Y�=��K<p�6=��>L�>>��=�R?�W?Tc߽o�`��+)<-꒽/}�=��(>�.�>��f<�*���x���>��>��-?;��>Լ�=~-����޾���=�[?@h6?�g�>�'u={p=� ���(UP=�;>[�e�5n��v˾�m��#���k�>
�]>�>��'���R?-tc?�?:��4����㣿��l�?}ξb�>�[?�^�>8�<�Z��O�AAa�k���R���=���-�J��|A$�\/�=q��>C�a>�S>x�j>�}�=��=	�=Kw-�rB�=�6�>�?ϵ�>o��>, @��Ͼ��H?Ƈ���������Aʾ+߼�1 >[�I>����?19�:�}��㥿Ц9����>�P�?��?ܫa?�iD�&���T>R=W>�>��#<Q�(�aj�����B,>9�=@���f��x��;mI>D]l>-⽂�ƾ�⾢,�3����r��`F���ྙ��M���\���Ü�g��j�B��<㾆ݽ	ҽ��A��Q@�Čc��������xH���?�˔?�)0>?��=DI�q��3��'���Q�U���ta��o��������>L�^��:�6��C������W�=��9������%�h��z���?P�s?����js��f0���>��&>z�?�?R������������>�Lh?��2?��	�aC�Z�S=������>���>��}�y��=ͺ4>J$M?"�7?*�<�qg�*� ���$=`
T?��? 85?� ��|�9����u$���	?_
?
��>!|��wؾZ����H?tx6?�:�>-�m�r���=�?��\?��=�b�=��>֟�>�'��d�)_�='5�������\>�q�<�J��{߾)�=��>��>{�=��¾�0��^��>D�$�N�#�H����$���ˏ<�?���6>�i>�H>ɸ(����a͉��"���L?���?��S?�k8?gb�����g���We�=��>
Ѭ>{��=U��r�>+��>+c��tr�Q�1�?#I�?y��?�]Z?�m�I��Õ�k
Ѿ�誾�w�;f1w>�tb>��=.�2=�dV�cb���""��>#�>��>���>q�>2AT>��>�6��k��i���y
���`��(��m��p���?x����g���7 ����_���ɼ�!�;
7q�b$��q⊽��Ⱦ0�=�U	?�k�>KM�>�l�>F�2>K]�����s1��9�T�P��w�S!��2̾�)j�;��9�C��zR�1��<I0��-�?6c�=+�<"��>��=�jz>���>A�=V��>ra}>m�w>���=�q>��	>��>�@>���Cb|>�z�=j��一�R:��|Q����;�mC?S]�豙�W�3��޾�䨾=��>ӑ?��S>�'������9y����>ϾG��Bc�L�˽��#��J�>@�>�F�=VV���A�}rw���㵶=e��>��>o_�w��������=ܲ>N¾Ro�?ɇ>�^3?`�c?�K?[�4>���>� �>OX>��=��>Z�>i�>c�?��4?�2?M��>\>�m���;�=$m>*³�*����i<�w=�����<>T̾�X=�!�=vM�<��罼�>n�]>E@�<�c*���?��7?pQe>L�>�偾-'��	�$���6�>�s��|�A>}`�>n�?vt>(��>��>B���ιʾ�T�u�>sgx=�)j���R�\��=֟�=��H>L	�?��^?J�RYe=��>Ծ����0>��0?tvW?���>0��>�F�=b$��������X�"g�P輽]�N>G/;=5_�Q�R������݈��F.��r��	A�>䋫>���>X��>+4�>zq�>���>�,�>0_ >Bj=L9M>Ǚ��{���ʔ��X�:
!=�U�ї��&H�<O�}<�f�� ��KX׽�����=��#?��?� �ļ�����KN���oo?��D?�X�>1�"?K >�1��:��;���2.��T�>f�~?���>���$ҟ=���J����>�P�>SA4>�S'��.F����sѵ=dԐ>�9?�9�>��H=��Y��z��仾P? L�=:�q����?�?�Q7��ξ��� �t�2-,����>,�l�>r��^��/���b��{	����\��z��>wJ�>7��?,�
:��:c��������`Ǿ������K�?���>�vȾ�ھnxN�]_��L��ežH�>�5�=YW�>	9	?w�>Dt?@M7?�I#?�u	>���>AB>��>
J�>oA?�`�>�Y�>�Ñ>���>���<��!�p潙埾����B����*&=$R>�{h>��=Y�= �ԍC= �e=W���rE<�̻>ߛ<�! ;>/�=F�?sL#?@|���Խ��>6�	��=>�#>��>�*��ئ=F���k��=�U?kM?�F�>Q�=��1�����E㾾�3=��
?x�,?+X
?��>}�=����1K�?7�>G�>��̽�#��.������7���X�>g@>��=\�>�D�?��k?PU�>�ڭ�L�t�Qܔ��GK��^�l�ٺ�1�>�!?O�B>��AGl�{=��ޢ��7n��v0��դ���<&�?=��_=/1 >��>	ߧ>@�
=�cm���,�|�ʽ�B��� ?���>�?�&�>�cA>�K���q2���J?+����R��ा:JȾWd��[>Ab>�b����>�ƽM�t�����&<�k��>{ �?2V�?��f?�RF�7I��  Z>>#N>;	>iI=�"<��,��r}��	I>	��=��^��*����&�]es>F�~>n+ͽ<?˾�Qо��<D����N�t-��Ѿ��p�b���-7��(NｹF����ڽR���������!����R�%�^䅾�>��cSr��W�?�[�?HQe>�-=I)������ᾁ��=A4��[�@˾#Uy�㖾��پr���_���C"�8���*����>ӉY�FA���|��(�����;�?>�5/?`ƾ�ϴ�]��y�g=Oa%>��<�:�*��������cW?��9?R�j+���Ὂ�>��?�t�>��%>�(��*5��&�>/94?e�-?�E켾��#:������]m�?N�? `@?�xK��B�T���=�L9?r?i��>@����˾Rݽ]�	?�*8?Ӈ�>�E��m�������>�Z?��M��`>�{�>�ٗ>¿�op���C�{Ŕ��4ͼۡA>ϫ�Z.�݂a�f<�r�=�+�>�<{>�^]�[��^��>D�$�N�#�H����$���ˏ<�?���6>�i>�H>ɸ(����a͉��"���L?���?��S?�k8?gb�����g���We�=��>
Ѭ>{��=U��r�>+��>+c��tr�Q�1�?#I�?y��?�]Z?�m�I��Õ�k
Ѿ�誾�w�;f1w>�tb>��=.�2=�dV�cb���""��>#�>��>���>q�>2AT>��>�6��k��i���y
���`��(��m��p���?x����g���7 ����_���ɼ�!�;
7q�b$��q⊽��Ⱦ0�=�U	?�k�>KM�>�l�>F�2>K]�����s1��9�T�P��w�S!��2̾�)j�;��9�C��zR�1��<I0��-�?6c�=+�<"��>��=�jz>���>A�=V��>ra}>m�w>���=�q>��	>��>�@>���Cb|>�z�=j��一�R:��|Q����;�mC?S]�豙�W�3��޾�䨾=��>ӑ?��S>�'������9y����>ϾG��Bc�L�˽��#��J�>@�>�F�=VV���A�}rw���㵶=e��>��>o_�w��������=ܲ>N¾Ro�?ɇ>�^3?`�c?�K?[�4>���>� �>OX>��=��>Z�>i�>c�?��4?�2?M��>\>�m���;�=$m>*³�*����i<�w=�����<>T̾�X=�!�=vM�<��罼�>n�]>E@�<�c*���?��7?pQe>L�>�偾-'��	�$���6�>�s��|�A>}`�>n�?vt>(��>��>B���ιʾ�T�u�>sgx=�)j���R�\��=֟�=��H>L	�?��^?J�RYe=��>Ծ����0>��0?tvW?���>0��>�F�=b$��������X�"g�P輽]�N>G/;=5_�Q�R������݈��F.��r��	A�>䋫>���>X��>+4�>zq�>���>�,�>0_ >Bj=L9M>Ǚ��{���ʔ��X�:
!=�U�ї��&H�<O�}<�f�� ��KX׽�����=��#?��?� �ļ�����KN���oo?��D?�X�>1�"?K >�1��:��;���2.��T�>f�~?���>���$ҟ=���J����>�P�>SA4>�S'��.F����sѵ=dԐ>�9?�9�>��H=��Y��z��仾P? L�=:�q����?�?�Q7��ξ��� �t�2-,����>,�l�>r��^��/���b��{	����\��z��>wJ�>7��?,�
:��:c��������`Ǿ������K�?���>�vȾ�ھnxN�]_��L��ežH�>�5�=YW�>	9	?w�>Dt?@M7?�I#?�u	>���>AB>��>
J�>oA?�`�>�Y�>�Ñ>���>���<��!�p潙埾����B����*&=$R>�{h>��=Y�= �ԍC= �e=W���rE<�̻>ߛ<�! ;>/�=F�?sL#?@|���Խ��>6�	��=>�#>��>�*��ئ=F���k��=�U?kM?�F�>Q�=��1�����E㾾�3=��
?x�,?+X
?��>}�=����1K�?7�>G�>��̽�#��.������7���X�>g@>��=\�>�D�?��k?PU�>�ڭ�L�t�Qܔ��GK��^�l�ٺ�1�>�!?O�B>��AGl�{=��ޢ��7n��v0��դ���<&�?=��_=/1 >��>	ߧ>@�
=�cm���,�|�ʽ�B��� ?���>�?�&�>�cA>�K���q2���J?+����R��ा:JȾWd��[>Ab>�b����>�ƽM�t�����&<�k��>{ �?2V�?��f?�RF�7I��  Z>>#N>;	>iI=�"<��,��r}��	I>	��=��^��*����&�]es>F�~>n+ͽ<?˾�Qо��<D����N�t-��Ѿ��p�b���-7��(NｹF����ڽR���������!����R�%�^䅾�>��cSr��W�?�[�?HQe>�-=I)������ᾁ��=A4��[�@˾#Uy�㖾��پr���_���C"�8���*����>ӉY�FA���|��(�����;�?>�5/?`ƾ�ϴ�]��y�g=Oa%>��<�:�*��������cW?��9?R�j+���Ὂ�>��?�t�>��%>�(��*5��&�>/94?e�-?�E켾��#:������]m�?N�? `@?�xK��B�T���=�L9?r?i��>@����˾Rݽ]�	?�*8?Ӈ�>�E��m�������>�Z?��M��`>�{�>�ٗ>¿�op���C�{Ŕ��4ͼۡA>ϫ�Z.�݂a�f<�r�=�+�>�<{>�^]�[��`��>\;��N���H�^����0i�<��?U��K>�/i>�P>�(�:���щ��?���L?6��?�S?yj8?oV����GΧ�뚐=���>zŬ>���=4��3ߞ>e��>V��or���Ӕ?�G�?���?AUZ?K�m��P�� ���:�:�ž��X=��>>���o7=����9<�=��н�Ǳ>C٪>�>���>�>>�L�=<�=>q̂��(������#��C��<ZǾ_�4��J������U�� ����%�����B�@�+=\�����f�,j׼�����>��?M�>s�>�dA> �,>����'�8r�U뱾՛���50��h>˾�<w�[�(�Ka�����QͲ�8y��?�`@<�h�=9s�>�J�M
>k�>��}=�v$>�B>g>�J>>s8>�
M>i�%>�X>[�=y�x>Mk'>b�����~�E�"��%Z�LT=)>T?~Z���B���:���#2��b`�>52?���>�C�����=F�����>��:�ܽ�	�tu��G+�>|��>B3K>H����?�=	Kƾ]�Y=k��:��>��u>f�=@ҫ��d˽Dc}>F#?!��W;��>�S ?�vB?��6?��>�#>�4.������� �b��=<��>��?�� ?��-?9ZB?b?�>�c�=4����&˼o�-=�z�4���5�<o��<e��<pE�RC>$�����=׽K>�+>E>���;���=L>g�>k�Q?.��>���>�ֽުE�"~;��p����e>� �y��>�}>�?�r�>z�>�-]>DM����k]1��V�>f�!>-Ft��ك�� ��[�>M�>S�?�;?Y+�=�˾��#��=��>`Z	?�0?�?�c�>��"���tӿ3$�!�!����o����;S�<�S N��a:7�-�q)��G'�<>�\>J�>a�p>7�D>ז> ?3>�?�>�,G>Dv�=�!�=R�;�;E�<�M=�3��WJ<�FP��;���kɼ�ԗ������J��@����9�ؼ�?�]?% )�ጽ f�����諭��>R��>>�>O��>���=9l��}U��GA�G�F��|�>��h?Ƙ�>��8��S�=�8/�#��:7�>T�>�>�b���������o�<P�>��?ou�>~��K[�_}o�ָ
� �>����v@��2�?b�?�+Q�����OBD���.��T����>X��>	����!�ӶG��>i�!]N�ۤZ�����c�>��?Ɨ�?3�3�g艼�پ? �������^��=��>B"�>@�>f����[L������Cs����>aEJ>�+�>5.�>�$?c�X?Mt$?�k?��8�ѽ�>�L���>�Q�>�Q?�?D��>��>���>�XA=V�옽�VL��KU��`���#�=��`>!�1>Il��p�=�<U=�t��:νT���=�W����J��3)>G�>Z��=�=?�n?]޽/��q�=�ҽ���=E��>Sv7>��=V������=��>e� ?�w#?�? �=}���+�����ˁR��Y?%�K?��>�"_>���=�	��OǾ.���pa>��)>5�L�Xc��Orξ��s�V��>�m�=��w=�}/��d�?0�_?��=����{���:��v���.�>��>�Ғ>��>�����r�)I��-���έ��T�v�����(��"�3>��=�X>�F�>'�;>��O>y�/�n�M=�����'���H�w��>�A>Wv?�[O>8@/>-v��M>�i�I?"���?������y�̾`��m >��=>�� ��?���-~�=���Ci;��r�>���?�!�?�zd?ӑB�"}� �Y>�Z>�>�9<��<����!�:�/>8��=�u�/����@����_>��~>�����ɾv��}
3�'�Ϳ�A����<^w�-���gp�FL��ϭ�沆�/i�/����E����Z�s�O�cҺ�1ئ�P�������9k��Ã?#�q?�\�>ݚ=L'�bw�ɏ����=oB���<�C,�?���1�)� �D
�TM=���E��x�2\����>�Y�~@����|���(��ŏ��?>B5/?�`ƾnʹ������g=�^%>©�<$<����	������bW?��9?�P�>*����o�>v�?3s�>��%>�'���3�.&�>�94?ޫ-?�V켽���9��ލ���l�?� �?3o??��P��}A����2���(?�<?"��>Χ���ϾM]�?D�:?ė�>5����#y��{�>�XZ?��J���^>A`�>��>�� �i:��Z�y�����ʼ?/>��:���'b�)8�bu�=�_�>�jz>�wa����4��>7B���N���H�/�����QU�<�?)��6>i>�@>/�(����Gω�~)���L?ߚ�?D�S?l8?%_��$��;���,��=���>�Ҭ>���=����>t��>�e�Lxr�u��?JJ�?���?\Z?��m�Vaпn����Ծ�o���[�<��<��5>��|��S�=އݽr����'�Z�=��>�ϱ>qa>�2\>���=���>e���Z�h	��(쯿J򃿢V<�#�	��5'���㾔蓾�1�ZѾ܌���	�  ���#!��3S��٬����;�s���e=m�?;��>J�>��C>�j>�{��6��P>�$é�%���^���待����pp����R�$�b�T��/�'��_O%?���<?��=|��>%�����>�ݐ>]�=�ZD>�EV>��=��>�LA>� >��='�>:�=r�x>��=�4���9��y�:�A�R���;E�C?P�\�y�����3�Ǜ߾1ҩ�`�>@�?WS>O'��}��L}x�!��>�F��lb�b�ν݋%�V�>��>Xֽ=�����w����ʔ�=�;�>t�
>>li���Ty�}ӗ=�W	?њ&���B�w9>��F?�W�?	W?F�>���;i�4>I��>�Aڻ�8�>dL�>篋>fW-?R�U?:�?;��>%�o=�W�s��y��=>�&�g�!����}zS�ͳ��B7�=�8E�����=�ݾ=�?�=��;�R�F�N�`�d���?@�d?�p�>(�>�m��W_u�_� ��W�=딬>F���;�=��?� �>�?-��>|rc>VW��t����x"����>�9�>z�8���u�V�>ò�>���?�?��������Ӳ=��@=��$>�Z>/�}?kz'?}��>"�>�����譿��F��od�����^���C�>�1��+>��>N�������y���>L��>�J>��n><�>�'�>9��>v��=��n>�~>В>�>�$��?ɽ'd���Q�=ݢ���<�-=��0�Y��	_=�_!=��,�J"j=�?	T3?E1�U�}�Q�����{��Y+?f�?�>3>�e�>ɔ>"���e�E���+�&X"=J�?7�i?�c?�*.���?=����i�ǽ5H�>�?;3�>���y��t(x��h0=�>�??���>�d�n�d�E�h�މ����>��D�f���?yc?�9,��2��Ǽ8���U��#���S>���=�'پk5-���Y��O� "8�e4M��V�DPR>g�?w��?5o��m��>�����������̹����!�r�����>�(}>i����S�	w��&�����`���ȼ���>L�x>�˰>E?%�d?��H?�?2?��p����>�&y<8�#?���>�c?�w"?U?W��>&��>�=�>LBͽ}�J�$~�=�e=B�->��?>�z<>%��R�V=��(=� >�.=y�5�9=1!2=rW��B�=1>sF�=�?-�#?X�H�V7���Q�=��	�ƈ�=<�_>5�=��X����?��<�;�>o?e$?$��>F~�=}������|��Ѽ�O	?�!>?a��>}�=���=���+䳾<@�=1�|>��6�&������{]������1�>.W�>�.ĻB��>��i?��%?��,?͚���1�Qޟ��Zl�T�=�;w�?���>.Y�/<a��c~������#��RǄ�S�B�MEԽ�R>ʆ�� �=-��>-vu<�3�>��=��=���	��T��{�}�D��>:�?��0?��>�b>��������I?�h���e�i����Vо���[�>��=>"����?_��B�}�����0=�Q{�>H��?#��?Z:d?m�C��L�\>V>6p>�.<8�>����d��b�3>���=Ty��ܕ���;��\>�Jy>;�ɽ��ʾ�S�F��淿.�x�@�͹7���
��	f���ݥ���`�H���b�;Zj;�"x�)�þ#P��ػ8=M�6�:�9�0kŽ4�����??�?0��>UV��,=���Ǿ^_о�b�=TUd��َ=�~:���s绾W���;$������(P��M��@�����>axY��>����|���(��c��р?>�=/?Eƾ`ٴ���G�g=q[%>o��<N-�k������y�
��bW?��9?Q쾧��9X���>Z�?{�>��%>�,��2�'�>�64?Y�-?������6���㓼kk�?���?�x@?��ܽ��9����'E����?��?��?�Q��ܾ��&���?��P?�ǲ>�8��b8m�������>�^a?�MN�P�+>�>��>�y��Z��_2<�>������k�>��m9�2��e;��F�|�=P��>��R>Ɍw��L��`��>\;��N���H�^����0i�<��?U��K>�/i>�P>�(�:���щ��?���L?6��?�S?yj8?oV����GΧ�뚐=���>zŬ>���=4��3ߞ>e��>V��or���Ӕ?�G�?���?AUZ?K�m��P�� ���:�:�ž��X=��>>���o7=����9<�=��н�Ǳ>C٪>�>���>�>>�L�=<�=>q̂��(������#��C��<ZǾ_�4��J������U�� ����%�����B�@�+=\�����f�,j׼�����>��?M�>s�>�dA> �,>����'�8r�U뱾՛���50��h>˾�<w�[�(�Ka�����QͲ�8y��?�`@<�h�=9s�>�J�M
>k�>��}=�v$>�B>g>�J>>s8>�
M>i�%>�X>[�=y�x>Mk'>b�����~�E�"��%Z�LT=)>T?~Z���B���:���#2��b`�>52?���>�C�����=F�����>��:�ܽ�	�tu��G+�>|��>B3K>H����?�=	Kƾ]�Y=k��:��>��u>f�=@ҫ��d˽Dc}>F#?!��W;��>�S ?�vB?��6?��>�#>�4.������� �b��=<��>��?�� ?��-?9ZB?b?�>�c�=4����&˼o�-=�z�4���5�<o��<e��<pE�RC>$�����=׽K>�+>E>���;���=L>g�>k�Q?.��>���>�ֽުE�"~;��p����e>� �y��>�}>�?�r�>z�>�-]>DM����k]1��V�>f�!>-Ft��ك�� ��[�>M�>S�?�;?Y+�=�˾��#��=��>`Z	?�0?�?�c�>��"���tӿ3$�!�!����o����;S�<�S N��a:7�-�q)��G'�<>�\>J�>a�p>7�D>ז> ?3>�?�>�,G>Dv�=�!�=R�;�;E�<�M=�3��WJ<�FP��;���kɼ�ԗ������J��@����9�ؼ�?�]?% )�ጽ f�����諭��>R��>>�>O��>���=9l��}U��GA�G�F��|�>��h?Ƙ�>��8��S�=�8/�#��:7�>T�>�>�b���������o�<P�>��?ou�>~��K[�_}o�ָ
� �>����v@��2�?b�?�+Q�����OBD���.��T����>X��>	����!�ӶG��>i�!]N�ۤZ�����c�>��?Ɨ�?3�3�g艼�پ? �������^��=��>B"�>@�>f����[L������Cs����>aEJ>�+�>5.�>�$?c�X?Mt$?�k?��8�ѽ�>�L���>�Q�>�Q?�?D��>��>���>�XA=V�옽�VL��KU��`���#�=��`>!�1>Il��p�=�<U=�t��:νT���=�W����J��3)>G�>Z��=�=?�n?]޽/��q�=�ҽ���=E��>Sv7>��=V������=��>e� ?�w#?�? �=}���+�����ˁR��Y?%�K?��>�"_>���=�	��OǾ.���pa>��)>5�L�Xc��Orξ��s�V��>�m�=��w=�}/��d�?0�_?��=����{���:��v���.�>��>�Ғ>��>�����r�)I��-���έ��T�v�����(��"�3>��=�X>�F�>'�;>��O>y�/�n�M=�����'���H�w��>�A>Wv?�[O>8@/>-v��M>�i�I?"���?������y�̾`��m >��=>�� ��?���-~�=���Ci;��r�>���?�!�?�zd?ӑB�"}� �Y>�Z>�>�9<��<����!�:�/>8��=�u�/����@����_>��~>�����ɾv��}
3�'�Ϳ�A����<^w�-���gp�FL��ϭ�沆�/i�/����E����Z�s�O�cҺ�1ئ�P�������9k��Ã?#�q?�\�>ݚ=L'�bw�ɏ����=oB���<�C,�?���1�)� �D
�TM=���E��x�2\����>�Y�~@����|���(��ŏ��?>B5/?�`ƾnʹ������g=�^%>©�<$<����	������bW?��9?�P�>*����o�>v�?3s�>��%>�'���3�.&�>�94?ޫ-?�V켽���9��ލ���l�?� �?3o??��P��}A����2���(?�<?"��>Χ���ϾM]�?D�:?ė�>5����#y��{�>�XZ?��J���^>A`�>��>�� �i:��Z�y�����ʼ?/>��:���'b�)8�bu�=�_�>�jz>�wa����4��>7B���N���H�/�����QU�<�?)��6>i>�@>/�(����Gω�~)���L?ߚ�?D�S?l8?%_��$��;���,��=���>�Ҭ>���=����>t��>�e�Lxr�u��?JJ�?���?\Z?��m�Vaпn����Ծ�o���[�<��<��5>��|��S�=އݽr����'�Z�=��>�ϱ>qa>�2\>���=���>e���Z�h	��(쯿J򃿢V<�#�	��5'���㾔蓾�1�ZѾ܌���	�  ���#!��3S��٬����;�s���e=m�?;��>J�>��C>�j>�{��6��P>�$é�%���^���待����pp����R�$�b�T��/�'��_O%?���<?��=|��>%�����>�ݐ>]�=�ZD>�EV>��=��>�LA>� >��='�>:�=r�x>��=�4���9��y�:�A�R���;E�C?P�\�y�����3�Ǜ߾1ҩ�`�>@�?WS>O'��}��L}x�!��>�F��lb�b�ν݋%�V�>��>Xֽ=�����w����ʔ�=�;�>t�
>>li���Ty�}ӗ=�W	?њ&���B�w9>��F?�W�?	W?F�>���;i�4>I��>�Aڻ�8�>dL�>篋>fW-?R�U?:�?;��>%�o=�W�s��y��=>�&�g�!����}zS�ͳ��B7�=�8E�����=�ݾ=�?�=��;�R�F�N�`�d���?@�d?�p�>(�>�m��W_u�_� ��W�=딬>F���;�=��?� �>�?-��>|rc>VW��t����x"����>�9�>z�8���u�V�>ò�>���?�?��������Ӳ=��@=��$>�Z>/�}?kz'?}��>"�>�����譿��F��od�����^���C�>�1��+>��>N�������y���>L��>�J>��n><�>�'�>9��>v��=��n>�~>В>�>�$��?ɽ'd���Q�=ݢ���<�-=��0�Y��	_=�_!=��,�J"j=�?	T3?E1�U�}�Q�����{��Y+?f�?�>3>�e�>ɔ>"���e�E���+�&X"=J�?7�i?�c?�*.���?=����i�ǽ5H�>�?;3�>���y��t(x��h0=�>�??���>�d�n�d�E�h�މ����>��D�f���?yc?�9,��2��Ǽ8���U��#���S>���=�'پk5-���Y��O� "8�e4M��V�DPR>g�?w��?5o��m��>�����������̹����!�r�����>�(}>i����S�	w��&�����`���ȼ���>L�x>�˰>E?%�d?��H?�?2?��p����>�&y<8�#?���>�c?�w"?U?W��>&��>�=�>LBͽ}�J�$~�=�e=B�->��?>�z<>%��R�V=��(=� >�.=y�5�9=1!2=rW��B�=1>sF�=�?-�#?X�H�V7���Q�=��	�ƈ�=<�_>5�=��X����?��<�;�>o?e$?$��>F~�=}������|��Ѽ�O	?�!>?a��>}�=���=���+䳾<@�=1�|>��6�&������{]������1�>.W�>�.ĻB��>��i?��%?��,?͚���1�Qޟ��Zl�T�=�;w�?���>.Y�/<a��c~������#��RǄ�S�B�MEԽ�R>ʆ�� �=-��>-vu<�3�>��=��=���	��T��{�}�D��>:�?��0?��>�b>��������I?�h���e�i����Vо���[�>��=>"����?_��B�}�����0=�Q{�>H��?#��?Z:d?m�C��L�\>V>6p>�.<8�>����d��b�3>���=Ty��ܕ���;��\>�Jy>;�ɽ��ʾ�S�F��淿.�x�@�͹7���
��	f���ݥ���`�H���b�;Zj;�"x�)�þ#P��ػ8=M�6�:�9�0kŽ4�����??�?0��>UV��,=���Ǿ^_о�b�=TUd��َ=�~:���s绾W���;$������(P��M��@�����>axY��>����|���(��c��р?>�=/?Eƾ`ٴ���G�g=q[%>o��<N-�k������y�
��bW?��9?Q쾧��9X���>Z�?{�>��%>�,��2�'�>�64?Y�-?������6���㓼kk�?���?�x@?��ܽ��9����'E����?��?��?�Q��ܾ��&���?��P?�ǲ>�8��b8m�������>�^a?�MN�P�+>�>��>�y��Z��_2<�>������k�>��m9�2��e;��F�|�=P��>��R>Ɍw��L��4��>7B���N���H�/�����QU�<�?)��6>i>�@>/�(����Gω�~)���L?ߚ�?D�S?l8?%_��$��;���,��=���>�Ҭ>���=����>t��>�e�Lxr�u��?JJ�?���?\Z?��m�Vaпn����Ծ�o���[�<��<��5>��|��S�=އݽr����'�Z�=��>�ϱ>qa>�2\>���=���>e���Z�h	��(쯿J򃿢V<�#�	��5'���㾔蓾�1�ZѾ܌���	�  ���#!��3S��٬����;�s���e=m�?;��>J�>��C>�j>�{��6��P>�$é�%���^���待����pp����R�$�b�T��/�'��_O%?���<?��=|��>%�����>�ݐ>]�=�ZD>�EV>��=��>�LA>� >��='�>:�=r�x>��=�4���9��y�:�A�R���;E�C?P�\�y�����3�Ǜ߾1ҩ�`�>@�?WS>O'��}��L}x�!��>�F��lb�b�ν݋%�V�>��>Xֽ=�����w����ʔ�=�;�>t�
>>li���Ty�}ӗ=�W	?њ&���B�w9>��F?�W�?	W?F�>���;i�4>I��>�Aڻ�8�>dL�>篋>fW-?R�U?:�?;��>%�o=�W�s��y��=>�&�g�!����}zS�ͳ��B7�=�8E�����=�ݾ=�?�=��;�R�F�N�`�d���?@�d?�p�>(�>�m��W_u�_� ��W�=딬>F���;�=��?� �>�?-��>|rc>VW��t����x"����>�9�>z�8���u�V�>ò�>���?�?��������Ӳ=��@=��$>�Z>/�}?kz'?}��>"�>�����譿��F��od�����^���C�>�1��+>��>N�������y���>L��>�J>��n><�>�'�>9��>v��=��n>�~>В>�>�$��?ɽ'd���Q�=ݢ���<�-=��0�Y��	_=�_!=��,�J"j=�?	T3?E1�U�}�Q�����{��Y+?f�?�>3>�e�>ɔ>"���e�E���+�&X"=J�?7�i?�c?�*.���?=����i�ǽ5H�>�?;3�>���y��t(x��h0=�>�??���>�d�n�d�E�h�މ����>��D�f���?yc?�9,��2��Ǽ8���U��#���S>���=�'پk5-���Y��O� "8�e4M��V�DPR>g�?w��?5o��m��>�����������̹����!�r�����>�(}>i����S�	w��&�����`���ȼ���>L�x>�˰>E?%�d?��H?�?2?��p����>�&y<8�#?���>�c?�w"?U?W��>&��>�=�>LBͽ}�J�$~�=�e=B�->��?>�z<>%��R�V=��(=� >�.=y�5�9=1!2=rW��B�=1>sF�=�?-�#?X�H�V7���Q�=��	�ƈ�=<�_>5�=��X����?��<�;�>o?e$?$��>F~�=}������|��Ѽ�O	?�!>?a��>}�=���=���+䳾<@�=1�|>��6�&������{]������1�>.W�>�.ĻB��>��i?��%?��,?͚���1�Qޟ��Zl�T�=�;w�?���>.Y�/<a��c~������#��RǄ�S�B�MEԽ�R>ʆ�� �=-��>-vu<�3�>��=��=���	��T��{�}�D��>:�?��0?��>�b>��������I?�h���e�i����Vо���[�>��=>"����?_��B�}�����0=�Q{�>H��?#��?Z:d?m�C��L�\>V>6p>�.<8�>����d��b�3>���=Ty��ܕ���;��\>�Jy>;�ɽ��ʾ�S�F��淿.�x�@�͹7���
��	f���ݥ���`�H���b�;Zj;�"x�)�þ#P��ػ8=M�6�:�9�0kŽ4�����??�?0��>UV��,=���Ǿ^_о�b�=TUd��َ=�~:���s绾W���;$������(P��M��@�����>axY��>����|���(��c��р?>�=/?Eƾ`ٴ���G�g=q[%>o��<N-�k������y�
��bW?��9?Q쾧��9X���>Z�?{�>��%>�,��2�'�>�64?Y�-?������6���㓼kk�?���?�x@?��ܽ��9����'E����?��?��?�Q��ܾ��&���?��P?�ǲ>�8��b8m�������>�^a?�MN�P�+>�>��>�y��Z��_2<�>������k�>��m9�2��e;��F�|�=P��>��R>Ɍw��L��S??��־,ޒ�i<�~ㅿm��=�<���>���=�}�>	]>p~c>����d��F�����޾��&?�O�?�Ԓ?��>:��%[�C�'�-��=?��>5��>��/=�JǾ��|>ø?����2:���˾y0?M��?1��?8�Q?Z�r��V׿����D��������=��D=@�->��^���^=1�+>�^;��-���>�q>���>�ӕ>�0>P�>YK>>�&�����{�����EA�� 	�ʖ�FK7���S�w������&ľ+
Ӿ�tȽ�S�白>�B�:x��;�;�6��>C�?dc	?92�>�]�����>{��e�F������b�YM�p���幾x��������T���'ƾv�p��0Ӿ.(	?��<��a�����>�ā�e�=L�>bs�>��>�!>l>t��>+�>�>�>؅�=lK�>�����,y>���=:#��� ���@2���O�QԼ�6?��R�������6���辠;���O�>
?fE>��,�⓿�{�lk�>cf� �j�?5��m���Y�>�z�>��=m�k_ü��y���,��=v>�>Ӥɼצ��¦���=�O�>$gϾ�br>~�>'-?d�m?4�A?{�>�$�>8�{=��>Ry��/�>��>5(�>��4?XFI?gM)?���>�L�='��=1hb<!T��j-��#U�����:����<���Ϗ����!��P����n={^=�N��[2�<��=�U�>�o?�E�><���H�����GR����0�4�>'�>��>�~�>^-?��8?��=�]=�X۾j����M>����>�>�>�q���i���^>'��>&��>�?$Y8?�������<'<�u�>FQe>	�2?m�,?K`>F`�=�ҽ���ڽ���횾���6�=���y%�=����N�m�ѽ�%��tþP~W����>4�?�#�>J?/>�A��w�����>��G><PI=
8>q��=+N�=/bz=/k�<M͔=�F�=��i��B&=^�=w@�=򓽸�j���3�P�^�ͼڽ��:?T�?����<����[��ޡ����B�?�!]>#r?�Q	?�듽���Q�X�c]M�WSھ��?p�?�Y4?����8�>�>�J�>'�!?`�L���P>bh1��q���:��tߝ��O�>�?��x>v���� \�m�����9���>/��;ĩ�(�?fvQ?;�B�hI���I��cT�"�9�u8>��>��l���i��#���T���Ѿ�;�4X�����'��>��?�ۖ���˽���w��=ê��v(�VH��O�>�-?��*>
ҹ����XA���D�Ug�������=��$=�t�<��?��?rT?#�?΀7?�nZ>�_�>[N�m�?�M�=��??��>�6?%&?4p?�S�>�z;O���ӕ��̙����n>�i>�}=�>{ݍ=�T���=l�ټ�Q\�op:=���&�=��=���<�>`��>�`Z?fҽ�[��ú>R�R����X�!��>�N �����=���>Aa?D?��>Ƥ��$�����:۾	Rb�[p?��O?料>a�� >1��<]Jj�q����U<�J��B��>��0�'����^u>�@�=�3>�>]>� �?��?4�"?��=�F�,�O�U|��<������8̼'�>d��=`���1��a��<���R�2���fz��o��睕>`c2>��=��W=�u�>[� >�DR�Qkj�:�$=0�#�� 8>���>2J?�+�=��=����+�)��N?Gݟ�$9��}��d۾��?<��>��U>���?-���\�x�������@�X�>�{�?4��?6�l?}���^	���l>�}X>ad>��y=��8�%�'�@A�9>���=@3g�Tם���f=�go>?hv>���ڈľ��ᾆ�K�T���Xt��Ҽ&4�����������I���?
�n�G���\ڽ�>���|G=h�-��AҼ����bP���䬾ɡ?�L?�]�>a���Bf���Ӿ<��Ɓ_=fO��*�½���e�3�S��������/���pF/�q�7�K��U�>�G罼Ҋ�+8�O0@��侨s�C�G?���=\|E�_�1�(��>8��=ē����!��ɟ��ۛ�KD�1�P?7f?�����=��s������"V?�>��=cS\>9������>�U?���>�ɯ��f��X>���/Ѽa	�?o��?�$@?0Xʽ��H�4�Ǿ���Z�>_�?���>���B�ܾ�k��`?!�?�B?>Ѝ��v��������>�sn?_��Z>��?�#�>�d۽7E]�aO��z0��6�H��=a5�*`.��e�F$����<�j�>�֨>0|¾5����6�>�B��O�K�H�]����x�<��?���">�ii>�,>T�(�����[Љ���ȧL?ȧ�?��S?�K8?�9�������� �=��>j٬>�8�=�4���>��>�p�iOr����?��?޺�?�CZ?n�m�v�ֿ����܊��_����=��=R�X>�5ɽ�M�=�dǼ�FG=N0�=a�=��>���>���>⥜>~z>�>p����B ��M�������.�,���v����C��Uy�T��#~������[;����Z�{ʈ�Ĉs� A�� v�}�����=$�>b��>�!�>�������>��&����4O���.�i/c�|Oݾ�:���g���A�=ё���v��y����jоZ�?Q��=ᵕ=�_�>&�/�QL�=�,p>GY�>k+�>*�h=-~=*��>	 ?w�>��ּ��K>Z����x>���=o��������}6��[U�1�s�X�B? s]�~��9�2�J�ݾm���T�>N�?/MR>C�%�Q��� x��9�>�'p�H�`������&��Y�>K��>߄�=�!&�n�+��;{����߾�=z�}>�Q>͌����<����=���>�	�,�
>,��>� %?�Gq?t�8?�ɟ=L��>}+W>Gf�>R�=�g4>�~s>�>s�?�[<?��*?-��>��=*_���<L=y.F��Ӛ���׽�:޼Gz��& =^�h��)f=T��=���;(-.=�1=�<{�޻�m<��>w�k?37�>����@�=�߾�i��,�"�:BQ=�]�>Q��>��>E��>�$?"rx>fO�=1�w�d��"X&���>���>��d�]Rg�&x�=em>q�>��E?
�1?�Mн�;��kO]=�A�&;�>,�>*��>�ۑ><�>��#���d?ӿ����p�^�ʼ�<H[1=b�+��##;,�0�q���޽���6\>�ϗ>.��>Z�K>��=K�>˪�>�\>LS=3��=�8�F~мۏ���fp=�tq<rM=�'�mqD<����3/�ڪ��������j'Q�'�ü�m?�H?-夽tҽޚd����<ɴ�|x�>1.�>{� ?,3�>��=�=��^��C��=@��+�>�NY?��?E�G�=�kǽ�<X�.�>�ʰ>?o>8D/���w�V��^�(=���>�Y?U�>�5I�|lM�F�r������z�>E=����J�M��?e�H?#d��^��!7�2-�R�R��u�>����ZE��,(�o� �]B	������P�]�ݾ����ѥ	?�N�?~<��|�����f����L��Ж�[��>o$�=�&?,G�>y޽�f۾Z�5�i喾�捾���Cc�>�:�4�>� N?�0G?��A?��>��*?��轆^�>��v�}�-??0�>O�?&x-?�D?��?�0?��<u_��� ���|���>�"=m�>T�i>F'�=� 8���<b`=�]>ܫ 9�ct�:s<�'�<��o>Q9>B>)q>E��>ݏ&?&���	˽<��<�Ƨ����ew>�>"ve����o�E=�>�|�>dx:?���>�i="��q�������:�V��>ne?cޮ>��=��>q
2��ǿ�b��6��=����^W�����D���k����>��!>�x0>}^>�@�?��>?Y�?��ܽ�Q)�ey���1���μ�!<�u�>�M�>]c�=�<ξR�3�
�o�_�c�-�./��&�=�ː="%�=�)>�qD> ��=�:>z*@=N��%�׽X��;�/�S�>'�>��?�fX>" �= �������I?���?h�A砾ikоA{�E�>J�<>��j�?��<�}����F=�I��>ʄ�?���?97d?o�C�-���\>;OV>0�>e�/<��>�"��Mh����3>(!�=�xy�*"���;G ]>2Ky>�ɽ��ʾ�+�0�H�춼�{:���5\=fEB��Z�����K��������I����=)�־����E�����z8=O�S���9��ؾ������?,H?Z��>+�,��H�֖	���%�k�9���n�=��Ѿ��׽Ɵ�=�(��Ӿ6���]]��%�B��L�?$���0���}���n7>E�P=�F?��<%��BB׾��>�iH�����_"��*d��螿;�,<�Iz?g�4?�����w�@�~ѳ���,?�s?�=�\r�~�a����><�?��>-7�>#�o�N,��������?��?&�d?��l�8�~�*�ƾ�9��Q?�)?�e�>��d��$�(�w��>��d>���(@��ޔ����\?6��?�z����N>R#�>!l�>.��=ƿ���Y">�ى�Q�u�"��GՔ���^���=	��V���%>]P�>�����S??��־,ޒ�i<�~ㅿm��=�<���>���=�}�>	]>p~c>����d��F�����޾��&?�O�?�Ԓ?��>:��%[�C�'�-��=?��>5��>��/=�JǾ��|>ø?����2:���˾y0?M��?1��?8�Q?Z�r��V׿����D��������=��D=@�->��^���^=1�+>�^;��-���>�q>���>�ӕ>�0>P�>YK>>�&�����{�����EA�� 	�ʖ�FK7���S�w������&ľ+
Ӿ�tȽ�S�白>�B�:x��;�;�6��>C�?dc	?92�>�]�����>{��e�F������b�YM�p���幾x��������T���'ƾv�p��0Ӿ.(	?��<��a�����>�ā�e�=L�>bs�>��>�!>l>t��>+�>�>�>؅�=lK�>�����,y>���=:#��� ���@2���O�QԼ�6?��R�������6���辠;���O�>
?fE>��,�⓿�{�lk�>cf� �j�?5��m���Y�>�z�>��=m�k_ü��y���,��=v>�>Ӥɼצ��¦���=�O�>$gϾ�br>~�>'-?d�m?4�A?{�>�$�>8�{=��>Ry��/�>��>5(�>��4?XFI?gM)?���>�L�='��=1hb<!T��j-��#U�����:����<���Ϗ����!��P����n={^=�N��[2�<��=�U�>�o?�E�><���H�����GR����0�4�>'�>��>�~�>^-?��8?��=�]=�X۾j����M>����>�>�>�q���i���^>'��>&��>�?$Y8?�������<'<�u�>FQe>	�2?m�,?K`>F`�=�ҽ���ڽ���횾���6�=���y%�=����N�m�ѽ�%��tþP~W����>4�?�#�>J?/>�A��w�����>��G><PI=
8>q��=+N�=/bz=/k�<M͔=�F�=��i��B&=^�=w@�=򓽸�j���3�P�^�ͼڽ��:?T�?����<����[��ޡ����B�?�!]>#r?�Q	?�듽���Q�X�c]M�WSھ��?p�?�Y4?����8�>�>�J�>'�!?`�L���P>bh1��q���:��tߝ��O�>�?��x>v���� \�m�����9���>/��;ĩ�(�?fvQ?;�B�hI���I��cT�"�9�u8>��>��l���i��#���T���Ѿ�;�4X�����'��>��?�ۖ���˽���w��=ê��v(�VH��O�>�-?��*>
ҹ����XA���D�Ug�������=��$=�t�<��?��?rT?#�?΀7?�nZ>�_�>[N�m�?�M�=��??��>�6?%&?4p?�S�>�z;O���ӕ��̙����n>�i>�}=�>{ݍ=�T���=l�ټ�Q\�op:=���&�=��=���<�>`��>�`Z?fҽ�[��ú>R�R����X�!��>�N �����=���>Aa?D?��>Ƥ��$�����:۾	Rb�[p?��O?料>a�� >1��<]Jj�q����U<�J��B��>��0�'����^u>�@�=�3>�>]>� �?��?4�"?��=�F�,�O�U|��<������8̼'�>d��=`���1��a��<���R�2���fz��o��睕>`c2>��=��W=�u�>[� >�DR�Qkj�:�$=0�#�� 8>���>2J?�+�=��=����+�)��N?Gݟ�$9��}��d۾��?<��>��U>���?-���\�x�������@�X�>�{�?4��?6�l?}���^	���l>�}X>ad>��y=��8�%�'�@A�9>���=@3g�Tם���f=�go>?hv>���ڈľ��ᾆ�K�T���Xt��Ҽ&4�����������I���?
�n�G���\ڽ�>���|G=h�-��AҼ����bP���䬾ɡ?�L?�]�>a���Bf���Ӿ<��Ɓ_=fO��*�½���e�3�S��������/���pF/�q�7�K��U�>�G罼Ҋ�+8�O0@��侨s�C�G?���=\|E�_�1�(��>8��=ē����!��ɟ��ۛ�KD�1�P?7f?�����=��s������"V?�>��=cS\>9������>�U?���>�ɯ��f��X>���/Ѽa	�?o��?�$@?0Xʽ��H�4�Ǿ���Z�>_�?���>���B�ܾ�k��`?!�?�B?>Ѝ��v��������>�sn?_��Z>��?�#�>�d۽7E]�aO��z0��6�H��=a5�*`.��e�F$����<�j�>�֨>0|¾5����-?����_�d����nH��U̼r1�S?� [>��>M$?he>pWC�F+���Yn��IϾe�B?�.�?AG�?�#?����Ҋ�AЉ�Ⱥ�>�	?��.>�H�����8>0�?'��u�b��1��H�/?r��?j5�?���?�w�'�п%���55��wؾA-;�Cg��z�>����^�=�0�>L?>
>�K>��>�-�>��>�=Z=�F>w���� ��˙��<���`�B �����%"��|
�����x�����	���a �i���8�����Z������,���;�Ps�>J��>��?��?��C�oo�>@Y��/
-�ϝ���߾��2��3� 4	�`x$��y�����=`��K�¾�)m��$��70?�.5=��=2�>ڷ��W�>�> �k>y��>:�!=�
>(��>k�>���>q�~>��=��ʼ�(>�p =O��\)���3��M�ک��r�!?�L�mt�>�;"羥a��n:�>�?h�">�[/�����K�v��P�>���hw��g���H,�DH�>�t�>�
>�=LEv����6�&�~7�=ɬ�>��=�.���@r�S߽Z�=^��>��Ⱦ�">p�+>O<?o�?<�{?_�>�>~#��a�>N�?>ל�>F�j>"K�>�?#�Q?l�?���>�o">�9[������ >�派ϙ����lT�٦/=���=�>l��=O�;>f�C���e��{�=�r+�;�2>Mx>B�>O}:?��C>z��<�1���,��q���&���¼s��<z�|>{H�>D�>�&?6�>S(<��@z��9���>1��>� r�G΀�d��=��>$�>���	?H�&?>]�>^�����?��؝��ep>�g?W�>D�`>�e�>�O��j��*�ſ���6"^��)��0<�^ͼ!�=��|�L.��@����[�����>j�>���>�k�=ൽ�D�;��={>�>�W>?l==�$�=ˠ>��>B��|��=H�+:�|{�A\������� H�����*a�h0]�� Ž'v%�+��)GA?���>��̾:y�qu]�8&&�+��y^�>d%?���>-�(?�!��tY��
v��mB�.y��_?�܊?��D?[˾E|?����� >7�>�����?65�=]����$)�W���(?uc?v}�>������8�WƏ�>>�[y�>�/i�>M�����?�rN?	��������X�3���,��mžA��� �=-�=�ξ�MQ��7�e�q�N��=�
?S�?Ld�d���>��'���Rp~�:����sn=��X>)�>���>
3�=o�|
�&Xﾄ�m��ಽ>,"�0��>��?0�K?`�~?��>��;?��-��;>=�<u0�>�-�>�4?4?�S?Id?_��>�7Ƽ��c��K���z���l�;��*��<��>�1T>��.=�1�=�4ҽ�-�	��=n�Y����=��.>��=,m_�;�:=�b>�/?�'1?Q7�08�����<x�v����t�c�c�+>v��=�Ծ	0 >�%Z=��>���>�Φ>������s2��9�R�H���$?H�b?�=�>
���n�R>I$��b�n	�r�>TՀ��B��0�/�P0̾ӭ｜>�D>�+f>�kc>��q?�t?D�?��2=�
w�2�%�U>'� 8H<��?>-�;>@#��2��xT$�Too�hh���)�i��./n���^�pC�=0��>	]C>��x�љ�>z�>^%<�,����=!���Z>�Ψ>�R�>��=� Z>Cݡ����9�h?��׾�M'�Y��ㄵ����=c_�<�>��#>ʭ�>�>����7���cT�
�>͆�?��?��?�G��s��q�T>�>&��=WD�<�
�(����9m�>V=��������?��T�=�>�>�����Bþ�W�i�E¸��to�3����޾�+w���!�/q��a�<U�K����mC�dI��j�"�ƽQ�J��	� �������Gq�7!�?UAF?��>�H=��z�'��;b��!�� r��)��Z�(�қ�طW�q=ɾ�,۾��?	�+ɾ���>
�/�	����*��RO��=�����=HZ\?o���������]��<��b;�9��	!�)�ɾ���
ؽ�h?�i?S"�����Y��[н��	?Z2�>D��>Ɣ'>���$"�>wk]?\G(?���[b��}���nv����?#z�?~#8?t�C�ǓT��b��/�-<ߚ>��?���>"E���2���7x� ?8� ?�>X�!�Js|��Q����>Pc?1���pl>��?���>'=+=����Z�<l��a�
����<9���Y *��G���(��T�̼��>S�>K�� =��?
� ���E����4I�$�̾�>h??�be�?ٞ>�?~��c�S������怿]L>9�J?�N�?�n?F�^?1�}�Z�Y�*qV�2�=�ĥ>�]�<L��=�2�>Qg�>�_�����#�kw�>���?;��?��?�5���̿������f�����="BG>�e�>X���>��>C�=$e;~�<>��>}`�>b�T>�
>8��=�>@���C'�҇�������T�����.�Y���FL� �?����]J���ʾ0E���a7��E�Um���y���۲��x����>j>�>v� ?}�>�8�=�\> �������(�m��������ݾ�(~���߾�=���`��#��M!��f���	k!?�=�K�< d�>9>�2�>�,�>�W�=ֽ�=�D>8F	>Ď]>�L&>�x=aˌ=��I>Q/*=&�������X*�n���x'���?�Zq��NL�R ����L�~�>���># �=��(�����ءw����>Q�x��#?����:̇��y_�>}�>�8>����q����\�G�.�Nya�.>�UK>�{��I������Ǥ	>s��>��о�>�8�>Ai-?�{?S�6?�̰=z��>�VZ>�N�>���=`SU>�h>��>*"?�o4?�+?ʧ�>�[�=�g�&��<s�)=��9��aJ�#׽/���q8�3��<�9�`S�<�Zh=��8=�Ɉ=��3=J�뼇$�K��<j}�>��?��e>�|�=����A�&�w�q���h�=\ I>�N�>�?A�?�?��3>%�<��\���Ͼ�s��t�>վ>4&|���h�
�8��"�>L��>�>#?]�,?NL=nvu��Y�5��>/�=>�7?���>�B�>�j>�%�����Zjӿ�$�v�!������R���;a�<��-N�i�,�Ś-�0����q�<�\>�>�vp>��D>m�>`63>�O�>IG>��=���=5��;��;O�E�1�M=����F<"�P�޲���Ƽ��������lI�-�>��0�ټ��(?��?$?���|����2�w9��LX���>辝>,�?	E ?0iD=�$��&K��A�
ѽ���>�3{?��<?�l���J�>]�X�>�f=��*?�E�=�o>�^�
ؾ�V*��f=��>��.?'�>�J�dv�u���o����>�1G�|��Җ?��X?�}�m䋾T,D�.�X�f�2�&#�=��<~s�����R��Yu?�7�������f�=�&?���?dྻ߽�9��8̤��q���o4>�u�=�T ?{P�>韋���s=K�^#��4b�$>��>� �4?��f?��6?f��?��e?��0?�Y>��>������>A��>TK9?�]B?B y?��>Nq�=P:�k ��d�����MT�D9���E	>Fl�>��>�������c}->�nv>�����`�=j,�>Л�=��(>��>d�>0A>���>Y?��6�ƒ	�����^l������=d>���,,d�(��==�> l�>��?�<�>��;=yؾ^�Y5�g׎=2�?C�:?GԹ>�Fἣ��=���ꅾ/Y�ia>�G�o����3�-�����׽�W>�$D>b�>:��=�-h?�� ?y�?R��;��"�Y�=�� �fGS��"���jŽ'׵><7O>q;�����V���:�p�*�"����Z���q>���=�X�=���=��>3>���B�U��}S�wg>�%�>'�>I5)?���=����������&3�?d���9�n[����0�����t�6>��D>��>���=aҞ�
㌿�෿�Z��ק=2A�?�4�?QǙ?��/�@���ua>���=ꉽ��B>>Y�⽇�̽�>�O��V��!���ʢ*>��=�>n��~��!B��7N���0��K"t��V���}���b��F��A��V�I�Jv���➺T,���Q����:H����x
�𔾾�O徹���ȍ|?��\?�H>�w�=zD1���_��ZQ�L�޾�3�ԗ��-轮o���k��#��&�ݾ�$������徑��>F�X��ё��{�R�(�s����=>E�.?��ƾ.������߻W=h�#>xV�<�﾿]�����
Q�W?�j:?�뾳W��'�O>�
?>&�>�S*>K������9��>q�3?��,?ύ� ���F����e�7��?A��?UQ0?��/�f�F�ŕ����M��>��?�B�>���������̽7?��%?���>���	�~�һ�=�>dna?螎�-�g>�?F?z䪽w��7�;��H��}���W\<49��O��'R��U֨��ң=���>��I>ڸ����%ѫ>H9���*3�U�@�����B������8��>s����i=Y�>���`�2�~Z���{�럽_�j?≲?��T?�,6?�u�NM	�w�i�s6>�ʆ>P�>Y�
>�Od=a�4>�,�>[��P�^�+��V6*?�:�?�g@�r[?A$^�9yԿ�	�����م���U>9��=I��=2�w���#>����j�� ��.?>���>�>=�>[89>��>�� >�v��
a!�C����$��O6����� �)������c���&*�਍�F�������!��P�\����p׽�D����% =L�>���>U�?�Ze>=v�A������b-<M;ľ�g$�8�2������Ǿ�s��h��`���߾N�$<йʾ���>/bL���=�%�>}VO=�7�>}��>�k�=n��=�O>�s>}�&=�5g>��,>���<�>�>t/>xV�>���=6������LRK��f���=��?�͚�����"1����!���v��>�~"?��>p���ӓ�ok��S�>�+=�|c��ܽꯌ=�W>l�>�%�=	�Ҽ�3=^����~۽�;>:�>�b">=��u�a��븽P��=5��>��վ�]�=P�z>��(?�w?5?�\�=���>�A`>��>�C�=H`I>��N>��>��?<g8?i71?	 �>�=��^�$�=��@=��:��]�aq�����- +�d��<	/���P=�$�=�/	<��Z=D=7=4�ȼ&2t;_�	=p�>��9?�S�>o��>��<�hd<��K���"��� >�;�-��>�#�>��?z��>��>�G>O�/�"¾wIܾ�]�>ʒE>��]��v�_஼M'|>i�j>�P?U`2?t��S_��=�3�=�Ʈ>��?U.'?(^�>�L>������	���ڿ��<����\�
=�p��lj���@u�����[9���1#�E*̽{�=�/>X,>��t>�0�>h>q>q//>h��>��>�>��> �(=��ۺ��	��能Qx��h=��`��aO�jG�n��af�IY��$I=p�ҽ˙����#?��>W�l��h����-�?�O��9�?q��>:W?�k�>/}/>9߲�#D]�vJ��#��lU�>�l�?�K2?�K�<qh�=]�j�?򐾘i�>��>$Z�><8=>!q�=�$վ�(U>و�>��E?��?<u�H���\0g�2d�"*�>�l=�����ώ?�
M?ϛ�+�V�NjG���W�X�|>6����#�^���o��"��ؾ󨼾�4>��>��?}�?��ľedӻ�v��2��3�&�)�@�>aZ>l+-?yn��O=f^���-��*����n<��E>H��><���I��>��R?�{Q?�RJ?f??��z>��=�i�=��*�<�.?�� ?X�?�Q�>O�W��ye�������������޽�s��������v�4>R5=m�2<�ѽh-p���<�#�=�<��<�[)=gQ���Ѧ=5��=�	?>F�>��1? �?�v㾡�� z���Q��g>�7'>&:>ǒ�=[ֵ�&1���>��!?6�k?��?8h>��	�J>��>G�Q�<��<?�iQ?��>��!��o�##�����Nr>�&���"�=Ԕ����8���>:���=ft�>�
P>Ƃi> ��?�J?�|*?�UM�}R��0?����.o���;%��>���>b,W>� ��9$��^��d��lP�:H�%���;�=>��>��m>oE>D@�=���=��=���/R�����I��;D��>`խ>�=�>#�=�|,��������%?�Q�<���h�˾�z���n!�`&D��$��$G>�ZþԹ��	ɪ��/��@'?�D�?���?�K-?3���1]L=��j=���<J�>@���=�ї=����>^H%>S������#!����>�d�>ϼU=Ͳ�,��Ͻ��qr��
��Y��K��<!9���k�����-�͞T������e�&�;�y����)���%:
�>������?��V?��>3� <��&��Y �2Ε�ܠ<�b˾:[ �{hʾ޾!��������������=�?� �ʾ��>��]��)��Z�z�[�3�K���t��>�4>?�����#������9/�=��>W�(=?k���!��P���nq�|Dr?�j7?����E����?�*g>�I4?�
?4�4>��a������PC>�>G?�z8?
��=�D�A��&ս��?�	�?4�i?K]־�U���9���Kw??$�?M�+?Q#->=J��^/��P�C?��`?�� ?�V��х�
�?�\Ç>��?M�(��9>��m>���=�㽨ߢ�u���Ug���*�=���=�+��*����$�i�)�>��?�!�>ܭ�6�W��>�=���N���H�p��<B���<1�?j���>שi>��>H�(��������:� �[�L?Xu�?�nS?Y8?^g��C4������=���>�X�>O��=���~�>���>�6�WUr�mP��S?�'�?<��?H�Z?�im�&Hǿ8z���w羖N.���x>U:)>���=R�	�&B�=�c�=��=f���=#�r>tgB>�fp>���=%tB=�Ƽ=��w���R�������������&�$����{���8J��K��;�����ѽ)����0��$Z���]�?#�+9޾Q>} ?��>})�>A�D>̘>��R��H�8u?�E���,~�Q^��t���J٭��p��0�t�o��͍�\C����?X�3���<��> �c<A��=���>�r�=U�>x�F>�B>�R>٭(>5Ň>�->�5>y�=�4�>ەh=�̀�s傿G��VF�S�=�dH?_�"��3[�Jc,���޾�굾?5t>��?��>��!��ē�� o�.e�>�y���ɒ�-z��d;��>I��>uP	>m=j%���$��ٽf�f=�4W>��>�G�m�=�H�=�>�O�M��=jq�>� .?)�m?��?0�=�>��]>�Vn>�T7>|�>�u>�5>�?�;?�=?`ձ>��=L)@��6=Hr}<��^�3..��̍�-�/��J��K��_)�1q�==d�=�i<�r=m=M!�<,���<Ps�>�l�>�6#?Ӈ�>�ﾳ�V��b�A@Ѿ$���D�꫷��}(>�U�>�X�>�5?��?�&>�iJ��ih��6�>�*>�XN����D���x�>3��>�T?�J#?�OM=n�3�%-0�L!3�N�>jf,?Б?�t�=�Y���2>�[��h���>K�e�Ӿ+��>��I>��`�������:m�Y>�Ѽ�	�����#-=���=��=,�=?{�=���<��>��_>*O>Y^=x�>(#�=�6�=��=�c=�q�=���x�<��Z�[�ٽ�-V���K��	=uM�=�==��?���>I�#�6+����4�z^"�^R��7��>�S�>"<�>�7?�+>��[{c�<JI����M[?�{?��?�}���=����Z�;�h�>�Zh>c�>�>=(���߾�O1��s�>ԛ0?/�?�&N��m������
�z'?<��<qn5�=g�?�q=?��!��떾I�"�,�V��Y���@;/kP�z���_���H��%�yR����ƾ�$'��f>U
?���?v���܎�=�_�����s!��֨�_%.<����3�>��<˝�$J@�mI����t��P��f�=OO�>$9!�>?	�+?q�2?��??��>3��>�� ��$?�]�� X�>�J�>xY�>4��>���>yLP>@�=_	��j��di���g����=	���>6� >qB�=|=��Ļ7�F=��>����u3�;��=��X<�=!��=PS>V��=%?|?I�=k���?��<ľc��:�P�=�| ��e��_���;\[>���>�?���>dK�>��A>`VѾ�`ݾ���0�l>�?jAK?�'m>�I��ғ=t!� ��ܺ=���=�
�~l�*��8Y���~�~^9>��>/h�=X�A=�Ġ?�?"?lt?Խ��ʩ�K��\�0�������,.z>�p�>�i�e�.��t$��w}�0qn� hm�e%�N���_"�=�A+>T�O>��<>�^�=���;�Q��S>ǉ^����=�R�;P�>/��>���>IR]>Y�=�a�|%���S?�Ť�K���v
�0;�0_>��>O��>��=�B?��6>d�^������ Z����>���?,[�?$P?+���H�;|=�:A�ҹ!=���>	\�>KF�9<˽�y�=��G�"�T>_���<Z�=�婽K����%�5Ľ���=��a=M㴿Ӳo�=h��9���T���)��wф�a/��u��^��+�X�?�������J���:��Gj��}���o����?� S?)�l>v��Bn�p| ��b���ɽ6SY�R�V��`B���}|�����#hX������վR���,��Ft�>8�o�E��W|�=��\7H�����?�>����U#�~��Z\C�NL�>���>GMW��d���k��C�=
O\?�Z>?Q-�D�PF�����>��?�ƒ>^�e>=i�%=_Ac>mN[?ȕe?A��=L����@���[�:]�?��?�F?Pݸ��o8����$�=��>�>JB?]R>b��� �>��P*?V�V?�@?	�&�H�a�>�ӾL�?v�?���:�>^�>��>��Z�ھ	u�=�������mv�>�͖���>.�D��$̳���f>� >?���P�z��>�n��*M��CE�%,�ˋ�R��<f1�>��K�>��a>�>�x&��׋�N刿����o�K?M��?_�R?!�6?ne����辢���#y=�4�><d�> V�=.��;��>Zs�>U�Bv��-��a?�\�?�t�?��U?�Ll�S�׿0�����j���8�=N{ >0>%��f��,�4���Z=��Խ�=T_X>��:>�*>��>%�>>e��=Be���!��v��oՁ�I/I��������0�:e�D8Ⱦ'4�3Ȫ��L���׽�ݽ,���=i?���O��z���ھ��>�l?w��>��>�E�=�LM>C\^��qʾav�?��8��P��&H��3kž�^�K8��4$��t�ɾ� A�����>K=�j0>R0?�hӻW�O>8(j>�8�<�]�<i�+=��=��>j��=f�">�Y$>��>��->~�>d��=F����m���5�d�%��]=A?n��g��0�4�^վ�梾B4�>,*?��O>�&��3��/#o�7��>i�L��.<����+񮽧��>���>R�=�߬=tE�;K�����ؽ��>�ų>�I>y*���i��x��9
<$_�>]'׾�]�=e�v>oS)?Z	w?�4?I5�=0��>d>�܎>���=�&P>��R>Ԙ�>�?��8?b]1?׾�>47�=��_�C�=٤2=[�=�oa[�1�L׼B"$���<l�)���`=�7u=�l�;iS\=��D=�T��0�;�Z�<��>�2?qG�>_��>.՜�y�T��P�d���o�1�bP����H>3fn>��>)��>f?���>�
>r@�����&�>�D>�v�·x��{u�8�z>�u�>��G?�e:?U��;��6�u~���->3��>~�?X0 ?vI>��>6� =�:��)ؿIZ9�(J���b���ʽ��s�o(��T���I�b5�D�I�����j>�(>J�U>�E>B�>qO>�ײ>
^6>��
>3�=�k�={������&\�<�J���>�ڠ��k��{p��]����������E���9���;�c8?@�>���� ��C�ֽ���Am��?@*�>��?pH7?�~�>����~��S�a��{�0?��g?��?7�����=�,ӽ+����?`N�>
"_�R�������2����/?}�??�>�!K�R:��Q❿��x-?u�:U�?����?�SJ?��)틾'�&���G��$3�rC�=�si��s���缾5L�A����@���yA��+>�C
?���?���x��=A������冿Ɓ������52���>H�5�&|$��}�,�������{����V=]��>�����޸>��7?���>��y?�?�=?y��>�}?J >��1?�� �L=zh=�Uj>� �>(����6�����X���b�����֢�r91>�1>O��=�0 >!��=���=�=�n�=^&=��=�h�=M[�=I�
>$�8>�4>��	?��5?�6�|�}.��#��܁>8�f>���>���=�+����>=�J�=�!�>��?���>�m�<�Z#��,,������>M� ?"�^?�Q�>�T���a)���6�M����=�G�>\����q����.}ھ�J½���>����.;>�L�<�f�?�1J?oL?7�����9����C5���P����>��>.���Tؾ�g���?��k���~�u��򑓾��=�]<>j�L=,b�>I�<�4e�Q�D�ԯڽ�����#>C�"�w:>�F`>�A�>��>G�|�U��;�f��K�6?�-�J<��Ž$S�`܃��tk>�h�;�@g�}P?s����4O�i`�������?��?2��?��3?!�A�3&o=,5�>��$���þo��='s)�W>݄�>M�>)�">1c>�O��1�U�N�+��<>%���y˸�<˾��ݼB���p�t��w=BE���7��u����ھ��<Dt��O��<_��.mU�V{��I��x�)��F���k������q�SX�?��H?�<[>ӏy��w^����������9�c羲�)����p9r�ͻ���뷾�s���������R ������>��??��I�d�F�[��	BG���c>H�վ//��nH�d:���>�?�1�=���Z8���W�=�;�?*�E?�k&�i㾹��=��g>U�'?Ճ�>�+�=�\�<H.-=�2>�n,?8�m?#p�>
��h֘��	�gT�?0(�?̆^?�����O�������u>q�>��½�%>��=�"̾j���C'W?v��?�?$&�6w���`�;w)?�%?�����4>�?���>㫲�"���"�>!����=O��=��ԽSnl;t�O��x	��a�=m�>2V>�(����/�%ѫ>H9���*3�U�@�����B������8��>s����i=Y�>���`�2�~Z���{�럽_�j?≲?��T?�,6?�u�NM	�w�i�s6>�ʆ>P�>Y�
>�Od=a�4>�,�>[��P�^�+��V6*?�:�?�g@�r[?A$^�9yԿ�	�����م���U>9��=I��=2�w���#>����j�� ��.?>���>�>=�>[89>��>�� >�v��
a!�C����$��O6����� �)������c���&*�਍�F�������!��P�\����p׽�D����% =L�>���>U�?�Ze>=v�A������b-<M;ľ�g$�8�2������Ǿ�s��h��`���߾N�$<йʾ���>/bL���=�%�>}VO=�7�>}��>�k�=n��=�O>�s>}�&=�5g>��,>���<�>�>t/>xV�>���=6������LRK��f���=��?�͚�����"1����!���v��>�~"?��>p���ӓ�ok��S�>�+=�|c��ܽꯌ=�W>l�>�%�=	�Ҽ�3=^����~۽�;>:�>�b">=��u�a��븽P��=5��>��վ�]�=P�z>��(?�w?5?�\�=���>�A`>��>�C�=H`I>��N>��>��?<g8?i71?	 �>�=��^�$�=��@=��:��]�aq�����- +�d��<	/���P=�$�=�/	<��Z=D=7=4�ȼ&2t;_�	=p�>��9?�S�>o��>��<�hd<��K���"��� >�;�-��>�#�>��?z��>��>�G>O�/�"¾wIܾ�]�>ʒE>��]��v�_஼M'|>i�j>�P?U`2?t��S_��=�3�=�Ʈ>��?U.'?(^�>�L>������	���ڿ��<����\�
=�p��lj���@u�����[9���1#�E*̽{�=�/>X,>��t>�0�>h>q>q//>h��>��>�>��> �(=��ۺ��	��能Qx��h=��`��aO�jG�n��af�IY��$I=p�ҽ˙����#?��>W�l��h����-�?�O��9�?q��>:W?�k�>/}/>9߲�#D]�vJ��#��lU�>�l�?�K2?�K�<qh�=]�j�?򐾘i�>��>$Z�><8=>!q�=�$վ�(U>و�>��E?��?<u�H���\0g�2d�"*�>�l=�����ώ?�
M?ϛ�+�V�NjG���W�X�|>6����#�^���o��"��ؾ󨼾�4>��>��?}�?��ľedӻ�v��2��3�&�)�@�>aZ>l+-?yn��O=f^���-��*����n<��E>H��><���I��>��R?�{Q?�RJ?f??��z>��=�i�=��*�<�.?�� ?X�?�Q�>O�W��ye�������������޽�s��������v�4>R5=m�2<�ѽh-p���<�#�=�<��<�[)=gQ���Ѧ=5��=�	?>F�>��1? �?�v㾡�� z���Q��g>�7'>&:>ǒ�=[ֵ�&1���>��!?6�k?��?8h>��	�J>��>G�Q�<��<?�iQ?��>��!��o�##�����Nr>�&���"�=Ԕ����8���>:���=ft�>�
P>Ƃi> ��?�J?�|*?�UM�}R��0?����.o���;%��>���>b,W>� ��9$��^��d��lP�:H�%���;�=>��>��m>oE>D@�=���=��=���/R�����I��;D��>`խ>�=�>#�=�|,��������%?�Q�<���h�˾�z���n!�`&D��$��$G>�ZþԹ��	ɪ��/��@'?�D�?���?�K-?3���1]L=��j=���<J�>@���=�ї=����>^H%>S������#!����>�d�>ϼU=Ͳ�,��Ͻ��qr��
��Y��K��<!9���k�����-�͞T������e�&�;�y����)���%:
�>������?��V?��>3� <��&��Y �2Ε�ܠ<�b˾:[ �{hʾ޾!��������������=�?� �ʾ��>��]��)��Z�z�[�3�K���t��>�4>?�����#������9/�=��>W�(=?k���!��P���nq�|Dr?�j7?����E����?�*g>�I4?�
?4�4>��a������PC>�>G?�z8?
��=�D�A��&ս��?�	�?4�i?K]־�U���9���Kw??$�?M�+?Q#->=J��^/��P�C?��`?�� ?�V��х�
�?�\Ç>��?M�(��9>��m>���=�㽨ߢ�u���Ug���*�=���=�+��*����$�i�)�>��?�!�>ܭ�6�W��C�>d���EK���H�R/��#�DQ6<�3�>s��X�>fQ_>��>(�d~���N����68K?�W�?=�R?��;?���#�Lu��5:}=�<�>�R�>�ݣ=��
�&`�>��>~�쾨rp�O����?r�?J.�?��Z?i�i��Qտ�[���F��G����">&,�=п'>T]㽷z�<_�!�j��,�]��=[Uy>�)H>��P>�r&>��	>L
>ve��.@�%���ǈ�[�4�xR�
q�D������S�$��teɾ�������H ��{ڽ0uj�wf�����Sa)�_ݚ>�	G?��?P��>�L�=�t=i;���&�a��p��6����꾗վio��K���4K��d��l����<KF�����>�뼴�p>l]�>�m�<iԏ=�I>��U=���=�Ի>4�=Ŭ>rn�=K�*>I�>sݚ>p�>=��>Iwh=Q���|��<Y@��>���<iD?�1��p����4�R[�"����^�>�3?�r>��%�>��Kq�"��>9�X� ������A�1��&�>�>o�=9�<ZB�t�R����=p�=@�i>�)�=<�|�_���0����=v��>Db��~�H=�$�>�C2?Ρb?�R?�B�=�,�>��>�y�>��>�9�>ٹ*>�,T>t�?�>?�P/?x�>��=��J�$L:=��<ۃT�9A����;}n����s�l6���,Ž�-=!É=,rF=A�S=e�?<�{��ʶ<�91< ?[�>E�>%$�>�D;�	�B!$�+���o�;���=��S���>X|�>[ ?i�9?���>���<>�	Yo�y��>�Q>�t�����=��
�>o� ?�^z?Y�R??U=5۾���Y�W�ؽ�Z�> ?i�?.>@"�<�r(=R���a��������j��=0���pg�1��	�����������O/P��C�=Y>3�=��!��=e�I=���>�<�XNh�$���\<�呼X��p2���'�=ϴ=��Z�{-=7ɘ��p��ӽw@:��"h�*��e�=��)?�h�>����ݫ�9��ޯ#�z�'�.�?V0�>���>(?�߅=L
��Jt�
�R��7K�Ɣ�>��?*(?0%�0R>�ͼ�(=���>���=GS���M�<�D�X�Y�z<��#�>/�*?ȶ�>�,ǋ��T��$'�2��>���<M0��0�?P�D?�2�8���В#���J��U�K��<$$��፾�籾(��C`1�ٞ����rO�9@>��?MA�?,���a�=����V���d-���Z���?�<��L���>��=�<��lY�nξ�	s� !��r�=aH�>.�.v�>�L?�U?Dv?��_?=��>�MD=���>q�~>+�?`ma>���=ږ�=�>1E>��Z>���o�߽�a��:��"sؽ{BY�(�j=�>>�0q>�t�=\�H>b� =z��잽��=���fG�<'�=g�=�^>�f�=L
?2�?���V���ۣ�rY����=�=�}���qؽ���>v�=6',>��>R"?�^�>��w==_�����c�͝>[�?�gD?<��>i �����A 7��Ӳ����=�&>�4�=��ɬɾ���w�K=��=�Q
=8f[>4z�=���?G�?k?���!G��3�G�,�)/=}8�=�T? ����<�Pe�@���QX���e���t��஽l䦾8|�=�=�>�>�B�>X�6>�Žg*O�>;��!.��;�=�[ؽki�>k܉>��>,M>֞�=�B�Kdھ�oK?x����\)���+��%�Y�g=P6�>m^E>��=Q4?�b@��l�^˔�_��!?���?餰?�y]?~,>*Z�=+�>q֢��������>�kŻS�Ƚ,��=sjb�����>55��［@��𸐽��F�UAؽ���CW�=�[���V����;%���:�y��qq���$�}W���N�5�ؾ����)r���<���V�g]3������ľj�v��T�?I�A?.#e>��m�D��&���i�}���D�s��`پ���Q����o��1ۖ���K�Nx۾V��������>=hr����;�e��]���5 ��ǚ>���Q&��6���.� :�>Nf?N[?�@�]�����dP>�Vc?hp??vtH��D�b�0;<�J>�:?j!>�=�<"!��内=�j>rgu?���?7�>�2���6��ox<���??�i?lV?���G	K�5v ��ȯ=�~/>���=��>�&>��A��z���:I?�*k?�w�>�H0�"�X���5 �>��>�W�Xі>��?���>�־P�����>����e�4��=N)��]c=��Y����,�>��A>+�*>HоZ���*=�>0a쾘�?���C�� �t7������>o�����=mH>}��=�.�;X��.7����սF=R?�`�?NlK?x�<?�ľ��߾m����=׳}>?ԑ>�e�=��P���>��>���4�{�8��h4?�?We�?�(U?	�a�0�ۿ眿1촾���*�=S�b=1�>je�=-!=��v=��M=R.�=�Nm>A�>�K">ɦA>�h:>9�A>#!>^����'�5L��{P���~A�v����-C�S��N���-��I��q����͈���z�m#��by��Ȭ�5炾��>��>?^�>�6�>�hX>��>�N�������i?�"�z��	���Ͼ����Y־.j����r�/����H������+� `�>O�=�!�<���>$�d=$�y>�$�>L��=�> F>��L>[��>��<>.SV>	iK>���>�L>�+�>C��>%���P^���,��e �ƀ=)\&?�s�=�|��/�8?��U>�}
�>��>&�=��1��0��]�}�M,�>Y߼�e��f�ܺ�=n|]>$��>1�=������E�Z����y;��+�=20�>���>q3�=�(^�aMJ��b���2�>J���۸�=7z�>�QY?���?ͅB?�ʼ��>��N>���>�>�=���>�9
>+t�>)�?�&*?aG5?�}?���=�4��>�#�<��G�B�K�90��^E���{(�v!+��3��Q�=��[=�ϻ��L>�j>^t>�$>���=��?.H?k�h>͍_>����HE2���E���'��j�>/�=��>3:�>Pg?���>>�z>���=�U%�l��O���h�>��P>(�f��	~�Z�<B��>��>rlS?:?�H��J3��1�=�
�>ϫ?@d?��#?�D�>��J��K�������ѿ��6�m��P�ü���= Q>��>E�==6O�=!�=7z4=b��>D�v>&�j>��,>/�>X��=�a>A0�>���=�]�<3�>�*5���>R����=G��=kf��AJ<.X����%�+ٕ;��B��X����鼔2��U�>�
?z!9?�+�L���������W��m+> ??� m>E��;;�9��%���d�Gq��5�>9z?�S�>d���c>_�ľVⒾ5��=�>�QZ>�2񽊈g>�I&>7��>L3U?��i?u�>n������ w��^X�W��>�<�Z���?�N?��3�<hJ��3)�y�4�̰�g$R����,��{˾w!�W�-���پv���Y����x=W5?�U�?a"�g�������KM��m8���8��J0P�O��;߳,>I�m��Ǿ_찾z���O�x���r=]s�>'�>׫���>��M?{MP?w<!?̟>?dW@�&�>k�>��	?Շ�>�b?�Rn>��=?�ؽ�HսfY4>v�o>�ݼ�����û�+��>� >���>>-�=]=���n5���ɽK�[�+U<%(�=�l�=g�>>"I�=��	?q�F?�"��羱eX�<*���[�7�>{V�=F���`�ؾ1R
�WE��*?�C?��>e^V��w��M�ɾ��:�N ?H�o?��6>�Oｸt�.ֵ��q����@�>� >�4���
,�_��!���m?>\�>:A̼�9�>��m?u�\?�/"?*t�>�1�ޠ_��a{����{��}�?��?���=���Xt5�0�|��}�rhn�J^���2D��sc���{=��e>V�o>���>�$>e��2!���Q�='艼{���;�>�r>x}�>�c>Z8�=ux��QU�[c?�P��SB�V����o��4�d˼>|�Ⱦc�U�ȭ=�{���W�
T�RA,?���?_��?9?u�=F���>Gj�=��c�yʼ>;���8��<g�O��|:>�Y�=ݰ]�V�V���;O�9>ߊE>x���}����:i��Y=�����2y���ɽ?�p���������;>�u�;ta�!C��e�2��T���*��wͽ���(� ��]��.ʘ?_dS?���>K�i��6|�����������F��*YC�����5���x�-�ؾ�ľ�I˾�b���r��_ƛ>�YY�KC����|�f�(�+ꏼ�q?>�./?�@ƾ�������(h=Jq%>���<�L�R��������7�ZW?��9?H쾙+��DG�u�>��?F��>��%>@+��HG�"�>�:4?G�-?2����-5���=��za�?���? �@?����-R�����#�?�?j�>�<�5C��+
��?��>?�>�H��R��� �s��>}!??j�I���T>p�>��>�ཽ3���� d���D�ko�=��� )/�-|�" �,�
>n��>b�s>��T�"Ӿ"��>�^���N���H������p+�<Č?���x�>�i>��>�(�����ǉ�e �u�L?ז�?ÀS?p8?;-����c����M�=Ǧ>f��>�i�=GK�cĞ>F��>d��ьr�!���?�G�?���?#SZ?�m�Eٿpz��fɾ�ؐ���>,c=9>U�o�ͧ=?n%��=��=��+>m�>��H>Zw>�O>�z+>QN>>B�����7:��P^��W�E�����-����5�������땾Wꬾ,ѽ~~Ž��� �1�DZ��&�!����>�!?{[�>�m�>�7B>c:> ����U���p�9��0����}�dԾ�&���>�[�t�b��?Τ��\��$��>)21<t*�=�6�>�ȻR�>�>d=vm">��=>)u>�f>�6>MeK>;�>��G>��>1�>8�>�/��:����&��ғ�[8��^5?Q|t��텾x�+���ľL�B��O�>�y�>���<�5��������D��>�ݼٔ��
� ���$=l.�>m��>eǽ������ >[�:��Y%�[p	=B�>cT�>��=�\�G ڽ�ڽ�M�>l�ؾ�v�=h~�>�0?��r?YX8?��=�ǹ>���>��>6>��R>�r>��>�k?08'?��2?�$?Gb�=A�N�E<�o=L"<�t����ֽ`<3���'���KN��ވ=��Q=�P�<V7�=�M= �d<b��<�c�<r��>k�B?N�>�|�>]$f�o�H��	7��� �O�X>�M����>@8�>�?�&�>�Fy>��G��>-�XG��8ھ���>�_�>��l�P����e=^J:>�[>ʰ0?V�=?���<j(���wZ��c�=Ѭ?��#?�:&?��>��=�M����ο�d�%(�|��ݼ�?=>e�X�ýSIO���潏�o� t=�r>�W>���>�
)>�>�`5>���>B�>.t�=�Ӽ=b�r���=������=�E�<:M9;#;���s��"<�x����9���\�����3Ğ<3�r����>}D?|�=Gt���U�iL��ؾ���>�.?t�?dd>h�$�kV��4��b�p�.�_��?�jl?��>��A��rU�^a５�+>�q>�_�>�<�>�+�+�_�`ȳ�&q�>|�?ԈY?�x�>Ң��]���7���I�)��>,*o��s���ϥ?�U?'�A��潺*#�v���8�
J���q��þ�D׾_��c�q�Ѿ��þ�%�Fs}=ʠ?D:�?'g����FӾ֘���o������6�<�����M�>|�A������r5���a��1��G��hi>�z>�*޽��>m�Q? �x?n�2?4H:?
�o�Jː>��>X?ϟ?o]?0?�p?�) >��4�	 �=E4�>�@4���E��������RG�=�D>�T>��>���=zAŽZ�Z�@��<�hN=z��=/}I=Mz-=�&�=��X>t1>C#?�5?O׾@I����:�3z��-#>ƫT����=M��>a<z;�<>�H�>Z!?d� ?�74>[�"���s�+�K�վ�����?	[[?9`�>���=�7>�y���L��0��= �>���=�(�����TF��A�=��m>�|�>w�~>��G>N_p?�*,?�j?�=�10 �e�K�B��]P��{�B��>G[�>w0>�sپ��V��́�^b�WH��n5�4��d)�=!�<7_�=�F�=���A�=�<J<΅/�����xG=:�=°�>���>s��>_ >- ���۾� �?}軚^(������ʾ�f���澩��>i�h�Wߑ=^�.�Y؜�㽿�	f�l%�>���?�.�?U�Y?Y������(]�>�U�F����>4�G��T�=l&��e��>��>������Jb= F
�ՠ��r�ɽg�����?�3P�,�ȿw�~�C�<E��"���S-����R��=ē�s�?�{�}��K�y�������{�����\m�&�R�=v���?a�<?���>���=�Y��ڗ���%se>E��ך����վH���ľCʾ9��� ﾫ�뾊
 �����bC�>��W�V����|���(�Ò���?>�j.?%�ž�����)��]k=Y&>g�<w��b���w���D� �V?`�9?ne쾠���Xݽ��>�?}��>)(>x���=?�3�>N4?{l-?� ������n�������X�?��?�@?����D�͜����4��>��?�e�>䄾�W��v����??9?�<�>0���Ɂ���K�>qgQ?��X��.>�$�>�s�>2�ɽ�8���\�xA�WG>�[�>�<�ǽ@}_�5e���=���>��k>�SY��r����>{�R�پ��A��~��4����[����>�н���>	�f�H�_��Li�i��h��L`���<?aʹ?L�Y?�?"?���Ⱦ�)Ƚ)>S]�> ��>:��Sx�=7?">��>ex ��~m��u���R?
��?�w�?LM�?k��d ��$7����ھ���FC�=�>��d>�<��=R�f>�=T�<>��>��>i��>'l>4W�>��(>U��<X^��9�#��ٙ��W��`�L �����V�L=�ı�nսC޾�a=����Ɋ����Ž~zu��\���B�����_ݨ��d�=@D?
�>9�>0�C>w9>��}��
�������t�Ps���Ϟ¾�Z`�[2���S�����,É����'?.I�V=�=6s�>�Fb����=hZ�>=�x;>�t>6�>@>Z;>��P>�q>�"Y>�o�=���>�D�>�����$����(�^�A�����+?�������'d�[���
�:/�>��%?[>��d�����	���2�>�cüع��UP���=�>��>F�<S���j�=�P�5>\���><��>��>�U>�������5���%��>p�վx8�=���>�L3?*�}?<�L?f�>Xu�>7��>QT�>�>d��>ֳi>ڙ>��?�X*?P�? 
�>���=w��H�㼲��=15ɽ�)+�Zzb��H��Q�h<�*>x5r<+>��)<8�=O��=G�=�fM<r��$m�=��?��E?P�>�p�>ޞX���<�#�N��~��<4>$�+���>1B�>�4?�a�>n�>R�i�]�F�RF��wg�����>/�t>��q��v��!�����>��Q>��W?��"?�꽺�ھ{Q仝�>?s?��N?9�6?�=>}=׿�0���ҿxk��J��C��=�y
>@&�>�i+>C�">�Zo���=u��=�ss>�K>��>0��>O/>�"�=����خ�>SM>~h�=T��c�>T��<���=*ӕ��!����F����	��fi�<�#�<~�;%�<X$����2r�=���>�?Q��=����d��'m�\�����>��
?_��>��>�s���,�˨e��J�w��z�>��k?��>'�$�/���=X{��ʊ>���>�	?40!>r���܊���¾�ɡ>��>��U?��>��@�(/w�q��� 7N����>�%�����<Y#�?n ?R�Z�����7���4�1�؂p=��(=Ci���
���D���f���W�ț����0�F��>���>�.�?ʆ½�=���=&���#d�V�Z��y�>Ӏ�>PEx>�l>� �����lB�Q�۾�sm�>A�=�u>�ߣ>�k�<��>*�E?m�b?�CN?�;P?��K=�>�a>�9?M?^�?�[?{�?}ԟ>�B>	�>�a:>>cӻ�`e�)k��jѽ���S�>��d>�Y�> 
}=��>���=�m7��́���\�=��<22�=9jw>�i�>�5"?N�D?��ʾ����fm>�`��֥�p����I��} ��T��Y�i=���>��,?�!?-p�>�=^�r�E�Q�J��-ݾLĎ��S?��~?�Z�>�Q�<n�N>V������7�š>>8�[� ���վ�bʽ���>%��> )3>�k>�Fl?XG7?e�?�k�:�!�D2j���#���Yw*�#��>��N>��|�(���e�L��k�_��{(��=�㡽;3">Y���Э@��V>�;s<�[%>�T5�����V�!�5WB=�> /�>���>��>��='��;s���V��q�6?ck�M��ێ˾ ���k?�����6'>� >ZO?�7��3���Q���?a��fJ>+��?��?��?�)n��h�@�*>Ȣ={�&>:q��;yp�A��=u�=��=��(<�y�z9����=�C�>,	�>������������dp��$&K�ϛu�t��Z�¾NC��I��k>-��'��
�I��ƅ���2��E��*Q�)�j=t�5�}���������Jt�?�=�?XJf>܎���u�^#�%O���<pþ���﩯��ɭ�H�ϾAdᾴ�侗-+�E���A�������>/�Y�JA����|��(�
����~?>�4/?�`ƾ�δ�{���g=�b%>ɱ<�9ﾲ���篚����aW?o�9?�O��)��3�$�>��?�q�>D�%>�(��B/��'�>.84?��-?�_�����9�������l�?�?��??�O��A���T��3?ũ?|��>�Ǌ�^�̾zN�"?�9?�ļ>��f��c=�u��>H�[?�GN��ib>���>�A�>��b����F&��@��������9>#�����Rh�)>��ڧ=�>�x>�$]������>�B�k�N���H�H�����U[�<ڇ?U��a6>�i>bB>�(����ω�f&���L?���?��S?�k8?�^��*��l������=^��>Ѭ>Y��=���b��>y��>�d��wr���d�?J�?���?(ZZ?ۙm��~ԿxV��YӾEo��`��=E�=<Ņ>߱�=��>��M>&K�<� >��>|	�>!�v>�cX>_u$>�Yz>?H >������(�K替?ג�Z�I�E��ʓ��r=�ƾ�P��������xv�`�)�#����<`�ٽvȽ��j=>+q��(>��?�~�>t��>�^R>�>����Qm�mb�}�@����=��^� �s[۾S.���)����9�(ⰾ�����R�c�?t+�=P��<��?���=��P>^y�>0�I;:�=m%�=5�g=�>>�#>w�?>�.> �>��=o�>��\>�Z����������쾷�e����>�����a�P�s�#�
����?��4?��>n������r�*�O�>L^4;��Y���9�⢩>��R>�3����=���W�o�}E��:�>7e�>�J>���:8Ar�ԗ��j9&�4s�>�~Ծ�I�=�b�>*�*?trq?�[9?��>+�>�Ѐ>�ܚ>��>~2W>��,>��{>{b
?��6?��-?���>���=)4j���$=X^5='O�VVȼ$̽����lC������L�y�w=D��=J�I<s�i=�2�=^Uڻ ⚺d�N<ʵ?��-?k��>�X�=�i$���z�7ll�6Z�(TA�q�����=u��=���>�8?�*?���>+�o�ж���q�'��>|�y>ؚj��Ꮏ�?	>w>��>�!?]?V�`=�G�������=G#�>�Z?o�+?�Ez>���<���<�������Cx�6���L��H>�~�>gɡ>h����>c9�<Ѱ=��>���<0�>��B>���>Y�>�3�>�k�>e?n>��<
��<��L;A[=W�9��MW�ċս�⼍���F�ƽ݁c�����C�*iI=�]�;�Gͼj�e��p#?��3?�)�U�g��j��������>���>e�
?;�>��7��'��k\��fw�#�ھU߫>D4�?N�?k~��`?>�#��3j�E��=�[�>���>2�<'�Ҿ�‾2

?��)?%,Y?�e?�Ƅ��̎�����#E�eP?1e�=�nu���?��I?��j������:��6�k���R	�B������i����N���
о�������=��?f��?�1��u� �ԏ���ſq��S��� ��3�w��X�=ˌp��͛���w�,ʙ��'=���ν�~�� ��>9��>?k�=Ƨ?�*a?�ln?��$?%4?�2>X��>��>�_!?�?�a�>Ų�=3���x7����=l"�=��,=�s_�(�A�V����D��V�=-4�=�h>�V�=W��=~a >��R=Uv�=.�>��S=�˖=d��=#K >�}�=��->E8?]}>?/;��&��D����2䤾���盽^�����Ծ)�����=�0?�hD?�Y?�J��u���ؾ j۾�g�=o�?`�h?ܔ>�L�=٦�<1�վ��:���=3�B>J��=H��:89�i��N{��>���>�y3�W��>���?��!?*}�>E񯽝�!��L��I���սp�:����> ��>)�^>�ɾ�<�=�o�������y����R�Y�y�,��V�>���>M?y>�p>��g>��:�����,��l�)<�;x��x�=�/i>L�>��?>�2=Zl��劻��F?������¾)������Ǿ����b�+��&u=��=�P(����!¿o<K��u�>k�?���?�4W?�ܾ>7A�3F�>��=���=aa�>�����b=�,�a��>H��>��o�'����Q���h��쓾g槾�����-�x��Ϭ���i��,��9��G�������Ϝ���N�h�� ���Ჾm��mL��`�M�-d8��@u��*?����Bx���H�?+P?��>|J�=��BZž�t4��/½I���X�����mF��ړb�GZ��]Z~���o%�{�;[��Xϛ>}dY�7��X}���(�t_���?>�/?Ɖƾ������e=�%%>�Z�<���T���9�����6oW?��9?o?�'?��Z����>!�?�R�>��%><�����"�>�74?�-?@��}���6���<���h�?���?XE?��G)I��v�;xL�D��>r��>�-�>�4��3���Zn��M�?U�3?��>E�����_/5��O�>K�@?�TU���>��>{��>�>������ּ�}6��Nʻ���=���Li��- ��-��cU>�Z�>Y�}>�?��� �F��>���ۑM�yBH�)����B�o<��?���:�>h>g>��(�\�������[��M?�{�?�S?��8?�t��y�쾅���9C�=@�>��>��=���0ǜ>e��>��p�r��K�C?3@�?���?l6Z?�um� �ӿ������F����V>�+0>ʼ�>���=23�>?c�=�DG=@�=�>��>rV>>�of>\=�>�^^>
W}>5c����#�N�������w�-��K�(�ھ�J����á�#HӾ[y��at��Jtk�xy��.�8+���!�}w��yFI�j>�"?<�>���>2�a>��	>;'���+���H�}�5�H����̾-�	��߾�؛�e8���,�i;�ɤ�M����>c�m<��F=I�? �=7+�>:ԟ>���;|�n>4�->?�=�Z�=D�>�xw>m�a>�T�>|��=w�>�Vv>ڶu��#���G&�{]��m;c����>��S�l\�]�����Y	�> �@?���>�^��eM��4�$���>[>�=𪴾<7^��@=�x�>H�>�սfre=��x>�뛽k�y��Oi����>�CP>%f=-�s�37F�C�<JR�>l�׾Y�?=�>Cd-?k~f?ɟI?��1>���>�V�>ꀯ>G�1>Urf>\Q>�9e>"��>��&?\�/?f.�>$�=Z�M��%{<\R�<�|I��F���A���S�<��<�a�=UCɼс[=�5�=��G=B�=��-=��%��@<�ʪ=��>aQ9?�9�>H��>�V��TP��T����e��=�8�[r�>Bj�>e��>��?���>�"x>~�+�<F޾oQ���>�j>wro�ʁ�^;R=T�c>�Mw>Kg8?k�*?��5��.a�j��<(d�=���>}?�@+?_��>q�=1�@�����vᲿxq#��!�{�=4x�>WC�>�fv>V��>��> �i/k=V�=�S�>0�>>
��=|>^jP>�}=�<�><Ug>O�=
�1=b'���=����\��J�ļ�oU=��/�Lh��ؖ!�����p�輄�8�4���](�g���Y�?_�D?M�1�N���~����Ty���=&Q�>���>z'�>�A������B���j����Aj�>x��?u� ?�/ͽ��=+ɵ��U��t�+>��e>�>G�2�V�J���n�Vʴ>YF]?��e?�F�>7fپ]6��N�����
����>��=�K�<:�?I?n2W�Kӽv�:�	���)��̼�н׏��������ph ����,ڢ��}��;aW=ѯ?S�?.K�`J&;M�ھ����n����$��C���P$�}�'>N��{���?þ�1���:I�,�w�7��=��C>�ǩ>�ϼ0��>��d?2V?�?��F?2�=N�3>���>�%?y?�C?v�>O.�=�,��Lџ=Ĳ�>!�>�f��v ���.������=3к=(zb>.U�=)Q�=�*=�Sx�_,I=Q�=V�>pi�=C��=�RB>�c)=WyU>Ix?�D?-��f���@��5�� J�i�c�����0�����J��N�D�?�A?Q?�}]�Q�H�V_��Ͼ�f:=��2?EAU?��>=��=S�>�ž�<��O�G>y��>@�Z���Ǿ�-��İ�J��zG�>[Ȇ>�����۵>h�v?-�/?��>�Bi��N��E]�ĄR���!�� �7��>Db�>i��>O���0K���k�J0���M��)��(��/�W�H>��>�>�M>�>��=���Y���jH<՜����5>=��>��>��V>�&=Xl�و�
�0?�!�=��s�D� �-t6�x2�)��]���f���Z� �q�3�bQ���.#�R�!?z��?���?� ?�ӽ�얽��>\"νL@�=-��>���o7�`�ӽ ��>�ģ��=ؾk�5���>���9u���7i�t/0�J$;�έ��Um���iZ��:ؾO
��I5���?0>�Ǹ�U]�����)�)��l=��*2;\ǽ�6���4�����y����?��I?	�>U˜=1U���,¾�&`���.>eƘ��v����<�¾�K���S{�����lp徚M־1T��'���>чY��@����|�F�(����/�?>%5/?�]ƾ�ʹ�s����g=�a%>ꗱ<�<�U���������7cW?��9?�Q�>)���� �>��?xq�>c�%>'���B��%�>L94?E�-?q$켎���9��r����k�?M �?m@?���'K�`b�H�*����>��>0��>�-i���ξ���E?�B?ـ�>s�������y+���>q�B?�S?���G>k��>>��>�����r��v������+N��V)>�8��!��K__��y½��!>��>��l>~	��%���1�>jҾv�H��1G�J���:U�J��<��?��侺�>��p>е >�5��C��끿����"f?9�?	�L?�4?������sP��6�=�f�>�Ҙ>.�$>�t����>rG�>��뾚zs��_��>L�?	�?A�_?O�c�g��� 5��P$о�rI���>dӄ>��>r@�!lZ=E��=�0�=�>x��>D;�>^P�>e(K>\�3>_�D=���=�q����&�����q��SC���1��$�\۽�#���m�&���վt(����ɽH���*�ٽ䌾mi;��Ry�.C���ݣ=!s�>
��>a�>g�Q>��]>�ZN��Ӿ�dL�Wܚ�'���h �a�Eɾ��f��'P�O���H���-������?s�<*�=��>Ng���=U^�>v��<��>�#i>9��=��B>�>�&>4�:>��h>OQ>�5�>�u�=�����ҁ�=�8��O��g%<#B?��N��4����3���۾�5���M�>�?&J>"-'�ﳔ��uw����>EX;��X�������ݣ�>Qr�>�ʹ=�>��ę�NKz�����7��=Gk�>4�>4|X��ҋ��E#�Gw=A`�>������v=��>��?#W|?��6?�4'>�h�>�q�> *�>��<�|�>z�{=��=m�	?�%2?�?!| ?H�=�GE�4��<D��=�w��$ =Rΐ��ͥ��Z�/U���*�=��J=�"�^>�<5>���f<��*=d�6>�^�>���>�[�>��M>���=��L���{���\6��W�;	)��-??(? k\?��>~1{��'�n�ȼ���R�>�">�]��9Y��Yн��=�~�>:U?�V8?��<>��<�����="L3=���>���>b��>��>#��7���Ͽ_9��.�e��=K�m=3c�=���=g����AI��8�Z�ľ7�F���=M�>���=�5N��[��w=����>ao>��^=��
>�;>���=v�x=��B<Ԣ�=Z�=BQ��{ݼ�����A��Y�����L����Uǽ�$�=l�$?�~2?���VGܾ�"��]M���p�����>�l*?�5?"o�>��$>�(���^���T�^�i��>dx?��?H���:>�@���>7��>�a>�@D���=�S����>�*:?^�>�y7�Z�k�����R����>b�ŽG�쳨?��g?j^��ʚ���3���H�]��nI�z����TA����b��6�˾��E�Q\���b��@p>=?�R�?�G��M���w�'��ul���,��@TK�Aּ>ʟ>�lu>�c����>i��� ����V�b�ף�>�>�a�>Y�>���>�?�dc?}�?���4�>�M�>M�R?+�>1�?M>*�d>�`�>*�]>�s~����>�^��;.������l=�'>��>�#X>6AY=��Cz�*=�����J =���<��4�=l�gS�=[�!>3��>� ?�KE?^��<��C��F��"?��.D_>�Y*>)�>��/>�Iv� ��.j�=�o�>� ?�.?y�<>R�����J���Gm>V�=?�G?d8q>�q���->��¾7��KJ+>��>z��'w��FϾ*�i�D��;�<�>S�>2�!�l>�~?T�>?�*?����-�xat�ä*��I�N��]O�>�ޤ>�d�=G�׾�7���s���_�c�2�XZ���F��s�<���=:�%>�C>[�==>a�=����#ٽ;��;��ȼ�b�>5�>c�?��e>�u�=�����w�[YI?Dn�v�������ھ�I��>��>4$Z��)?�4�fs��v���<��q�>��?N�?8sv?Բ8���̽�؇>��;>&�8�A��:[p���%����>-6�>�>:�W��v�߼V��=s>lͼ#�ž�����A��*�ƿ�z���s�r 9�,#k��0}��f�3j&<�v�a�S�?��n���s���è.���)���f�˾h辵X����}?��H?�1�>���>e+��V#��U����p<����������tF��㲬��թ�h���Ǿ�a�͗�}
�q��>\���$)n�3��:����%	=��	?�辒�Ҿ#�#�b��=��0>�>hp���T������W��dQ?��9?���}	����-�
U>��>���>�+�=���� ����>��B?��D?�5<=6 ��F���f��D�?Z��?;�>?'	����>���/�֗;���>���>\�>o<�������L�`�#?��=?/�>�B��l���| �'�>�� ?VB�/E]>���>��>U����RS���=}	X����*�=}�ŋ�"���օ��p=>�b�> �>f��H��ƥ�>���`�K���D����%�N�`<PA?���Q��=De>-
>�*�+��
]��m� �kM?�A�?Z�Q?��8?7��B�Oï��w�=,�>
]�>���=[x
��ޜ>3�>$��p��p�#�?���?���?�4[?j�l��ο�ࡿ���Q,��}�D>�&�>o_8>�e�]>��s=ܡ�=��n=�0> �>�X�>�>�M>xom>��>%��o�)�V#���`���'7�v&�����᧾J(�gx��ie)��
ھW��y��f;�+ҟ<�R��H�8n=꾬ʼ7!?#~?�?Q�>�e�>a<`�W䍾��������N�LX��Q�����὾�U���&�e)��ٍ=l�����?S\�>6�=��w>�=�8���:�Ԁ>��#=���<]�>����H=l��9=���=�Zk>l�K>vBw>E�=�	��1y����8�qVH���;B�A?�	`��O����2��ݾy���Lރ>�R?�K>�Q(�H
���y��Z�>st.�yNS���¹����>���>_1�=�����:w�����F�=L̃>��>�?��9}�������=� �>vz;���=l1y>�j(?c�o?.�4?2ʑ=!�>аY>t�>/��=n�>>�GN>,�>�?�Q;?�t2?���>���=�b�
��<O�=��>�e�d�D�����E����<��ӼȈf=�]=�F<�a=Ù4==��Q��;���<�/�>��,?1j?�l�>�T,>E�	��̓�y#�?��K8������q�>�� ?}�j?�AP?�T�>#����ƽ8�=�>0i�=)q��@1����:Q]>\�>@?_�?D�<X9'��W�=`;>s�]>u�
?�I?�B�>��>��ǻ�j��}�ֿ�e{�}{T�t->c�g>���=X��)_��yp��7���s����=�F�>8]�>�)V>;Ĥ>����>�M�>��a>߰=�T= �=8>���z��$�=/�pE<�9�������;�<�=<��xӊ��/K���}�d�*?+s?M78���`�+��xb ���]�ˇ�>�'?�D?�!?Œ>�~Ͼ�T�a4L�IzY�6�>�[\?��?[��Ł�=A|G�t>?�q>���>��d�����y��c���#��Kz?�
G?P��>�%����y� ꂿr�E�ß
?b��3vi��ئ?���?8��Y������6����V�V���\��ǆ���(�m�2���/�~)��q�sX��J6����?W�?�d-��qk=���`���.ᑿ��
�jG��8��d�>}~�=���~�i�#�Ѿ�E��\J>��>F��>1$�=(�>8n???J_?�1?_?ak���?^�=��>sn�>u�?|�?��>�#�>M�>t|a=a�X�*���9��_��;=���=�%>Zn&>Cd<��Q=?m=�g=j~�C#���<��<3��<���=��=�}>o�?c& ?�B#�=�x�=��c�L5���,���!D�z�;�����ս��=�?��F?�&?)VU>�����-��~�ƾ�e�=��>��?���>�U׽�}K>)Ҿ�nu�	��=2��>�u ��G���-޾^����<�dM�>�>q+���>g�?my3?
?����{���a������>�>��!?{Qv>dv�>�A�}�;���|�(�^���_b�=��C��!:�p�>*NR>q�>h~���:��=���=9�3��B
<~�B=�n>'$�>m�?��>6�=T��WҾ��=?����T�����D�^���_�5�5=���>MB��O�>j=��k�V��a��-I�k��>S5�?���?l/?�����A-=Yp><,�=&��9;��	�=|n�Nf��-��>�?�?ֽ��{=��=L��>)�L>��ּK����#���'��1M���X�W��ڱ�9F��(U����ղ���wS�+�꽙仾q���I�=��T��5��1�U���} �����Ǌ?�
�?:X�>G��=İ�󋪾j�o�A��=����3��";����皾�о�ǵ�� �~N<�׭,�q~����>֨T��s��;�{���%�Ey�lK1>d+?MUɾ�	�������q=�n'>�L=$�O����e���}X?W9?o��?����׽�H>��?���>R�>:������!��>e4?`"/?o��������p������!��?�?'�L?��="���E������>ޝ?�?���� >�dn>	eO?��Q?��==�M��k�ʙ+�ԇj>�$?�U��u>�H�>
�Y>�@� ��=��,>�����!=D1=�*�>q���˻���%����=��>��>����ң�
��>#꾇�N���H�7���d�WR�<a�?ۏ���>o�h>o>�(����U��������L?��?�lS?t[8?��������3܏=�Ԧ>��>Eɰ=,L���>Z�>�u辛}r�.'�Ɗ?�D�?7��?�YZ?)�m�Cۿ�ƨ�8i��6����>"">��L>9fƽ��=�T>d2=>�P�s�">Nd�>h�d>q|>(2x>ЦJ>�Z�>�ʅ�@b�����L��1�I�s:$�����s�Q��n ���L���þ[���[I_�����JqA�]����/��2��l���m�=с!?�+�>��r>�>���>p����J��.Bv���9�������lM��g!k��.��!����=/*�iZ*?��>Aͼ>��>42�:�HҽRҁ>r��>af�?�|>�Q{=�G>D��=Z+�=-<>܍J>_K>0J|>U��=8儿U����0:��KS�:��;�`C?��\�EV���_3��޾ō���>t�?\R>Pp'�u����y����>9C�R-`�n�ǽ���Y��>>-�>|��=�:����G�s�j��P�=��>��>sX���������r�=��>��Ӿ��=�~>Y'?�0w?ޭ6?�z�=Wt�>��i>]A�>	�=�O>�}K>�5�>��?�r8?/�.?���>ꌽ=�6`��=��:=T=�gE��ͬ��\̼���h�<�����A=F�q=j9%<B\=]�==�Q�����;���<�
?��!?J>�>��>�i�C�B���T���E���(�&�p�Z��=(vN>�Ķ>�?k0?˾�>fS�=�!��<�����>?0H>=W��e~�ܕ˽Px�>��=��-?x E?�2>�ᑽ���=�H�6^�>� ?{%�>���>j�>�Y����.׿�C��p7�����=gKA=��>�!����۽����oE��O�=uS/>ἄ>]X�>�4I>��=��.>[=�>5�>EA>r^�=�����s=ڃ����(=1���pG����1��1?R�*ߜ�PÛ���[��۩�}���'�K��'?�-9?�f�gd�q�z�����	����?��?I^'?pB�>�h�>����YU���>��
���>k�?��%?JDt����=�e��=K�R�>�j�>��=����7(�����0���֤?��Q?e׀>�|���t��뗿v�8�q�?�	+;��뾾4�?K�?; ���O&־!W��4�;̽�Z���b������J�n~���)龟/`���=l�	?<�?�!��7��=9z��ǖ�R-��>:��@�y��L���v�>J�	>Y�H�Յ6�~P����Ŵ=��g>� �>�K�=?��>ó�>C#?�t�>�#?�f1?���=R�C?G(�>�k]?{�>T��>�p=�>�O>��> V�\Q>���G���Y�ǻ��F���=9�>���=-�^�Z=�Ю=EP<֬�A�V���=@��=�'�=/��="�&>s�=5�?L/-?ʦ$���޼�ן����=K�L>"�Q;�:�<�0���U�(�a>0)�>8?o�?A:�=3�{��ξ�T�[>%(?ak<?���>��0YT>����eR��d>O�>�(��S�X���/c���r�={��>�i>�>���>C�}?S�&?�B	?Z�0�+�2E�ۑ	�b.=H��=���>|�>�[�=�����@�9�e��J��=�����.Ā���&=��#>M܂>�*>�>>��.>F�b=���'�� �>��C�>N�>�v�>�<>��=���a�ؾ}#G?^��h��ؤ����#Y��C����>��ؽM��>D���v[����-a��?SL�?Y��?Kk?�r��F��&��>��;�t��Ȅ>|�=��h��~���$�>S��>1�W���4�=�x�>=��>�O�wO��.������<Ļ�?KT�g������ o����H��l��.�����~�޹̾^ڛ��ş�˖2���k�?�����Q^Ҿ&��X��?2ez?���>�I�<C��e���G���P>�4��s4��Nľ��E��yľ4�Ⱦ�پ�,���-�d^4��[����>���	"f�B{��n��,2�=��r�)AG>��U8ƾ��=��L>��>q��>ف������˟�)�U�Y�??��/?�$�V#�'Zg����>�(�>��>5�P>	�����轆C�=I�Y?��Z?��1>����/�������?ZB�?�ZD?�?��Ĝ=�B*3�;�>Ib>>�b�<���=��;�s߾Iƾ��s?��g?��?/�Ӿ�F��"kP���>��?�=���ʏ=q��>��?�d����	�z<�>��
�X[��2�=�U��c���ե��^���IW<?X�>O'�>𦺾�N����>A�龸�N���G���������<�y?���t.>fd>'�>��(����i���| ���L?�>�?�S?*S8?i��U�쫽���=똨>���>���=�Dל>/A�>���$�p�?K�By?#�?O��?L�Y?��m�1u���ᐿ1���Dh�%5>�F>���>�%<�I>OI�=㹄=	�}<�]=���>�1g>�W>�N;>�6>b��>tv����%�1Ē���n���~��bS���i�����呾��.�dP��)$�g�L�zj�H��ËI��rk���=���|P�>۬3>��>�=0ټ�/�mh��z��f����
�|�F�h��O�H7]��	>�K�>/��=�b��zV=�)���5�>ӛ'�1ߖ=�+�>ieѼDe�=E4>�)�>�ě>$��>�m��ޒ?>��>F��>,�>el�>�֓=�X�=R�>��h�,xl���E����~_��?l���о��>��*�,4��E�>�7?���>�@ʾ+��G|K����>&E=H8̾7���nH��v+>�>�>81>
U>"1����K�Zf%�rC�=r>+�>:��	ӽE6r��	S=�q�>�����hl>M�>��(?a+�?�;?���<�;�>�x>��>ȁ%=�&�>#SK>�~>)��>��?M�?���>S�>"�����>$4n>w��Q�D=����� �U����vy����Ao�=�П=(�ʽk}���G�P� ��W����Q��>mr8?~5�>���>)K^�`�>�8&M�(O(�h��=*���3�>Ll�>Q�>���>EV�>�i>C�z��þ�e־��>Z�L>jqe��{o�+�ļ]ch>��d>�aL?<�9?�ȏ���d�@b�<���=_Ν>i1�>j/?��>o�(>���B��Mjӿ�$���!�����v�qW�;C�<��/N�iD^�k�-�E���`-�<Ƅ\>K�>�p>SE>��>=3>�Q�>SG>SɄ=�ӥ=93�;��;�1F��kM=K0���F<��P��2��	�ż̏����WI�̘>�E@�}Mټ# �>u�?o��7��l�������R�%?�\�>��"?h��>̥~>�[��rZ��`���z�|G�>ߘ�?�A?xs�=!^ߺ�>�a㾴��>M�R>��=N�B>�Q��4�<�:X++?f�>?#�?���xFp�>���\v<�
�>	�4=���xq�?�W_?�t��L{�Q+ ���G���F?=�׽�7[�'��0�!��9��U�����g�s����=;�>벤?���E�=�ں����a��"U��Q,q=�]=g��>C�D>g'5������aҾ�L�q͜<C�>
��>a�$=N�p?��U?�ue?*fo?f�?�_Q��� ?/3<T|??'x�>K�.?� �>��>#3x�� �����E@����5=T�����={">-�[>^�]>-.�>�[�=��<F�+���Ҽlk�*˒�R�<�V=%삼Hf>P�N=��U=���>�-?�P���w�7��=��T�lHj���_>�K>�.>��I�/>��><N!?�/?���>�Xi=i�����Ʌ�:$^>
+?��N?�{c>�Rd��n�=ٹ����h�����?Rb��6�y������h�H�C;�y�>e��>��m>o�g>Ҕ~?�WB?:�!?����.� ;w�� +�%�����?��g�>���>M��=6۾q�6�Hfs�'�`��m1�+9���F��y�<Be�=�>7�A>6b�=;>�=ٳ����ٽZ%+<�N��侮>�	�>�:?F,\>2=ڪ��n��o2?aZf���=i����Ծ�����=�A>,\�zk�>P�C�I��*���'<����>�_�?��?�Ub?��P�m�ܽQW>��
>�>��=W����!�=�|
�>��!>�xT��~���m��t�=�G(>[�����&,��+�1���ſ�1z�]�� m�c�1���75��/����rB�e*��z����޾��^���^�x���Q��di���Q�k?�
�?�D��
��<��Z��r:��7������̾����+�����UgоǸ��Ʀ���๾����F�"�>��X��#��*'}���(��Ś��=>�n/?1kƾ?˳��z�Ӧp=,C&>	r�<Q*𾬹��㟚���
��W?��9?��쾂����1���>�T?/2�>�Q%>H����{��>�}4?�.?��߼Ꮏ� ���	���ۻ?d{�?ے>?jZ9�p�G���?���=��>i��>�?��?��{��&��h�I??V?��?=�#�7���ۘ*���Z>��(?,kC�}�
>�?->Mu�>�*U<�ڵ�ٰ�=�������=D�B>X�X�C�<�ש6��~��Y�>��>��>�����JÝ>�i쾯�+�H�/�a��F��+�&�û�>�#����=��>�Q�=��5��O���̆�B~���H\?�|�?YA?��@?�y������"�I�>Tެ><W>�C�=�/ѽS�>���>1����a��p� ?u3�?A��?��L?tEk��cӿ���F���ⴾJ��=���=@i?>�x޽-%�=�OK=������C��>�9�>�n>`�w>��T>��;>�Q.>?�����#��ɤ�h����AB��������5g��i	�J�y�P��u���m2���y��a��;����xG�:���=��#���k?>�D?��?.��>B���μ?>�{&��!$�5ӈ������<�F���ݾӤ��B㽄�򺻴ƽ�R������]�?��=�"?����>-���gow>���>��=!��=R��>���=��=��=Kz�=)Of>#�>ۆ�=N0\>�Cj=��\�W������<��ɽ�=�?9���sr���I?�S��>���d��>�?~��>��/�;�t��>p~���v������=q��>�6�>J� ��Jν�'���<�ֽfJ>ԑ�>���>���%辒���6x	>>��>�E־���=��v>��(?��v?��5?)=���>��`>yÏ>l�=:�M>��R>�u�> �?[.9?�e1?"��>��=a��<=�>=%�?��U�g����ۼ{"%�;O�<��2��MI=b�t=y�<z`=L�?=>sļ�q�;��=cX�>�|?Oݒ>B��>�8��S��_V�]i����� ��ΥC>
b>�:�>	\?�?ވN>���x0�zd+�B��>��S>VQ��M��������=%W�>[�l?2�>?ʄ�=���v�	>��J��c�<	��>�?yS�>@-�>Π�0��mӿh$��!��삽9J����;�<�@�M�Iǡ7��-�(���Õ�<h�\>�>�p>�E>�>�;3>�R�>XGG>�τ=F�=�9�;�;��E���M=d
�C8G<�P�����e+Ƽ՟��p��5�I���>�r:��6ټH	.?�?����u��1�~H��<��'�?���>Cs,?}��>^�u>#����d�@�U�=���v��>��?�?B#g�]�=�VŽgh��3C�>t|�>�_>A�C�Oq�z�����=�H9?T0?��>����]/c��Qs�������>���,���A�?��f?!��4���f��3=��������,0�_�V��_���!�[�>�Y��/[Ӿ�]<��N�=J�?I4�?y�T���;EЭ����c4���3��Z==��=�8�>���=��7��������K��s��\�>.�>%�B=��>I��>�_?<x�>M	?��?֞P�~h;?��l>�T?F�>��'?��b>��>S�=F�>�i��ú����y��g�;�6�<~L�=F}U>�x=�NY=�:>�<���<.�=������y%��t�=ϣ�=�˺=O�=p�>���>��?n5��ϓ��R^==!������=
��<�=%=������<���>;�>�/?`�>e7��ln��	���d2�P�=>�0(?��7?wԓ>)��]��>S�p�����5�o�.��>䳰��y��<�о�fƾmɽ��>���>Y`=g>!�~?ضA?�U!?�����`.��t��*��\���)���>*�>�C�=�/ھ�6��"r��_�s�1���J���M�J�=��=�N>��?>�K�=�9>�6={O��ƫ�wnl<$ؽ�Yw�>i��>��?�bY>�T�=񚨾k����?���y����������^��#���>�����>�:����{�4�����$����>E��?r�?@hE?�����b�Uq�>P�>:=�cL>x
��,ϽK�%����=o�W>(;x����n�=�_�>n}?�<�=F�����\5ͽ�ֿ֬���=�t��@���'s�d[4�
vK���P�����󰺾o�2��H�W���]�X&����m���쾡~龎�?�?�;>"��=ogC�"�F�P���ľ&���پB����@���^ƾ�Ԅ�&�����*����;P���w�>K�P���|������ɾ�4�=:���$l�>���j.˾�����	�3�g>��x>9�~�aj����6E��ZP?�,?���`����� ��R3>vb?�ڈ>�ю=y������`�>;1,?�E?�/�=/N|�����&yi����?���?&�S?N��
tE��*0�ܤ�h?�O�>5�>��E��5���g�M|B?zgS?=P�>�M���}�)|$�u�y>)�X?�U�� �=�w�>���>c�n�a���>s�M��=Y��=l+���$�oV��Y߽&O>���>�u>�N��g.��%�>�k��7��	#�"_��J��������>�����=��>����P?��ʔ�{����S=zS?)1�?g�>? -?��D�Z���ޥ���>-b>ڈ'>gA=pD��߆>:� >��� 0������?�_�?k�@���?�p}��߿�����]���q��,��>�v�=�k>^��=W踻��=�)�=3�6�
O�>�8�>�,�>��=:�>!��;�h�>l�~�V�'�=:�����W��(���v��_v��	��$�:4�C����/0�*y� 6�g	C�D��*��=����4u�=��!?�_�>$%>>&�T>e�6=P���o;;����ھn��T��^־��޾�;��C��q0��[*���i�3پ���>�q=+�K=D�>��[=
0:>,W�>�o7=�*U>��>CA&>$\�>8�M>�>�b?=��>�>���>���=Z�������0r�[l"�$�>�e?ZF��ݾ2�j�D�|�|C	?�=?���=4c0�6��{є�Hm�>�Ԓ<'U����l���K=6��>|��>���=T2>�]3�Ugc��Aʼp�;s�>��>�=�J�Rxo:�5�a��>�Ծ$_�=0�>I�*?3\y?ҭ1?�W�=Nb�>0dU>��>\r�=��X>��U>���>@�?eP4?�-?�*�>���=��X�,u"=�J=M(�dkl������w���-�(�<�3#�~�c=��l=w�;�.=~m=G��u�&��' =��?�+?E�>2mj>��������y��d���D��>	�?�ֵ>]�>���>��9>�l½&t��O�J�x�{y?���=�\��� ��:�;���>�)?⌐?UN?�𾾠`���\�=���>��6?ӱ`?)0%?���>��?��N1�D�ĿK^2�}�)>δ>�ս=�
��4��>�>k0��_ӽ�8�>�0 �s�e>d
>V��=�ļ���>�v�>~�>�k>�a�<~�ڻ�l=�U���O�:�"�=��5=bQ���p�=�6��Y�������x�=Q�[<==���z$?4�?}h>
�
=����X�&y��w8>F#Ѽ�2�>GI�>�8���(5��h��V��r���>^t?�>�	��8��=���>�%���,>_��>��E>��+��=��)�ƽ8��=�I�>�G?@�>���=؃��3�����r�>���=�<��?��M?Lx�Y�������5�|�Ⱦ���=������9�F ��C��]yJ�b����L//�j>�v?y��? ����&�=�cʾ-J����C�ؼ;���ߜW>,;�>ܡ�=.�[������Q)��*��<8�>���>�T=:ٛ>)-�>֢r?D�8?�\h?��>�s�=~N)?�����
?���>�?H�)?�E	?��A>�?y=&_��V>l�k�B���/=N,=��=��>?�m���d=f�+>�>s4�<�CR�K��nɮ�E���L�+�<��>>�.Q>6!?!�T?���;ޣ�c�F�v�þ�	?~�=b��<xo��#�> ̑>pb�>
7?T?��>�H��f���ɮ��w��b>��)?��Y?�_�>8�v��L2��=��{��Ԥ�k�->�ڑ=<�!��NӾm�����=$�{>���>>:@�>�xd?(l??��_�g�0�B�o��l���K�?�>�t5>�	�>���Î�O�ʻ��H�g��ץ%>'�սA?<ǈ5=���=j�C>�(�q��>�B����<\��=�y&=�(I=Ӽ>	k�>\Դ>8F�=U��}���$����F?�X�=���������=v���i��^?Ƚ��}����=��*�3����V�r��%�����?��?���?��ؾ�$M��%7=��=�q<>LA"�*:���v��N������=�q=jPҽw���3>K�->���=j�Z��>������7��hu����D��@b�~���?��ڀ�b~���ɷ;�CĽA���� �F�X+?��g7�n"��I6�F�y�����6pž���?��W?�j:>p�> �5��������ܙ=����� ����о�d�������n��$���%�.��c��Ǜ>�~Y�L:��&�|���(������?>W>/?YDƾ/״������g=$h%>t�<� �F������-��NW?��9?>�"'�����>��?
e�>�%>3�����;�>�-4?f�-?���p���2��/���wj�?>��?M@?^I�^bB�}�����o�?�?�j�>�e����ʾ�G�*?��9?�@�>E+�fބ�����>IcY?`Q�*rc>�0�>�ٙ>���N���w�"������Ns�\=>���<��f�OjA�mh�=t�>�Dv><�X�YϪ�q��>�¾D��>�(��f�Wt��~���>��ĵ}>p	�>(Ϸ���1�H,���ꋿs缦�S?�1�?eQN???-N�������%�K2>�$�>��>,��>D�׽�I(>P�>)�������n̾ڬ,?�?A�@��q?LO��Ŀ���W-���/�z<>���=��d>;�C�:�=nZ@>���=,T�=�EO>��>��><�>ʳ9>��q>���>��}�)�z<���Y���@��c#�(��AY��c��70�Y��;w��]�����k�����P��L��J������S���@?�K�>�J�>���= ��=��߾�~)�����쾖�"�"A�h��`���־5�Ҿ�ܾM��b�J=�<��,�>5aV=�!P�M��>�>�$>�P">ؚ:>��p>	�>���=x>�<���= b>��=N��>O�
>r��>��=k���]e��Hv����=�R�>��s?��">.��WwL�!�!�������?7'?�J>B*8��j���M����>܋q�����l�H�D�]��>�0�>�@=4a|>��E��];}=�L뼑�[>k��>�X@><�1�:D����d��>�C�����=o~�>�2/?��?<�0?���=���><��=Ƚ�>���>aݔ>	q>��=�?Fh=?	�Q?r�5?;[>���\��<_8<���x�=��׽�~<U�/a��CW��N�>�Il>~��<2>,o�;����
!�:�(>��?ϗ(?s
�>ix�>��ľF�$� _��Q�<>�V>��?r��>4M?$C�>C2>�7�rT��_��Zw���^?���=�Y�� C��y�B�o��>�2+?fM�?O�]?���Sg@�%<�=�>Zy9?�?�%?K�>��!�R!��V@��ܿs��b���޽�&�<R'�=%�n�Q���8>F�K��@��Ǯ�=9�0>*�_>�
_>�?>˞�>vQu>C��>��>�<�=�4>�#=���=zۮ�fts>0kY�漛�]�0˽BO���,�=�)���ֽ�Q=(��'�9��#?l�?,>f��=e�� p����4>n�9>���>t�>��!>�.�s�e�Mm;��n��/�>�Ax?��>�O�A՜=�uN;(><�P�>��l>Zx�>�h��bg�:��t�>M�>C;1?v��>+Ny��]��S`�ϊ��S��>BZ�<���ɧ�?��D?zo�����R�$�:�e��y1�\Tc>��'�q����׾\�R�F�H�7}����R�:����<>��><��?��i�j��=Dqվ�ʄ��+Y�BHl�C@=�_>�I?�id=?%(�����<i�8�P���@=׿�>K�?���=��>,��>U?�AA?T�?	?�B����!?�,S�):�>�0?%s#?�g1?���>Iĵ=ޢ ��+��k�>��f���M,=ƛ�=�M>�Ͳ>��p=͕��=o��=u|��K� ��޽|/>���<�\､XT=���=U�>m "?�	=?�T���䜾@�=P���0<QR�>�|�>�8�\�U>#2����x>��>0�>���>�Z�=1	�V}�я ��m>l�4?��9?ʻ�>Sp���2�'2���Ѿ���>hu�>;�Q���u��e�r��e���a�=��>ۙ>;�i><3~?�=?#$?�(�v�2�:n��,�]�^���<Yq�>w��>�z=O վw>3���n��\�|m%��漍(F���=�g>�*8>�d(>.)�=��+>��<B�r�7]��&#<�V�<$y�>.�>O�? GP>�A=賏����;;?�L�<� ���9��=�=c���ȼ�!��>/]���=�=�ھJ���m���h#��![?Tu�?���?>h<?��9��'�;�m>�{�<Tc�B>{�4���C�������>B�aW���C���%���>s�>��<�i���-��([�ζ�I�X���{=H���<g�4������ �Hܐ���-<����z�\���_���B��Uԡ�����ʾx'��hD�?_%}?!�>;���k�����=��  F=�¾��Q����<ݸ�zK���S��V�������P�~DQ��XH���>fWY�II��/�|���(�ϋ��C@>�W/?4�ž<�����i=��%>���<������g���Bu��W?&�9?����8��'h�Z�>��?���>��%>�^���}�Ą�>74?B�-?Z�N���'��W/���T�?���?.�F?�;�zMM�����e�.q?0?eH�>4���۾�#�$�?��=?Z;�>����pz����T�>�A<?wR�5(�>��>&�}>�*y�0���L߽���D嗼��U>��<ij*��w�w�r����=B�>ӑ�>r�L�l����Z�>�3�����(�2��~#�l������T�=??,�H�>\��>Q�d�M"T��ᓿ�3���{���U?���?lmB?׃??p#��<�Πf���>��=m�O>�o>>�m/=���<M�>���� j��#���a>+�?�@�K�?�����Ͽ�˙�Ū�>i���� >�8>�A>�6	��Z�=};=�����b��=�/�><�2>`l�>y�$>rU6>�GK>{����)� 槿ť����8����q��ݕ���/ap�#��M���Xd�����x��r����X�胳��Z�:�پ�����8?�vn>'W>��=�C=��B���&�:�)�Y��.`"����������ܾߍ޾Yl������򗾂\�</ߩ�e#�>}*�e�X��Z�>�%`��cP>���>���<�
>���>�J>|~>���>1�S>�`�=��A>�c,>S��>���<O��򴁿w�U�R�c>�>�>�,b?�ٰ=�����U�H���5�u����>�cA?q�F<y�/�������9���>�${���N�w�>q�w��>�z?�}3=$,>]�n�;D�й$=�v>E��>P��>�Pe>��h�ݍ��{��ZJ�>�Z־�=<[y>�)?i�v?~�5?� �=���>�ta><��>x�=�uL>=�Q>�a�>�?K9?�H1?F�>V��=��`��v=�!;=��=�i[V����3���'����<�(2���C=q=�<��^=YgD=�mļ$%�;F  =���>�:?!��>���>H?���>�.�E�(���>��s�>T�>�L?d��>uC�>4:>E
��Aþ�\;���>�pI>�`�)�u�����=�>�O�>	AM? 2?���+j�G��=c��=�ݷ>(�	?J�&?��>�>����N���
޿�^�#�6�Ĵ�b���C��>G��B����	>�2��5ü�Kk=�.�>���>��>ܦ�=��)=|�*>a}�>D��=��>(���|=�i�=�	��*3>Rz#�ws
>�U�S=ׂ���6��)jQ��n��A>ҼcYL�eIL�b�#?��?���e贽y���b0��L־E�?��G=��@?J�?����I��HP��V�����{B�>��[?�:?���;�T�=��v�xh��S>�ћ>G��>�J2>�*X�6�X��n�=R8?J�?��?�⫻b�~���s�%��@�?8��6��3�?f�:?,�#�bG��D~/���"�eQ$��~#>\�#�YI��Ĺ���5�h@2�oY�*��e�Y��>+�?yP�?q{����,��쾄ӂ�i|��3��3�=Jp2>:e?�fJ=�HY�<�P���ﾓt������>�>nd��h;�>_� ?�N?T�o?�M�>�M�>4���t�?�޽}�"?�V?$?�>Y?���>��>	i��䈺�.�=)ýmu��N\��f�*�A`�=�6�=�G�<�"�.҇=��=��<�7�����hԽ<�3�|q<+ʠ=�5>@h�=�u!?��I?e���F�=~!=�1���mJ�>h�#�.tǽV��<W�7�*n�=�p ?�M?�]G?o�>�[�ݐK��[9�B�%�"��>˺C?��2?]#�>�"��Sv�����4٣����=y��>�}�<3i��\��V���p����%>M>���>�$f>�ƀ?�;A?ž#?�����/��bq�*�-��v��+Sռ��>�5�>��=(�;��0��-n�]�`��M2���;�'�R�5�9=���=�>�.J>�A�=�>G�t=#EZ��L����<�պ<�>(-�>�l?w:T>��=钝��' ��.?�N|�I�"�ȹ�Yx���7�������r>�c ==��=;��x^���䘿,[���k��%�?u0�?��?h���z�)�">cOV>i%�>w�d�Z���<��5��=�=>h�'Q�2dp>�i�>��x>�6��`о�`��A��}߾�	9|�*�*>�������о7CԾ�	��K�\=ư�<x��໾����K�#�;�װ���羜o3�t��?l��?Uħ>��1=�)��7�	�Ǿ��==�����%�MJ� ƾ�I��k���\�P�vt&�����9��ǹ>A� ���~,���/�@"F=�1>�[7?O&��' ��kS��_�=�7J>��S=ľL��	I��� "��Y?�5?o����"C���}=�?��>V~">��O��'1��7=>��;?�T0?�ġ=��|���{�?����?���?>�b?t�1���y�Y_�᱾?�>?P7L? �'?�9<J`!�V��;)?�G?�?��a�|���)�w�>;",?[F�
�>�3�>��t>�y<��r��v;!������>9t<�{�:v�����Ό�>P]�>�i>�c���_
���>'������0�?2�k�\�����b��>f���U->��>�mG�Yt�dܘ�����ydн�EG?볮?�1?�G?w���1���)�V�=#�9>�=>�������BM�>�.�>4�
��`{�>!Ծ$(?|��?��?��j?A5X��Dҿ����������gm*>T�=|D>�r�����Ij�=��	>3�<"�>tk�>m�<>�,w>���>�}�>���=�j����%�^������v+�0���c�����o���M�-���}ľ粴�3�[�;��:�����I�$o̾���<R?�r�>C�>N�>��=n���������y�;�D+.��W�H� �W��Q���@۾6�ﾖ1���=�rоԿ�>Wy�A�Hة>7��=b�d>�rP>ר���=j��H�>N��=�|=7>u�=?eI>�9,>O�>Ļ�=5���d6��3]� ��/�??��_�꟞���3���⾞밾hx�>�?W�e>�E#��.
v��W�>��6��g��"½?���ˈ>a��>4U�=s��;���v���ڽf�=Ä>�v>#儼�������J0�=���>J־]�=�xx>��(?4�v?_�5?���=���>��a>b�>M[�=�K>!P>�V�>�?Z�9?�1?Ir�>J$�=H�`�.�=|'9=M�>�W�G�����ox)�-��<b�1�R�F=��r=��<��_=�U?=��ż���;�& =]��>>~8?u��>��>�Z2�!@�Z�M��I�{�>��7��U�>E�>�?/�>r�>?D>�n5�xž!�߾@ �>��A>.D_�M�u�#�Xx>�s>�HM?��2?�n�)�^��=m��=��>�?V!'?�$�>o�>�0���J�!�Կ���#�"���m���F�ώ��R���g�>������-N=�u>���>�Lc>��>�	_>�=>���>�u>#M2>ᚮ��*/�63|<5���_>��4=�p�=��4��>���н��@�L�q��)'�k��?�Z�A=�B?��
?�m%>ZsK>vߎ�����t���+�>6��>!v+?j�<k��=�%��+�h�zr]�\�<��'?Č�?��J?�	=��%��Խ����|�>u��>�?�[�=���XM�<'kQ>���>�^\?J��>��9��Tw��V�|�W��?�z�;��[��.�?9?Z���D|�^&�")%�_2�s��<�At��$��
���=4��H��s���6o����=��??�?~)�����=����8ؕ������ξ�B��P�>l��>�b>���؟ž���AI��4�/=�wr>�F�>H
Ҽ�g?��
?��j?��4?���>�9�>�o����>��ɼA��>���>[�?P?c�&>���<(B½�&��>�"�{�/��G����=V>��>!WF>���=��=*�>�!�<�7�<�=@.����i�`�< =j=F}�=� >�k�=�?A�N?=#�=����Z�>{�N���w��=G�=av\�(�d>���;%T�;��?C�<?l�>��2>���X��y�+�9>w� ?�51?��=@�-�������
�$Φ���&>�3&>v�0�b�\��׾�1��R��.T>�n�>c>=:�e>M/�?X�5?��?V���-��e��4����2O<���>�m�>*;>S��E2�I�j�Nb���-��֍���[���D<��&>%gJ>� >�
�=^s>�1<@Ä�S�$h�����<���>�#�>O� ?��O>#�=�@����۾�:?r�x�����O���Jg�&ľIヾ��<Y�Ѿ��=6�H�����^����.��"4?Z�?���?:]?]
�����>V_;���.>�Aa>��
�ӽ��p���>h.��]6R����?�Ú�>��>��=L9��'	�ř8=�d��1�\�;�O=��վk�{��a����˾e��|C����=�R�g ��N`���r|�9����	��F6���Iپ����{�?�iq?*T�>��-<L���F�V۶�`:=�ߺ�+nG�(׾�zw�nИ�-�Ͼ���/<H��0�Q��d��>��5����}U��>�*�beλd��>!l:?3{��C�;�������=�u�>�?=�b�E�������֥�Q�{?�;?:���6�.IR��S >�,?&�?�nj>��?�.e|���>�P?��2?Nt�=~}�7,��ߩ��'͢?���?�[p?q��j����W���?�C�?@o?��>ֳ%��༚�o?�F?UP?�gr��q����/���>�<8?i��MI>,��={t>8V>>
<�T���bD��uμ�d���}{��_)��u�	�3��Q�>���>�Yz>�yž��9�k�>�Ⱦ���F�(�q���<����@��u
?��!�>La>m.>jh����e쒿:������lp[?&(�?ջ9?��F?�����^�3�*��>�?n>��}>�P�=D�x��d>�#�>�����L��Km���u?l>�?K�@��Q?�iR���տ�����C��@=��YÙ=�y��I,�=��뽢�<X;K<��\=)�=B�>9�>��>E�>E�a>��0>��>w��w�!�]@���@��.J>�,/��Z ��Ռ�v**�L8Y�Wh�����X �������p��K��*�����1���u����>'r?��>��>Ҋ�=䖼=ҧu�����5�2]�^�!�J���	���׾����}���6�,Ë�S ���޾�H�>�DA=D�G=��>$Z����=�ȭ>���=��B>�1>l%$>�=c>�G>�>��>�FY>��!>�ă>"��=�{������0��d���U�@?|�a�B�����4�x�����$��>�?�+v>S��\��d�u�g��>^G��H]�˴��I�M��X�>���>�D�=�Y�!���QBx�&��=��>k�>��G��Ñ����.�=H��>g`־?B�=V�|>"i)?�Fw?��5?��=��>��_>�ѐ>&�=a�K>�kP>��>�?Z29?�2?(��>ZM�=��_���=
v==.<=��I�{-���`��<�(�^\�<��2�b�O=��v==��;y1]=�ZB=��ɼ�μ;6�<��>�8?���>S��>��9���>�,M�v�׹>L�����>E��>�r?X��>_�>�f5>�\���¾���`�>��@>��_�"�w�����x>�]s>7_O?��1?��f��Ob�Ʌ�<7��=�>m�?t4)?`û>Ƞ>dZ��D�j[ۿ�L���EW�=;�,�<,���$��_/�c�>�[=b���Ȗ+=�sb�=O>[!>G>�Y(>3=�>xY�>�=��>MM=rT�=��>QSW�\->W����=8����� �O!Z��*���S�n�<ح�<��W���
?&?U.�=7=>�'
�� �o ���(*>��>}+?�7�<hq����1�h�}�]�`����<�>GJ?K�(?��=�A9=鳭��s����I>[��>ڭ�>��=kf�<ec�j+�>]� ?�Ug?79�>��h�w�n�^5g��ƾJ�$?�kn;q'�~�?u�N?L� ��"��a�����=�̈́����7�����8���1��������Z���;\=z`?md�?��k���	>����}��jo�cR��|M3<'߻=Ȅ�>q��=[t�AZ��8"������=�b>O+�>獏�G�>�g�>� e? XJ?i"�>>�>��޾��2?�.�O�:?�+?}3?�?�J�=���=�ؽ�!�=I��3�P�r��=Ff2=��(>��<>��;�b!>X��=�&�:� ;L��������C	�"��<M�=��=��I> �b>�?A�]?%��o횾�V�=��?�+cE>��5����=��@������f=��W>�?�a?9�>A�:��V�W5�D�����=�BR?�AP?��>Dy(�j��6n4�)3����[>���>��E�=�QžZP�4�p���j>��><��c�j>�}?v�@?[Z"?���h�,�T/r�˫1��a�Ӱ���)�>ST�>�,�=�!о�6�07p�z�_��1�%׃�.�H��@�<F�>@+#>�M=>�\�=-�>��=^L��'
�D�C<��+��L�>�]�>d�?�S>*:k=d2���A���	=?��<)�ݾ9բ�����G0оk�;BҜ>cP�6y">��Ͼ�e��c��Uf'�z@i?��?��?(=�>U���	���.9>��>�{�=5n���i��&����B˽���>`a>��{Ⱦ�:�:���"r�=�nV>������̾a�̾C2���@���eo�E9r>5ݾ��鑽��սD��;7ؽ���i@B=��־�����p�P�������������~��2���X��?��?��!>�K�=�����aې��>:�r����_���۾z�O��m���#��,��D�@���)�K���r�>E���-�������[/���>�B�q>ވ6?2��V�;/ ��M�=�>!I�;�}�j%���o���PN� �?�8?�=߾��!g���V>pi$?X� ?׌�>&��z�����>��c?~<2?Z�>Q�s�d�����ý�c�?��?@l?�9V�®���� �v�PCs?f�?�S_?�Qo>�KQ�#lp�@~_?�<??�E?�����Ӊ��E�5��>N�@?�%B���C>��=��%> <"�Ľ�fm=5Ϧ����=; ��ķ<��2�X�徖e�=���>	�?7�M>crܾ�I�5��>���,N��I��������<��>����Bh�=��a>[�>!)�?W���'���$�D?z��?!�R?�T2?�G��+��xf�>�=�۝>|L�>by�=}p�%�>��>s�߾�q��v���?���?���?~�R?�Hq�Iӿ�
��������)��=2 �=��>>i�޽h˭=-�K=����=�'z>��>�o>f8x>�T>��<>~�.>�����#��ˤ�ؒ�xZB�3�=��eg�x	� y�ʡ�ʴ��񽾮���	���nԓ�*�G���=e>��Y���y%>��?���> (�>K�>w�)>J�����3�p�"���<�����wF��Ѿ*؁��-�	���Ј����ƽ����?��<=1��=���>�J���(>�f�>B��=��?>�V>z�9>�l�>�%a>�&]>]+D>��H>�r�=I\{>Jf�=&,�����.w:��.Q����;�C?Cw]��q��-�3�#o߾d���{�>x�?j�S>.�'�������x��>
cH��>b�p�ʽ���9/�>���>�=�=�,ػp���w�ܠ�P�=]Q�>y�
>�k��ӏ�i�F̘=�B?	K���=��E��>TNR?��W?���>C�?��>��?}u�>���>v�>5��>֢,?oT?��?�q>T0N=i߽�R�nB���H����<��=�5=�j/�w꼔 �x=vM���꽈؋=el����0�[+�=3�|�N�>15;?��?���>F���#��$�_�D���X��=F�?�x�>�q.?�@�>[T�>.=U>����&t�K1�:sn>E/k>�1���n���`>(�>�[�=��?��L?�x��������`>b�9>���>�y ?�Q/?~�>]M�=%"�fu�_�Ϳ2���0�ڲG�+�e�Y�3=�S��G�����Ž��B�߈�n�;,|'>�0}>r�j>z�S>c>�H1>�D�>�>>2x�==>+܁<c�~<
�^}�<�%�^���4`�xE�3��M�`:C�ݽ�3��M����ǼD2�4�>�O?��ל��I��񴃾�|)�)����S=3�
?�#�=� ��څ#��`%�$.n��u#���>{��?�a?M:��>��)�ɽ�Џ>��>�� >���=S�������7>=�X>KV$?�̊>"��<CM���R�Hľ��C>�I2�n�A�t�g?,�z?�= ���-��I�Z?�"愾�L��HѾp���՞K�2nM�^�ޝ��'��/f�=[9�>���?��#��1��N��5/x��������ҳ�RxúMB�>X�>r���Kɕ�fh�x. �gʋ�Y��>s#�>T�n>���=U�?���>.'k?�I?�v�>6ӌ>�G?h�]=���>=?�L?��??i�>'�>2ܛ=o��Mr��Ѝ�*���#.ӽ����R'=��$>L�=���=��W<��=%�O�T�|��=�.��T-=慾=,�>��8>��?�?k��=�o�<xI=<rü4&���7>���>E�d=g���+�'>z��>٫�>��G?�$�>q��=\9����:�"�и�<�w�>1�?a!>?�a#>��@>7���+=zW{="~�c2���d��;g���t½Qi�>�_]>��r>�>8�i?]�6?%�4?b�����.�'�4�m���C
�z���̘>)�=��4�~���=�$k_�Y�U���9��Zy��� ���>�F�>�k<�>�4�h>�ˆ>N쟽��]=L�k>�m>@��>��?r,?�'�>
Q�>y�о�"*���I?����)l��꠾rdоjH�*�>��<>�
�=�?���G�}�����@=����>E��?���?�2d?��C��$�o�\>�PV>��>k/<��>�����y����3>���=�wy�����B�;.�\>w�x>m�ɽz�ʾ� �*9H�	�ο����_�g���������*҅�8���?�<�F��s�I-㾟��8~��ޒL�T��ם������$���-�?6�>�d��o>N��6K�E������l����G4�g������=���a�� ޾����-�W�1�.��y��>�ݽ=���/*x�~ ��;1�<Q��>��
����:���P�����~ڽ�G��䐿}G���WͼI�s?��'?TԔ�����-����>��?�	�>4j�=!㕾�b�=a�>1?U% ?Ͱ>Pr�������T=�"�?��?�S.?�o�<�9F���4�����?�?h�>��(>�h���FȾ$�`�-4�>��?�d'>R�&�]���0�C��9?��q?@����i�=���>���>%"-��+���f>��,�[̼6�ʽRX�=#R=|�v��F˾��=yH�>7M\=��}��5��>���,N��I��������<��>����Bh�=��a>[�>!)�?W���'���$�D?z��?!�R?�T2?�G��+��xf�>�=�۝>|L�>by�=}p�%�>��>s�߾�q��v���?���?���?~�R?�Hq�Iӿ�
��������)��=2 �=��>>i�޽h˭=-�K=����=�'z>��>�o>f8x>�T>��<>~�.>�����#��ˤ�ؒ�xZB�3�=��eg�x	� y�ʡ�ʴ��񽾮���	���nԓ�*�G���=e>��Y���y%>��?���> (�>K�>w�)>J�����3�p�"���<�����wF��Ѿ*؁��-�	���Ј����ƽ����?��<=1��=���>�J���(>�f�>B��=��?>�V>z�9>�l�>�%a>�&]>]+D>��H>�r�=I\{>Jf�=&,�����.w:��.Q����;�C?Cw]��q��-�3�#o߾d���{�>x�?j�S>.�'�������x��>
cH��>b�p�ʽ���9/�>���>�=�=�,ػp���w�ܠ�P�=]Q�>y�
>�k��ӏ�i�F̘=�B?	K���=��E��>TNR?��W?���>C�?��>��?}u�>���>v�>5��>֢,?oT?��?�q>T0N=i߽�R�nB���H����<��=�5=�j/�w꼔 �x=vM���꽈؋=el����0�[+�=3�|�N�>15;?��?���>F���#��$�_�D���X��=F�?�x�>�q.?�@�>[T�>.=U>����&t�K1�:sn>E/k>�1���n���`>(�>�[�=��?��L?�x��������`>b�9>���>�y ?�Q/?~�>]M�=%"�fu�_�Ϳ2���0�ڲG�+�e�Y�3=�S��G�����Ž��B�߈�n�;,|'>�0}>r�j>z�S>c>�H1>�D�>�>>2x�==>+܁<c�~<
�^}�<�%�^���4`�xE�3��M�`:C�ݽ�3��M����ǼD2�4�>�O?��ל��I��񴃾�|)�)����S=3�
?�#�=� ��څ#��`%�$.n��u#���>{��?�a?M:��>��)�ɽ�Џ>��>�� >���=S�������7>=�X>KV$?�̊>"��<CM���R�Hľ��C>�I2�n�A�t�g?,�z?�= ���-��I�Z?�"愾�L��HѾp���՞K�2nM�^�ޝ��'��/f�=[9�>���?��#��1��N��5/x��������ҳ�RxúMB�>X�>r���Kɕ�fh�x. �gʋ�Y��>s#�>T�n>���=U�?���>.'k?�I?�v�>6ӌ>�G?h�]=���>=?�L?��??i�>'�>2ܛ=o��Mr��Ѝ�*���#.ӽ����R'=��$>L�=���=��W<��=%�O�T�|��=�.��T-=慾=,�>��8>��?�?k��=�o�<xI=<rü4&���7>���>E�d=g���+�'>z��>٫�>��G?�$�>q��=\9����:�"�и�<�w�>1�?a!>?�a#>��@>7���+=zW{="~�c2���d��;g���t½Qi�>�_]>��r>�>8�i?]�6?%�4?b�����.�'�4�m���C
�z���̘>)�=��4�~���=�$k_�Y�U���9��Zy��� ���>�F�>�k<�>�4�h>�ˆ>N쟽��]=L�k>�m>@��>��?r,?�'�>
Q�>y�о�"*���I?����)l��꠾rdоjH�*�>��<>�
�=�?���G�}�����@=����>E��?���?�2d?��C��$�o�\>�PV>��>k/<��>�����y����3>���=�wy�����B�;.�\>w�x>m�ɽz�ʾ� �*9H�	�ο����_�g���������*҅�8���?�<�F��s�I-㾟��8~��ޒL�T��ם������$���-�?6�>�d��o>N��6K�E������l����G4�g������=���a�� ޾����-�W�1�.��y��>�ݽ=���/*x�~ ��;1�<Q��>��
����:���P�����~ڽ�G��䐿}G���WͼI�s?��'?TԔ�����-����>��?�	�>4j�=!㕾�b�=a�>1?U% ?Ͱ>Pr�������T=�"�?��?�S.?�o�<�9F���4�����?�?h�>��(>�h���FȾ$�`�-4�>��?�d'>R�&�]���0�C��9?��q?@����i�=���>���>%"-��+���f>��,�[̼6�ʽRX�=#R=|�v��F˾��=yH�>7M\=��}��[�"=�H�v�e�,G~��3��9<�����	�:�7���I�����gkP���p�
A���Δ�3���g|?�*�?�?�6?�P��F�������>==�>��G>�=/��<N$?��>���J;��n5�7(�>���?��?X}e?��9�Ȁ���∿:��{.�����=�S�=���=s�Ͻ��=ZL<P�<-�T;8��=���>I}X>�Pr>�y^>�!#>Ќ9>/���i'��C��2w��A������'��\����;�����z/�p.��ڸ��6M��s����W�� ����l�6�9�ѵ��D~>�i?��>@f>����>Gꊾ�&���x��֙��&��޾�޷���ݾ����pe�s+žSQ�������z�@��>¿6>퇀��:D>	&D=y�F>O�*>i_�=��>6Ӷ>5�>L�&>�H�=KA�>隡>sK>Ζ�;L\|>�{�=���%���R5:��kQ�ɕ�;/�C?\��显Ϥ3�_�޾����>�?	iT>}s'�$���,�x����>�2F��7b��˽5^#���>�a�>ʦ�=G���We��w�K��	k�=jw�>�u>��]��ُ�I-�4I�=k9$?l�������$>3��>�@?S�Q?��>��&?,?��>�ڼ>�>�=���>(e&?*��>���>ꎋ>/t>������Q=�V�<�PH��@�KZ.����<�b��RI�<��n;d3>�N�=�v =a!>>�!>&ὺ|Bp��L}=z�>�Zh?�')?�]�>{W�V�V�Y"]��P�﫠=�ڹ�[?���>��?��>���>�d:>��ݼʞ�x?���>���=��k���Y�fȣ>�~)?8�>�o\?��E?��н;�Ͼ��I>�J>.x>�?�J5?���>��!>�&�=����lӿ�$���!��킽J�)�;��<���M�Q-�7��-�����j��<4�\>:�>$�p>�E>�>V<3>vR�>|IG>Qӄ=��=`3�;��;��E�5�M=x��%G<M�P�����Ƽ����>�� �I��>�%9��8ټ T�>D35?X�z�1�þF=��H��� ��DT=�c:>�Z�>|.>H������7U���^�E�Ծ��?�֌?��/?;���S>3mx>M>��D>�I>*�>��I;��%���|�=��>�E:?`0�=�����	]���Y,� �j>� ��х��X�?�rD?�3���
�h�#��gU��??�ó��q	/�,��\%��`3�ÊY��18���8�����s@=�I�>�͞?l�����Y=mɾF[���g�҂��( >�>d��>�<{>�����r���:��Ey��^?޽ȕ�<
�>�M<�EK>/��>͎K?j^?�?g�>��?D��>&3�>�y?��?��#?Y�?�>�>�і=d����bl�<��t��zqZ��w.=�sb>{;
>&P=���=���<0����@a��	���� >�W��Q��1
�<R=?>J��=�?�y?���1�1�>��4'��	�=|qo>���>��>= ],��$�=^��>51?��F?Oh?�%�=B��
ھܾO��=��?�?�m�>�Y��0=z�羡����)>�N�>#����2���F������tZ0���>��>��=��3>�ȁ?N?�S ?��'��'B���w�j�(����=�����>	o�>	�=I�۾D�1��n�"�_�¼4�A��R�%���=��,>�@>��H>̖�=�~�=a=�<�1��� \=ڿ�=�m�>��>��?�s>�&$=�7�����2�I?>�����x�� �Ͼ�d� �>��;>7g��s?���w�}�/
��%=����>Q�?���?�od?�B�o����\>NV>�>1^1<��>��o�X��>;4> �=��x�@5��Wʭ;�\>y>��ɽ�	˾$侾�H�b���|gy��b�<	i���A��Zľmn�Q�4�P���6�� ����ɖ���Q��Eb���{�C����Pƾ�:����5?�L?��(=r".=Y�=����`��/��$��P�����=���g�澆4����5�B�9�z�(�-:�.�t>\?�T��/y�(�5���Z��h�=�7?dݾ_Fܾ�*��6<��=u�P�_7�o����Օ�Vܽ�w`?�96?��̾Hj�o�J�>M.>��?�>Ã >����@��4nt>�,?"�#?y{�Y͈�����/=sx�?�P�?'@?YQ�<!A���������?O.?��>���Bɾ&b�.�?�:?�E�>�-�����vt��V�>��Y?d�K�?�c>X*�>�ޓ>V���h����9���n�8��U5>I�6�Z��_k���<�4d�=p#�>T�u>9[�C����N�>�8�l�N��6H�[#�^<��W�<��?�K��a�=%�g>�	>�(��=���ى�|����J?��?c�R?@�7?�����|�SU��Y��=)�>�m�>!�=�%��ڜ>��>��rr�6r��S?ƥ�?�C�?�3Z?&�m��/��І�Ս��<�G�:��=�v>��u>�f&�|i9>��=�^=���<S� >���>��~>�v�>q:�>DB>c2>,���"��̙��Ox�;A�<�!�0?�h������w5˾�/��(��-��?�ҽ.&m���� ˾\���k��7Tž�s3>R�?���>W}3>q@ ��E8>�aپk8�S�˾.�'��q�B]���|߾�Ͼ ��Cf�|�y��s���V�;(Vʾys
?O�A>���=΅>?�k<����=�U8>mpt>	]�>�QB>g��>�w�>t��>���>(��<z.�11P>��=��������'� �H� ����N3?�f�����(/��߾l����>�O�>�E�=&A.������T����>Y�:�@�%�����oQ?>Wj�>.�=mp�-0
�z�\���4�m3�=�l{>��>Hw�땾��ӽ����`?�W ��nQ=ƾ�=]%?>�`?��_?���>�i?
*�>Po�>�K�>\�>IA�>���>H?,�j?e�c?u�?��>>E�P�aG8��j�=�PP�kF������>:8;�=]=%�3�.%�=V�:=|D�;Ѡ�= X�=�M�=�">���>��I?���>��>�ھ�F��6�v�]���I<59�=G�&?n��>;��>E�	?ݫ?�r�>���Pߣ��[(����>Il�>~�$���n�.�~�i��>��R>��X?준?��3=��A��?~=�b~>t�>J9
?��9?���>F�>�v�=��
mӿ�$��!�M�Q�K݈;��<���M��H�7��-�O���"��<5�\>:�>o�p>�E>Z�>`<3>�R�>�HG>ф=0�=9�;�;d�E���M=�CG<�P�����)#Ƽ:�������I���>��:��;ټ7�?�??Os�j����V�����Eb��R��>��>���>�W�>���={��_�W�k�C�	kU����>�Oc?��?Ѓ1�0��=#�Q�uj�;�D�>�,�>6X>��>��p�F��R3�<���>?�8�>�b��Y�Am���	����>�0�<R	
��C�?��[?�/�W�x���!�H�G�~	���=Or�?�q�XԻ�m�!��9�^����h���+n�=�a�>�z�?Zt���=��������D����\=��{=i�>r�P>�2�"����p��]޾�]G���=~�>�t=bɟ>7�;?��?C~g?�:?�`?6�-<O�?�>5�>Y��>�s=?��?��?B��>!��>��7>�x���ҽ�v���~�=?�Q=�L�=�>˓>��=��=�C�=ʬ�滷=er/;��#�Z'=a�=�U�=��=4�>��?��#?9|ݽS�O�������h�<�s>n0N>�V��3e�%�-�X	Y>N�?��/?�,�>rp=>�۾* �)	�%��=,�?}f2?e,�>���; �=J_�nՁ��#�='cU>�Wb�Ӻ��Qt辖�������-�>�ύ>y��=��>�x?r�?�K�>`���ٜ"���x�;"�%��\�μ���>��p>hw�<l��h�F��_y�-�_���-�Uh\=!���ۿ<��>�Fx>��=>{�β\>r=_P�rJ�{s�<�Q���m�>ޣ�>���>�VJ>�)&==��Q���J?�ʡ�6v������fо���o>��=>S�9�?!�� �}�e勵@=���>���?4��?�cd?�DC����8�\>L�U>+>"�3<��>�{��mӅ��3>&��=4�x�8��3��;��\>�x>�[ɽ��ʾ�VH�	`���U_��/��R>�gd��Nо�黾zU�(����[�n"�ڿ�?2ξb�ǽ�<��=2�yJξ�}����2�>?�m?4���g[���#�ԗ��	���ɽ�ž�?�:�����������w+$�+�
�zQ;�2G���5���ӾR�=���{���
\��̤ܾ{�>�νG�>�[���뤾�X)�<�Q�졽w"y��q�
:��`���\r�in`?��-?��u��*��ɒ�p��>*��>M�n>KR>�z��[�����>�>?^�"?3��~K��R��X�!����?~�?��9?�*:���F���t��{?�?F4�>�A����Ͼo���?��3?V��>�$
��)�������>&�[?��F���Z>�z�>q�>Î��ؚ�����厾�B��$>�>��(�Li�g�4�0��=�ۛ>�j>?�G����[�"=�H�v�e�,G~��3��9<�����	�:�7���I�����gkP���p�
A���Δ�3���g|?�*�?�?�6?�P��F�������>==�>��G>�=/��<N$?��>���J;��n5�7(�>���?��?X}e?��9�Ȁ���∿:��{.�����=�S�=���=s�Ͻ��=ZL<P�<-�T;8��=���>I}X>�Pr>�y^>�!#>Ќ9>/���i'��C��2w��A������'��\����;�����z/�p.��ڸ��6M��s����W�� ����l�6�9�ѵ��D~>�i?��>@f>����>Gꊾ�&���x��֙��&��޾�޷���ݾ����pe�s+žSQ�������z�@��>¿6>퇀��:D>	&D=y�F>O�*>i_�=��>6Ӷ>5�>L�&>�H�=KA�>隡>sK>Ζ�;L\|>�{�=���%���R5:��kQ�ɕ�;/�C?\��显Ϥ3�_�޾����>�?	iT>}s'�$���,�x����>�2F��7b��˽5^#���>�a�>ʦ�=G���We��w�K��	k�=jw�>�u>��]��ُ�I-�4I�=k9$?l�������$>3��>�@?S�Q?��>��&?,?��>�ڼ>�>�=���>(e&?*��>���>ꎋ>/t>������Q=�V�<�PH��@�KZ.����<�b��RI�<��n;d3>�N�=�v =a!>>�!>&ὺ|Bp��L}=z�>�Zh?�')?�]�>{W�V�V�Y"]��P�﫠=�ڹ�[?���>��?��>���>�d:>��ݼʞ�x?���>���=��k���Y�fȣ>�~)?8�>�o\?��E?��н;�Ͼ��I>�J>.x>�?�J5?���>��!>�&�=����lӿ�$���!��킽J�)�;��<���M�Q-�7��-�����j��<4�\>:�>$�p>�E>�>V<3>vR�>|IG>Qӄ=��=`3�;��;��E�5�M=x��%G<M�P�����Ƽ����>�� �I��>�%9��8ټ T�>D35?X�z�1�þF=��H��� ��DT=�c:>�Z�>|.>H������7U���^�E�Ծ��?�֌?��/?;���S>3mx>M>��D>�I>*�>��I;��%���|�=��>�E:?`0�=�����	]���Y,� �j>� ��х��X�?�rD?�3���
�h�#��gU��??�ó��q	/�,��\%��`3�ÊY��18���8�����s@=�I�>�͞?l�����Y=mɾF[���g�҂��( >�>d��>�<{>�����r���:��Ey��^?޽ȕ�<
�>�M<�EK>/��>͎K?j^?�?g�>��?D��>&3�>�y?��?��#?Y�?�>�>�і=d����bl�<��t��zqZ��w.=�sb>{;
>&P=���=���<0����@a��	���� >�W��Q��1
�<R=?>J��=�?�y?���1�1�>��4'��	�=|qo>���>��>= ],��$�=^��>51?��F?Oh?�%�=B��
ھܾO��=��?�?�m�>�Y��0=z�羡����)>�N�>#����2���F������tZ0���>��>��=��3>�ȁ?N?�S ?��'��'B���w�j�(����=�����>	o�>	�=I�۾D�1��n�"�_�¼4�A��R�%���=��,>�@>��H>̖�=�~�=a=�<�1��� \=ڿ�=�m�>��>��?�s>�&$=�7�����2�I?>�����x�� �Ͼ�d� �>��;>7g��s?���w�}�/
��%=����>Q�?���?�od?�B�o����\>NV>�>1^1<��>��o�X��>;4> �=��x�@5��Wʭ;�\>y>��ɽ�	˾$侾�H�b���|gy��b�<	i���A��Zľmn�Q�4�P���6�� ����ɖ���Q��Eb���{�C����Pƾ�:����5?�L?��(=r".=Y�=����`��/��$��P�����=���g�澆4����5�B�9�z�(�-:�.�t>\?�T��/y�(�5���Z��h�=�7?dݾ_Fܾ�*��6<��=u�P�_7�o����Օ�Vܽ�w`?�96?��̾Hj�o�J�>M.>��?�>Ã >����@��4nt>�,?"�#?y{�Y͈�����/=sx�?�P�?'@?YQ�<!A���������?O.?��>���Bɾ&b�.�?�:?�E�>�-�����vt��V�>��Y?d�K�?�c>X*�>�ޓ>V���h����9���n�8��U5>I�6�Z��_k���<�4d�=p#�>T�u>9[�C������>>�o��+��[r���Ǿ@�`��I �US2>�e���1?k8h<,�+}m�����H룿Y����yA?r|�?��@?�<4?��׾RN$�� 뽅s�>!��>P��=����y�=�~l>Pk�Š#��:�w�����>t��?׾@�M�?͔���CͿ����`ݪ��������=�4�=#$F>�Vͽ��=�q~=���<���& >�S�>O>��>X%G>m-:>eqN>������(��^���|���!J���-�����������W����G���վ�Ҿ�������dQL��7�]z �A�M� ŝ����=Em�>� �>�И>g�$>��C>��^��� �y�������[��j쾩Eݾ����uY�h���I`�| p�F�B����F��>��_=�PL� �?�ͼ�ԝ�=X�>φ�=�n
>J|�>���=��!>�]9>B'>�=�� >w,&>���>�u�>ō�8����)�G����Ͽ�Ǐ_?����Bv��N�B�2n��A�>���>l�=vqW����$%���>��<AV<�����<><��>�;�>h�=-.�w᷽����^+7�Gt�=���>O�U>?�>"r�_
�P�g�閸>�/پ|��=Łi>�{$?�6o?�X2?��=E��>�M>��>,��=x�`>�h>h�>��?]�7?��)?�3�>���=g�O��IK=�iT=�qN��н��ǽ.��Ti���2�<%A��W�=��Z<�N<'W=���<�Gj�y���p=�??1UH?��>���>�x���1n�.L��.�����>���=�>ZB?=��>v �>�
|>VK)��Vc����.���k��>�7>��=����b��ξ>�˸=
um?��>�+�������;�Pj�oN?��"?��1?�U>Le���¾��Կ�ʳ����[R��G)���輫/>�y���D�ؾ���.���k �����=W��>V��>L�	?ܒ�>��N>��>�Z�>}->}rM=�]�=�х<���=��R��e=�{�<�k�;0V��[�=��,=(5��q���>�q Z�=�仚�_��"<?��/?ܖҾ���>�Y����I�?�J�Cq�>ҽL>�
�>Ǥ=>�Ҽk-þC��.k9�m���6w�>�;m?�?�p(�ҷ�=C:����=�^+>Y��oH�>o�\�nv�=�me��j>՚&?H��?z�>�ǂ��L���Sw��e�oy�>i�=�˴�v��?V�P?������W�*_�9���z�о��>O㈾����}p3���8�K�����[�D=O��ꕾhŨ>v}
?��?�q�=8p�$���}���7�� ����4�>�j
?�G��s��^�	���f��_&��d����>%G�>B>�4>�>zF?UEU?�vE?B�,?pr�>��->�t��H??���>H-?�_	?.?��=���=%���P6(>y�7�_z`���n�ѻ� �;�=K��=����sZ=Q��Ţ��c� �x)t=B�=�u�<N��:��=���=��='�(?��D?S���C��)�=�%.�[�1>�?Q�>m�Z>�K=(��>4jH=��>G�?Lk�>
|�5����J�f���V9�$�6?ks@?���>cj>=>/žC^��F�=�^�>�\�:�jt��LѾެ��-���>���>���>��>�?�?�=?U��VR��le�S� �s��=�l=f�>���>:J@>�$��2B�1��D�_�0���G��tB��f�<>�d=�7>hc�=B"�<��s<S�'=A�潤�l=<��=��q>Mn�>_5?2p>���<�㾒��S?��$;w�����+�޽���k,��["��P����>����晿F����Ӈ��zŽ"f�?s�?m�?�^%��V�#<sD�<�n�>M9d�+m���-�>�fI>�mC�� ���� ���:X@U=Zۉ=O�
?�p˼!���]о���=m���P�ֻ�q���oϾ󞗾ԑ�ON7���'��/�������6����Ͻ(E�����{t�nͯ�.Z�7L�?�O?�a>�Z�=�#S�B����߾�qq������<Ә�Ƽ;�״Ǿ�%ľ�PӾ�# �s�5��%����肛>��Y��,��H�|�]�(������?>��.?�ƾ��W���rj=%>5��<$�������-�ccW?��9?��y����߽'�>\"?�*�>e�">�_��
���m�>,_4?�M-?����(���M��=�?���?;�??�NM�keA����a��/?]�?m��>����\̾x��k1?�/:?i��>. �9u���T����>@E[?�"O�Y`>��>�m�>,��$A��s�5��w��!ч�Ն9>�ݻ��� g�1:<�H��=�U�>�Ww>r_�����8	�>����M1���M����y||��蜾�(�>z����2�>�Y�=�c���D���������"Yн��(?ȣ�?e�Z?�!?{����ؾw�����n>\"?6��=\y�=�Aպ	�t>��\>���5�k�������?�&�?���?q��?�����Ϳ�
��=f��� ��_1�=���=F>Z�����=��P=T+ =h[�B�>��>�>}�z>�2B>�&M>�]G>�u���&�t������aG�r*�Y���i���^�s���Gb���㿾�4��韇���L�F��jM�<"����"4>��>���>�Ƃ>6�=�0>>D�L���!Ns���1L�4���J�}
���Ӿ��e�[^�U�j��gQ������?
Z���s"<���>B���?C�=�?�>�-c=�3�=��>%F>�K>��b>X]3>��=�\>;`�=�>�">V�~������r'���-��q��o?/�&���ܾ�S:�g����d���>��?��>>�HL�Ye���l���Ӛ>��y�)ኾl���B>Oح>��>	<h��w��U�;e��H�=� h>�k> *�=
�f�u���v�h��>�\Ͼ�����"�>��A?��t?�mB?ƌq���>%�F=��>�ݶ=��u>�Ҁ>R�:>�r?٘7??P?Y��>���=��z��+��>�%=ZH��ʤ�*�����(�����68=mb@<�4�=���=��\=�ax=�}�=yp�dL<�@Ǽ�9?�5?��>�[�>K����C��TD�,�9>��B>���<�ݜ>�~!?3 �>��>u��>�!�S�������$N�*��>ɶy>�Q�᜗��/>oè>�y3<_s�?�1?J�V�(�F�N>�>��'?�9?# G?��(>�b��4��Tj���տ�����4)��Ƞ<��Y=�I����� p�R���2�W` =]�>��>C�>e_>E>n_�>���>���<��=5�=�%����<Z����/��K��<�9>����>g�=6�&��4�E���y_���;T�=<j
?˗ ?���[]>Q��C�E��+����>��h��?rJ>�_��e�H�^	i��M�W����?�O?`�>����F�<2C���0>�g�>�'>�@�>�E>�Z��X���3�E>�~�>��1?#J�>3�=�Ր�\S���)4��E�>j�<���o�?��t??J>�dL�n��}l3�V
.�=D�>k�[�#뽾�,��+�<�q[����S��
u��>l?��?,Zž�?���P�)=���c��"�;���=Qۗ�ˣ�>����F�f� 4`�V��}����=bg�>�U�=Dߋ>��>m��>O�s?sNB?��H?�q��7�?���7�=?�>�.?jYC?���> ��>�	k>��K��v��y"���{�!���5�=�$O=?�=n_{>�ؽ�o=�"���=S>�J#����̾=NѼ=Ta>�ʂ<)�=8�G>�?;�)?���V�ξ��\>��2ʽ��>�'�>gJ���3�*�~>�Č>m]�>��7?�4�>꘺�j�$�uA���v���~.:?Ae1?�V�>¦=SI>�K-��S���>��>Җ3�F�&��
��ϟ��r/�\'�>��>��D>�l>�x?Jm;?�(?��%�G�3��g����=I���̙����>RϘ>X�(=X:��.�Er���`���)������D$�03<?>]c�=�>��=���=W� =-��<��ýH}���:i=��>�
�>Nw?ǏS>ٟ�<�ۙ��n��D?��L��EvǾ��վ���ݱ8��(�=d>#=�J?���Y���@��VZ���=�z�?fS�?���?P��%+	�w>�>�ɦ>�do��q��n�=B��Έ�=<��=�<����}��)ؽ%�L>�`>*�N�'�8�]\����|N�����G#��o�i����[|h���X�jb�,�@�Y~>�b�F��1/�J��S�/<��9��<p�xga�;��؟?��N?���>@1>SsM�l� �D��b��=Xɹ��/>��	���i�%�4�y����߾��R��/�@z�*j�>�Z�P6����|���(�xŎ���?>/?�Gƾ]�������h=<�%>�<(�͙��?���j�
�soW?�9?�u����#a��!>��?�q�>��%>����N��Α>/64?��-?��1��42�������d�?d��?��??<�O�ǢA������?3�?k"�>�Ǌ��;���A!?��9?
��>5� e���K����>v[?qPN��2b>���>��>���@~�� &��@���m��B�9>�-�
��Th�z>����=Z�>�Xx>�Z]�	��CR�>i���#�F��h(�?����j��k�?����c�>fL�=�$���Vb��莿� ��F&Ͻ��D?�q�?��B?��9?Tm��qn��ym��z�=e�>���>c�>�5>�0>]�8>v1	��NN�������+?��?�V @_?ဿ�Kܿq��ndx�M꽾e��=e�>�Ђ>��׽P�>6�<s��<T�=�!I>0�>�"�>ˉ�>�g>(54>�Ȉ>�}����$��_��A�����:��z�Y��\q~����%@_�Ch�X�Ծ�dþƽ`<�<��.<����	�<��=R���s>�3?ZE�>�p�>z�E>��=>,���z��`�t�S������Wg�����=ž~��xd/�bgp���������:��_^?���<�c�=���>��� >��>�ug=��+>614>R
>ȘY>�x4>m�G>">h�K>Q��=�֥>��r><ɂ�!������Q�K���b?X۾�.ɾJ.��kP��~���u�=�i?��d��^��R���ǐ����>xhj�2�h<��-�>��>�p�>�"�=��=�%,<�e4��%��	<쀰>�B�>���>$�6��l��;"�w�>���P�>�i�>)?j?MJ7?�7d��r>V)�(��>��>�T(>D��>��j>c�>���>�k?j��>A">3�X�C����^���/���	���!�~~%������Q=�(d<yq`=��/=���;�s�=�}�;P��?Z�@�0�US�>�;?��>�q�>^<r��=��@X��$��9͂=/����y�><�>7��>��>4{�>_cʺ΅�K�¾����>�9>��Y�?ɋ�|R=R��>Λg>c�g?�u?����(�ެ,=��=,��>�0?��+?��z>��=����`��Ϳ�����6���缂�[<���=��
�7ཽ�������=g�>P*�>jT�>��B>��#>�,�>\1�>|5>����+��=iXļ��^�����͠>���<�)�=�]�=���<A��<����*� ���T���
��O��W?�*?_�����= ����+��ǹ�B�>�d`>�F?w?�>>Օ=�t'��y�fMV��4���?o5N?��>Us��z�=I��=N�I=%�>��H>mR"=a�������Nj�I
�dH?]�.?}bs;��0�Ʌ�.�~���X����>;��w��:�?S�W?bB��l���z0��2U�>��}�>{��U�Ⱦ���H<$���g�&�
�@�c^߽3C�>{��>�^�?��?�zh4>Ꝿ*��������_5�Jf=�X��W?���>(&�WP�πg�}�����$�羗>�L>Җ�=�Y >n{�>��>�MR?F'A?��?�`���>�dL���1?2O�>!,?w�<?'� ?�M5>�۬�X��c��<�ϽT�T��<��=�_;=��b>�|�=��ּy�=��Y���	>4*�\�p=��=��P�[��=�i�=6�z>�@�>.�	?�5'?4���x��8>� �ߋ;F�_>6C=.��� ����N>�">0��>��+?P�>R����2 ���-�/�����<�9C?V�V?�3�>#�D=��>k�
��6h�i�b><l>I�#��Z$�>)z�b	��v�ν��>HT�>ar�>-�z>��?I�?��.?fCt��SY�f�f�+xP�j ����=�;�y�>�=ƐG���X�~���I�5���@��Hs�ݜ4��r�;8>9@,�6c=F*�>�KD<V>�1A<b���-���|X�=���>��>�E?���f������j�4��na?9a�<��H��)���'����f��.(?B�>��?���{�������^1��q<^�?��?���?�.��V�r�s"y>	/���q>�R�=#�	��N�>����mڼ�=�C���D�<��=վ=��Z>C�T���rϾxq(�ӻ�
��Ke����lоV�k��~����/��nR���$>�v��'��B��pip�
�=��<�$f^�n���,.=���?++?	��>d��~�Q��p���}x�=!�M����>zqD��~]�Z����վ�x�-������l�ƛ>GY��5����|���(�M���X�>>!/?xƾaʹ�ѩ���h=YU%>a��<�_��������K��"W?k�9?�<�#��[Z�h�>��?(H�>��&>�P����K�>�24?w�-?�o�v����-�� �rZ�?6��?8�=?�V\�iA��� �+����z?�
?u�>�e��w�Ҿu$���N?hE6?S�>[����-�������>FU?i<J��)o>Ԏ�>گ{>2��cI����$�����t��U+S>���p��*�B�ր!��%�=�J�>Lr>�`��þ:%�>5D޾^/�J�8�և�ŘQ�Q�
� �>���G/�= j+>RF=KC��H��H턿�����RO?zl�?��D?�@7?6�����������D?>w3�>ŉ�>�',>���&�H>B��>�]龄Em�C���zi?zC�?�?�+Y?L!w�O�̿kL��Ϣ�v:��]	�=y])>+�?>7A�u�=l�D>�Ͽ<��nfB>�Z�>�[2>�_>�4j>ז>�>6���fU"�U瞿1ٔ���O�}C��(�*���0��ߎ�n�Rc��Jr����9�C
F�*����1�ǡ��\��4�>�s?l��>�7�>�D>`�(>�倾����m4n����C�B���� ���̾區��X/�W�i�D᏾�� ���?s��<���=�"�>���> ͚>���=9�+>�;>W>%E>;�8>D/M>�9+>ScW>���=��>��=�(�6�g�$Rᾝň�9����>۸�jkƾ��[�
�P���ya�><�Q?h{
?7dA�@��-	t���>0�ͽ�>���Q��Q��K_>�2�>��Q�jG��ѽ�W�7�>��=�	?7p�>����8��,���^�>���>�_Ծ�b�=�\v>�p(?��v?P6?	 �=��>aX^>�{�>	"�=��N>�zP>���>��?�+9?<1?&q�>&׾=��a���
=�l5=�m?�|�W��b��R|���="��,�<β-���Q=��o=���;`�d=�OI=x˼�g�;���<Rl?�e-?e=�> ?`��2�[�.�M�B]�Jݲ<U3�wq>N��>r?�?B�?2��>�qŽ:�Ծ:\��r8�>�lM>sR�֥/�ݨ���F<�H?�<R?�G6?���=fRP���n>\r�>}��>�	?�Q�>.^>���'O���Ϳ���h5�qup�^��=�<����nb��<�`���oK��;E>|��>�?�>�P>�>l
>jي>��>���<�"�=�>�G�=9ѹ:3��7���?�V����O�Ke�oL`=
X�<e��=%��e��;���=�??�V�>X����ؽfkƾK8���?���2?1&?kgJ?t�?���>�"#�8�]�i��ѭ��Y�>��b?m@'?�����f(>���;�o�>5��>�Z���(>p�*��q�o��<z�7?�}S?��>3۽�����Z ���>�= ����S�?�^?J�_�ϒU���#�t:���%�,d>�\����;����I�/"�F渾�0;��ۻ���=�:?���?-�*��wd=�ޕ�GV��o=��p�o����[��x��>��&���f��J���I��rQ�FT�>�,>K� ��@?�u?�;�>�"4?̜4?#D5?:g<�I2?�
f���M?,]�>]�?��>xG�X�V��n�=q���x�>� �I���gԅ=�E,<�����R0>�d>����8�=S�	=�X�<n1��P;�=%�Y=�8y�V�=���=�:�=�zO=Ю?��?�����>X=<f��7��9��L��5�_ӎ�t�׾d���>5'1?(iP?)��>��)������iz��`N�<���>L�V?��>�û�!�>;�¾�r�<���>���>�����ӈ�����$�žO�W��?���>}�*��"x>��?�`-?Y�?���<�p���`�7���}�K��<{��>��>Z��=�P�[1�'x��b��m>��p���u��I�=�?>�Ӏ>�q�>�)F>��E>R��;�f�<�����(>s����>�`�>��?$2M>�">�%���G��(�D?�# �����%=B��W˯��콖�w>��F��h�>3Ӿ}w���f���N��w�>`M�?���?ր�?�d�47=,�9>X���Y�B��H>�>�����&>�%�>��=�{��	�<�h�=8�/>�:U>vRQ��ݾ��Ӿ��A�쀲��}�-*S�N�������2�)t��Ba����RPϽe�р7��f�=�rJ�D����W5��w�&b��"ʣ?�D9?z��>C׃=G�e���:� �Q��>:G��.4�=���L�����qL�l����P��#��6��B�1�>�W��ᑿ��z��&&��¼�0>،+?�ʾ������V�o=,�#>nn=İ�1���Aɚ�V'��X?��8?��N�����½�>�?NP�>ZW*>)捾`r�ʫ�>s4?�.?�$�u�������6��N�?���?Q�M?���g�F�V�<��ּK��>P �>�I,?�\,�0R�����|K?�+?_�U>���fW��ܓb�/�>��?�ƭ�y�>m��>�=�>|�(�׎����m�i���"��Z,|�>c�LM��}����M�����>;#�>�f�=�j������\�>��dD5�Pq-�CM��Y���_��#^�>�8��1_>�,>\:.�N�����$V��k�m�4�N?M�?�kF?�|9?��̾� ���ν�<=>kk�>��@>U>�4 ���)>�]�>SD�._q��B�$C?dQ�?	z�?o�Q?&�=Gӿ�� ��������=%�=��>>��޽�ɭ=�K=uȘ�%Z=�t�>~��>o>?;x>w�T>ћ<>��.>q�����#��ʤ�3ْ��[B�� ���wg��{	��y�����ȴ���K�������9Г�x�G�`���T>��m׾*I>gr'?���>���>V�E>��<>��n��Ʊ�su��|�*��~Eྣ2Ҿf�˾�������Y8 �D��ꕼ� 	�+�?db>���;Z'�>[tP�k�>q��>-��<mZ	=�Г>�b�=��$>G�b>*h�>4DX>>J>��->3��> ���p��Pd����b]]�n����"?a,���8龋�?�i�׾`=M�E�>|>8?��>W�.�u؍���H�[2�>����hQo�9?=�|�󽾠�>�3�>�|�<m��e���X�=��Za��)�>�?m$�>*L���߾ >�����>���>�վz�='Iv>]�(?�w?�D6?{�=��> wa>�W�>�w�=��L>�zP>�P�>_�?�9?i�1?p�>��=��`�_�=�9=L�>���V��I��1�9Z(�@S�<tB3�_DH=�u=�	<�`=D�A= Mȼ@��;͑ =n�>t�?%��>�;?記���K��J�C���6>F*�;n>��>���>��>d� ?<��>.�z>}��I7߾�%�>�1>�nR�<���*5���>��>�Wl?_!Q?��=:n>�@%��x�����>y"d>�w?��>;�>��e��U��&ֿK��U�*�����s�J��<�&������P����V�p>wł>o�>��f>#�>r�=�<�>�8�>dZ5>�%V=��F=8�ؼ�"�j���i�=�Հ����<�K���`�h�o�xĽ�˲���5�Mc��2�Ѽ�x<%�B?���>����
��\��.�����[�D�P?RY?�_ ?��?�N�>���QF�E�Nq@��E�>R�?�[?Y���S�=�瘽�9:�q��>,��>��z=��_ۤ��,l��+>M�	?W'?XmQ>
;i��e��	{�����G}�>'���x��Ac�?�Da?��J��ꖾ���l�3�W���\>�!���,4�p^��*��/�����;i�"9D���{>�?�?�[��~�
=��{�h��m��H��&KR��`<ߡ�>�nս�sѾ��s�����
Y�I��>�ģ>Ƒ&��T??���>暦=��W?�U?�{O?�`K��2?�g��6B?:��>�?��>�n2=h���B>|V>���Q��CJо�q�=�D���ۖ����=���=@�ŽKli=*�<�t�ü�M[�1�YBb=.U=�#=�0�=U�y=v�=#?���>�{��1�>�hF=Dm������N���:��=��>N�>EQ ?��n?,[?lU>��
��� ��G�y��=č?	�T?Z?�ƻ�r�=d��?W��F�>~�G>��[��Ā��$5��߰��8.<=V?N�m<$�$��uu>a�?�0?Cg?�g���7���V�{����Y�=���>e�>ݨ�=,��<:��9z��~]�@�+���۽z���>��>��~>OmY>Z��=�->�X��K�=������V<�y��b�>�[�>ǎ
?�+�>��=�堾oK�c	<?�c��l���T̽I;A_��
�a��>�+-�JA�>�1���r��v	���%�@߭>���?T{�?\�J?�İ��$>�`t=Dy	���p���'=a�=>a��;f	�>dSj>ޭ@��˻<����n+>5N�>�=�>#5R=U�dv���o�����Y���>>�|�?#پ-K��r�|���7����i�ӽݪ�]ʾ�ाPܽ6Y�x恾W��i�y��ך?��Z?���>��_=�q?�����㘾���=�y��|^�<������{䎾���������Z���w(�a�s�ȾJ�>*˂�,��-�t����U���"�<g�?W�� ��mG"�I���|ʐ>j��>t��&kl���c��m_?}3?�ZܾU�*Խ� �<u<�>�f�>��>r���_-���L\>�+?K� ?/<�=�s���������Q��?L�?�mS?yb9���K�g�������>�z�>��?���%��g���@!,?��6?f��>�nԾt|y�}8�Π�>Ďg?V�ܾQ�>��>o��>�,i=?$�]�
>��ؾ�ݛ����>3�A� �b���n�ad����=��p=o�k>A����ž`��>y�꾏�N�߅H����	P����<i?���>@�h>�>ɶ(�U
���ˉ��<���L?ꑱ?߄S?gm8?�������7ަ���=C��>զ�>��=���l��>��>��rjr�r���?J�?��?FRZ?Z�m�M�ƿ[ڋ��(��6?վ�/>%�>~�W>�����<%d�=я=��?:�b>�Cd>9P�=5}!>��=�T�>�̆>s���p�RM��a��1@�<����5�h�+��(��O�����E����"�1�U�ؕk��ϻ�]e���F�=p{ܾeQӽi�#?7��>pj�>W�>�D�>(��'�7�B^A������[�;_�-��;�'��D@�V�o���⽵G=sE4���?�_�>Ѓν��>ֳ�j1{=���>��;Xr>h��>`ۅ>��>.�=b�>�<�wd>��f�L�>4��=8>��p�}���*�ʖm�n<����J?������%�3��i׾W���l>��?�}>�A#��ݑ��k����>H�Ҽ b�..ֽ� �a�i>>�>�a>M�<dd�y�s��yѽ�B{=��T>��>	�}�E�O���-���J=���>����LW>6N>��2?k$�?��Z?B��<��>e�>��>�0�>N�>ϖl>�xU>��>�V?��L?e�>%>�����=">��ʽ�ׇ���<B�X<3غӹ>g>�<}=[�=l	�CV=���<4j�>_�"��=3�?ԇ?�Q}>wk�>�[��ш+��2]��`	�F��=�p�M�8>��9>�)?l(?��?MD�>}�o�؞�*鮾��>��>n���鍿�}�>>�>PѮ��9w?�#(?�&�#n���g�=S�M>�|.>f<9?=W?l\�D��b������ÿM�;��j>��P�=�>�ȭ>O]�t�����ѽI�9����`�=�(J=��[�Ǆ%�RtV�K��=��>���>Pa�=2�G=�}�<��E�ݖs>��=��T;����0��ϽK���[��=��3��cB��e�<O���,j��G����?��?HT�e�=����ݠ���	��p��>�?x0?�"?�6^>6!�~�N�UQF��������>��c?���>�FO��H>�2�@I`���>hE�>
f<�G>��$�X����0>V�>��/?2�>�*��5^�KVl�K�����>Ǣ<G齾��?ȅ?��B��m���eؾ��Z��C��Z�p����������L��$4)�dα������e���@�=�*?9�?W{���y�=�������'Ɂ��ꆾ�>L>)��=�(�>�<8;��ټ�mE�i���W=�L�"=�S>��v>��>���>7��>!��>ͯq?�o�>E�>j7=�?w��>�!?�4?��>z]?��>#�v=�U�>i^>+䪾��C�{�$�^>K�<�7Y=�eA>�ƃ>�����<׺l�[S�=��;��=��ʢ�
Pݽ�2>�v&>�29>e�>�Q?*(=?L��}8ֽ�5�=�:���ƾ�Ǭ>v3�>.xl��S�����؛�<#_�>y�c?��?�:�>%-"��‾.ӷ�S�Y=�j?��$?�>	�=�ֽ>]��C���c��>�C>[������B��I� �򍾉��>lP�>&�=bh>�r~?��A?�^"?4���ݙ.�7Gv�+������&� �>�(�>Y;�=��۾�6��s��`�ԯ0��AG�X�E��R�<l�=*�>U�@>ݵ=��>�[=�����ؽPZG<i\��"�>i?�>�?�Y>�Ƈ=/䪾 ���?E?L�������VtӾ�	[���>�>�u���> ��'��l.��=�7����>���?�w�?��`?>9����+�\>��l>�$>�=1�:�WYƻ�z��չ
>��=(މ��E���3<-�A>%�h>E����Ѿϑ˾�3��mÿ�T��EL�c��4����Zžk��� Y��K����ɽv�ɾX�V��fa��*8��0F��x~�D���
j�^M���}?�vd?(�=�0Q��(�(����̾�� >D���OlW�a��3~?�@0��	Ỿˮ��l�p'��]&�r������>�I[�s-��H8}��<(�ݽ���d@>�.?��Ǿ���3-�f8e=;%>'�<uN�p����Κ����&�W?�?8?�������E�X�>�?5I�>$�&>�m��:��3'�>m3?�h,?QX��֎�LG���ۤ�rǻ?���?XkL?2�ϽݓK������{X�>x]�>�W
?�
W��o��C�<��>-�6?���>	�𾩓�� �A5�>�t�>�yG�a�0>U�>fN_>5�z=%ᅾ��,Dy�1C��>)�6�|N����Bɬ�jB?>�ɕ>f��>Z�m��l�f��>�EAS�`�K�$.�/�LG=ha?��w�>�}t>6�>W*�{������5����Q?�,�?��U?R6?���Q�`���c�=<��>Fx�>�@�=�x�G-�>���>r9ܾ;6m�>��
?u
�?��?��P?i�o��}ǿU������4��w½���<y�Z>;jȽ�>u-l>C�d>���/�	>Y�U>́>��X>A�>Jp�>ɠ>s���$����q���Q� � ��T��?��G���� �߹ʾ�T��99�?���M��Q�r��=UI�=�k���G�>t��>(Q?�>�.�>�X���e�����~�+�s��^��3o���ݾJ��Pzp�`	����A�@�N=���n��>��#>�M>�q��>|���(�<Q��>þ>h�O>|��>Fd>�a�>��=[��=T�=a>�>�*�>J�>���y��� ���]��y�R?��o�[3���9�ע��}m/��d�>�?&*>��.�]W��] v����>�"@��fY��^��d,�<�@�>ί�>���=~@�<�G����PA0����<�lv>ۚ>t�=3�[�ϗ2�4����>9�ܾ=L�j>��'?S�w?p�5?Z!�=�>�Vg>b?�>:0�=К6>#4<>�|>��?
9?E�2?4�>p�=c�`�sM4=�t=@-B��X/���Ƚ���=��ǧ�;�+�r{a=E��=��<�V=A9=ׁͼ�K|�2�<�`?N;?�<k>�>�.��P+k��O��+*<�ࡶ��q��S��<�]>JQ?-�F?y+?*��>xǹ�)�������̼>�ͦ>3�~������p�>�82>Nr�=~?H��>�4���7���j>Xx�>9�{>��5?nR?,���ғý��B�=�w���O�5E��(�����=t�D>�6<��۾:��<>���=��B�O���sY����Y��=�l?SM$?�)�>�6�>���=�R>igb>A�X>�K>���=B0	�5㽉�+��\5����Zɽ/��D<�����2���4��(�K9?G?� <Ӽ�nP�h�������>�d�>�u�>�C�>Yn=�!��"[�[w;� ?�98�>�I?�V�>��I�m�=��8=�O�bG�>�ܫ>�A>�Ĩ���O��Z����=���>,�?^�>ɪB���m��X���]��a�>��=b_Y��?yˉ?�88��cཉ���{o�����<��ďL�����v�پ��,��q¾/������>)�?��?9ؽ!�g�=��kl��|�؆�O�g��O�;�j�>��Ž��%=�LS��U����?<������=A�>�j;>ߕ�>��\?	}+?�Qa?@�?/�!?8J3�3�?}�0>7�	?K<?JN�>���>Q��>��=��=�]�;�[�+:��8���>�L�=p��>�f?>� !�����>.>��p=�A=3�<M�L=Ͷ^=K!s�F[�<�~a>�-�>{�(?�@?����K�~Q�>~=p�4_�< ��>�J,>f�2���پEw#����>:�>�(:?5��>ҵ齱�
�Yh.��\Ҿm�܌?Yu.?\�_>P>���>��;u�:>i��>f��>�I�������J�XBӽ��
?���>n����>z>_Y~?��A?cd?w!���q+��6i���$�Z�k�J��;���>Tx�>�ڵ=6cܾ�3�3qs�(�_��1�Hd��(3��}�<&�=�J>;.>7o�=��>���<�@�����Q�_<�&c��t�>��>gR?j F>��=}���� ���G?+NJ����|���߾�5�n�>?1p>�h��G�>l�Ǆ�7���Ǆ6�!��>��?X��?+8[?�O�
��c�G>�Ɣ>�aP>m�F�@�6O	=��9��Dl>x�S>l�սrꂾ[�$�	>��_=�Ô�{�`V�%�H�����C+d����
����a��P�4������#���i���s�������"��� ���_��7���̢��O�����?<XL?��=�_�=Y�Q��� ����'=om��S��������	u��:��2h��NϾ�����6�K
����>j�Y��B����|���(�%B��6�?>�4/?Pƾ ���j���g=�P%>��<�8ﾊ������ �
��gW?V�9?�P��;���὾�>��?!x�>��%>K��GP��	�>{34?5�-?����6���Γ��m�?���?GC?��&��O@��Q�0������>�?���>yń�y�žx	���?A~@?��>!���(ȅ��^��>o�I?�eP���U>M��>>I�>�}��b����Zt�-I���Y��*>'\	�S+1�i�s��Z!�ɸ�=��>uw>�l��࿾`��>y�꾏�N�߅H����	P����<i?���>@�h>�>ɶ(�U
���ˉ��<���L?ꑱ?߄S?gm8?�������7ަ���=C��>զ�>��=���l��>��>��rjr�r���?J�?��?FRZ?Z�m�M�ƿ[ڋ��(��6?վ�/>%�>~�W>�����<%d�=я=��?:�b>�Cd>9P�=5}!>��=�T�>�̆>s���p�RM��a��1@�<����5�h�+��(��O�����E����"�1�U�ؕk��ϻ�]e���F�=p{ܾeQӽi�#?7��>pj�>W�>�D�>(��'�7�B^A������[�;_�-��;�'��D@�V�o���⽵G=sE4���?�_�>Ѓν��>ֳ�j1{=���>��;Xr>h��>`ۅ>��>.�=b�>�<�wd>��f�L�>4��=8>��p�}���*�ʖm�n<����J?������%�3��i׾W���l>��?�}>�A#��ݑ��k����>H�Ҽ b�..ֽ� �a�i>>�>�a>M�<dd�y�s��yѽ�B{=��T>��>	�}�E�O���-���J=���>����LW>6N>��2?k$�?��Z?B��<��>e�>��>�0�>N�>ϖl>�xU>��>�V?��L?e�>%>�����=">��ʽ�ׇ���<B�X<3غӹ>g>�<}=[�=l	�CV=���<4j�>_�"��=3�?ԇ?�Q}>wk�>�[��ш+��2]��`	�F��=�p�M�8>��9>�)?l(?��?MD�>}�o�؞�*鮾��>��>n���鍿�}�>>�>PѮ��9w?�#(?�&�#n���g�=S�M>�|.>f<9?=W?l\�D��b������ÿM�;��j>��P�=�>�ȭ>O]�t�����ѽI�9����`�=�(J=��[�Ǆ%�RtV�K��=��>���>Pa�=2�G=�}�<��E�ݖs>��=��T;����0��ϽK���[��=��3��cB��e�<O���,j��G����?��?HT�e�=����ݠ���	��p��>�?x0?�"?�6^>6!�~�N�UQF��������>��c?���>�FO��H>�2�@I`���>hE�>
f<�G>��$�X����0>V�>��/?2�>�*��5^�KVl�K�����>Ǣ<G齾��?ȅ?��B��m���eؾ��Z��C��Z�p����������L��$4)�dα������e���@�=�*?9�?W{���y�=�������'Ɂ��ꆾ�>L>)��=�(�>�<8;��ټ�mE�i���W=�L�"=�S>��v>��>���>7��>!��>ͯq?�o�>E�>j7=�?w��>�!?�4?��>z]?��>#�v=�U�>i^>+䪾��C�{�$�^>K�<�7Y=�eA>�ƃ>�����<׺l�[S�=��;��=��ʢ�
Pݽ�2>�v&>�29>e�>�Q?*(=?L��}8ֽ�5�=�:���ƾ�Ǭ>v3�>.xl��S�����؛�<#_�>y�c?��?�:�>%-"��‾.ӷ�S�Y=�j?��$?�>	�=�ֽ>]��C���c��>�C>[������B��I� �򍾉��>lP�>&�=bh>�r~?��A?�^"?4���ݙ.�7Gv�+������&� �>�(�>Y;�=��۾�6��s��`�ԯ0��AG�X�E��R�<l�=*�>U�@>ݵ=��>�[=�����ؽPZG<i\��"�>i?�>�?�Y>�Ƈ=/䪾 ���?E?L�������VtӾ�	[���>�>�u���> ��'��l.��=�7����>���?�w�?��`?>9����+�\>��l>�$>�=1�:�WYƻ�z��չ
>��=(މ��E���3<-�A>%�h>E����Ѿϑ˾�3��mÿ�T��EL�c��4����Zžk��� Y��K����ɽv�ɾX�V��fa��*8��0F��x~�D���
j�^M���}?�vd?(�=�0Q��(�(����̾�� >D���OlW�a��3~?�@0��	Ỿˮ��l�p'��]&�r������>�I[�s-��H8}��<(�ݽ���d@>�.?��Ǿ���3-�f8e=;%>'�<uN�p����Κ����&�W?�?8?�������E�X�>�?5I�>$�&>�m��:��3'�>m3?�h,?QX��֎�LG���ۤ�rǻ?���?XkL?2�ϽݓK������{X�>x]�>�W
?�
W��o��C�<��>-�6?���>	�𾩓�� �A5�>�t�>�yG�a�0>U�>fN_>5�z=%ᅾ��,Dy�1C��>)�6�|N����Bɬ�jB?>�ɕ>f��>Z�m��l�f��>�EAS�`�K�$.�/�LG=ha?��w�>�}t>6�>W*�{������5����Q?�,�?��U?R6?���Q�`���c�=<��>Fx�>�@�=�x�G-�>���>r9ܾ;6m�>��
?u
�?��?��P?i�o��}ǿU������4��w½���<y�Z>;jȽ�>u-l>C�d>���/�	>Y�U>́>��X>A�>Jp�>ɠ>s���$����q���Q� � ��T��?��G���� �߹ʾ�T��99�?���M��Q�r��=UI�=�k���G�>t��>(Q?�>�.�>�X���e�����~�+�s��^��3o���ݾJ��Pzp�`	����A�@�N=���n��>��#>�M>�q��>|���(�<Q��>þ>h�O>|��>Fd>�a�>��=[��=T�=a>�>�*�>J�>���y��� ���]��y�R?��o�[3���9�ע��}m/��d�>�?&*>��.�]W��] v����>�"@��fY��^��d,�<�@�>ί�>���=~@�<�G����PA0����<�lv>ۚ>t�=3�[�ϗ2�4����>9�ܾ=L�j>��'?S�w?p�5?Z!�=�>�Vg>b?�>:0�=К6>#4<>�|>��?
9?E�2?4�>p�=c�`�sM4=�t=@-B��X/���Ƚ���=��ǧ�;�+�r{a=E��=��<�V=A9=ׁͼ�K|�2�<�`?N;?�<k>�>�.��P+k��O��+*<�ࡶ��q��S��<�]>JQ?-�F?y+?*��>xǹ�)�������̼>�ͦ>3�~������p�>�82>Nr�=~?H��>�4���7���j>Xx�>9�{>��5?nR?,���ғý��B�=�w���O�5E��(�����=t�D>�6<��۾:��<>���=��B�O���sY����Y��=�l?SM$?�)�>�6�>���=�R>igb>A�X>�K>���=B0	�5㽉�+��\5����Zɽ/��D<�����2���4��(�K9?G?� <Ӽ�nP�h�������>�d�>�u�>�C�>Yn=�!��"[�[w;� ?�98�>�I?�V�>��I�m�=��8=�O�bG�>�ܫ>�A>�Ĩ���O��Z����=���>,�?^�>ɪB���m��X���]��a�>��=b_Y��?yˉ?�88��cཉ���{o�����<��ďL�����v�پ��,��q¾/������>)�?��?9ؽ!�g�=��kl��|�؆�O�g��O�;�j�>��Ž��%=�LS��U����?<������=A�>�j;>ߕ�>��\?	}+?�Qa?@�?/�!?8J3�3�?}�0>7�	?K<?JN�>���>Q��>��=��=�]�;�[�+:��8���>�L�=p��>�f?>� !�����>.>��p=�A=3�<M�L=Ͷ^=K!s�F[�<�~a>�-�>{�(?�@?����K�~Q�>~=p�4_�< ��>�J,>f�2���پEw#����>:�>�(:?5��>ҵ齱�
�Yh.��\Ҿm�܌?Yu.?\�_>P>���>��;u�:>i��>f��>�I�������J�XBӽ��
?���>n����>z>_Y~?��A?cd?w!���q+��6i���$�Z�k�J��;���>Tx�>�ڵ=6cܾ�3�3qs�(�_��1�Hd��(3��}�<&�=�J>;.>7o�=��>���<�@�����Q�_<�&c��t�>��>gR?j F>��=}���� ���G?+NJ����|���߾�5�n�>?1p>�h��G�>l�Ǆ�7���Ǆ6�!��>��?X��?+8[?�O�
��c�G>�Ɣ>�aP>m�F�@�6O	=��9��Dl>x�S>l�սrꂾ[�$�	>��_=�Ô�{�`V�%�H�����C+d����
����a��P�4������#���i���s�������"��� ���_��7���̢��O�����?<XL?��=�_�=Y�Q��� ����'=om��S��������	u��:��2h��NϾ�����6�K
����>j�Y��B����|���(�%B��6�?>�4/?Pƾ ���j���g=�P%>��<�8ﾊ������ �
��gW?V�9?�P��;���὾�>��?!x�>��%>K��GP��	�>{34?5�-?����6���Γ��m�?���?GC?��&��O@��Q�0������>�?���>yń�y�žx	���?A~@?��>!���(ȅ��^��>o�I?�eP���U>M��>>I�>�}��b����Zt�-I���Y��*>'\	�S+1�i�s��Z!�ɸ�=��>uw>�l��࿾f��>�EAS�`�K�$.�/�LG=ha?��w�>�}t>6�>W*�{������5����Q?�,�?��U?R6?���Q�`���c�=<��>Fx�>�@�=�x�G-�>���>r9ܾ;6m�>��
?u
�?��?��P?i�o��}ǿU������4��w½���<y�Z>;jȽ�>u-l>C�d>���/�	>Y�U>́>��X>A�>Jp�>ɠ>s���$����q���Q� � ��T��?��G���� �߹ʾ�T��99�?���M��Q�r��=UI�=�k���G�>t��>(Q?�>�.�>�X���e�����~�+�s��^��3o���ݾJ��Pzp�`	����A�@�N=���n��>��#>�M>�q��>|���(�<Q��>þ>h�O>|��>Fd>�a�>��=[��=T�=a>�>�*�>J�>���y��� ���]��y�R?��o�[3���9�ע��}m/��d�>�?&*>��.�]W��] v����>�"@��fY��^��d,�<�@�>ί�>���=~@�<�G����PA0����<�lv>ۚ>t�=3�[�ϗ2�4����>9�ܾ=L�j>��'?S�w?p�5?Z!�=�>�Vg>b?�>:0�=К6>#4<>�|>��?
9?E�2?4�>p�=c�`�sM4=�t=@-B��X/���Ƚ���=��ǧ�;�+�r{a=E��=��<�V=A9=ׁͼ�K|�2�<�`?N;?�<k>�>�.��P+k��O��+*<�ࡶ��q��S��<�]>JQ?-�F?y+?*��>xǹ�)�������̼>�ͦ>3�~������p�>�82>Nr�=~?H��>�4���7���j>Xx�>9�{>��5?nR?,���ғý��B�=�w���O�5E��(�����=t�D>�6<��۾:��<>���=��B�O���sY����Y��=�l?SM$?�)�>�6�>���=�R>igb>A�X>�K>���=B0	�5㽉�+��\5����Zɽ/��D<�����2���4��(�K9?G?� <Ӽ�nP�h�������>�d�>�u�>�C�>Yn=�!��"[�[w;� ?�98�>�I?�V�>��I�m�=��8=�O�bG�>�ܫ>�A>�Ĩ���O��Z����=���>,�?^�>ɪB���m��X���]��a�>��=b_Y��?yˉ?�88��cཉ���{o�����<��ďL�����v�پ��,��q¾/������>)�?��?9ؽ!�g�=��kl��|�؆�O�g��O�;�j�>��Ž��%=�LS��U����?<������=A�>�j;>ߕ�>��\?	}+?�Qa?@�?/�!?8J3�3�?}�0>7�	?K<?JN�>���>Q��>��=��=�]�;�[�+:��8���>�L�=p��>�f?>� !�����>.>��p=�A=3�<M�L=Ͷ^=K!s�F[�<�~a>�-�>{�(?�@?����K�~Q�>~=p�4_�< ��>�J,>f�2���پEw#����>:�>�(:?5��>ҵ齱�
�Yh.��\Ҿm�܌?Yu.?\�_>P>���>��;u�:>i��>f��>�I�������J�XBӽ��
?���>n����>z>_Y~?��A?cd?w!���q+��6i���$�Z�k�J��;���>Tx�>�ڵ=6cܾ�3�3qs�(�_��1�Hd��(3��}�<&�=�J>;.>7o�=��>���<�@�����Q�_<�&c��t�>��>gR?j F>��=}���� ���G?+NJ����|���߾�5�n�>?1p>�h��G�>l�Ǆ�7���Ǆ6�!��>��?X��?+8[?�O�
��c�G>�Ɣ>�aP>m�F�@�6O	=��9��Dl>x�S>l�սrꂾ[�$�	>��_=�Ô�{�`V�%�H�����C+d����
����a��P�4������#���i���s�������"��� ���_��7���̢��O�����?<XL?��=�_�=Y�Q��� ����'=om��S��������	u��:��2h��NϾ�����6�K
����>j�Y��B����|���(�%B��6�?>�4/?Pƾ ���j���g=�P%>��<�8ﾊ������ �
��gW?V�9?�P��;���὾�>��?!x�>��%>K��GP��	�>{34?5�-?����6���Γ��m�?���?GC?��&��O@��Q�0������>�?���>yń�y�žx	���?A~@?��>!���(ȅ��^��>o�I?�eP���U>M��>>I�>�}��b����Zt�-I���Y��*>'\	�S+1�i�s��Z!�ɸ�=��>uw>�l��࿾�8�>�;��N�ʳG�J0������<*4?��.>�nj>�\>��(��������,��
]L?���?�oS?�h8?#6��B�좩�QH�=S��>��>��=�k���>���>�����q�����?۩�?��?��Y?l�m��ؿ�ʚ��mӾ-����=���=��$>�E��h=�=
�=f<
	�= ��>��=Q�>��>�5>R�>>V̆��d$��S������F�խ�~�	�i������
ݐ��#�>�������|;��0��G�r���@Z���C���ܾ�UI=��>�l�>G��>*��=Y�W>*�����-���R4�����^�����(���F�����V(��c�
Z�� ��#?%��<���;��>�ޏ���=C�>��}>d)�=�>΀>2T=z�>�Ã>/Ǜ>��>��u>l��>X.�>C���.��r�k�CU�֕�f�S?�[��I��m��O�c�����S>S��>pBK�pnN��X��OӒ��*�>T�*=kؾd�oD�=�$~>�)?�P����>&��ٟ�<]/�;O�5>,�+?��>�η>�#
��/�=�r��?���[�G>_�?�H%?�c_?w�W?���>ͩ�>����>��=���=2>~I.?��7?�{^?��=?*T�=:껽��=�+K=��[��c���_=Fa�<\�ػ�=5�ҽh`�(ms��6��>-�=�8����p=���<��>�@?��?wo�>��g��C���D��0��-��=�L!�d�>��?�qB?͍�>7�>�{���I�<$9��\
���>ܲ2>bs��t���;ff�>K]�>�>?=�"?�A�ɮ�oY>}&�=�H�>��>��?=�>
�s>}E�=-s
���ҿh-�����d��t���4c=7�i�}'ۼ���=i;+�0@!�ܣ ��>�#�>J:�>n�>�J1>��>L��>0��=
�>zx�=?4�c�E=yyͽm�c=�
���S�=/}Ž݅�=!�<�҆�R���B����<¡P��=x�G�?R?��'��b��f�;����������>��>CY�>ճ�>,�=�%��hU��vA�wG��E�>
qh?,��>l�8�_��=8�0��PT:�γ>4��>��>�`�2���U���>�<9��>͔?�O�>��V:[��to�c�
��/�>��\�v�is�?�K?c��DQ�nO�/~8�k�K��i�<���	`,�aۆ���c�@�`��N��O����YK=��>�<�?	�G��җ�dؾ�����=����j�	%,=p�>$NE>Yv%=�����Y�� RB��|>�Ք��$��K_�<=!�=��> r?�?��_?Z8?Mk
?7y�����>�p�>�L%?2!	?��>�?��>'"�>�.�>� �=(�=��!�hƮ���;2��=�x= ��<5��=}f=K��=�{=�>�v�|��}\=>=��"=m��= e=�L>�@�>��K?KB��H���^��0rT�wx����-�]�>��=q�׽��=���>��6?�O5?���>�<��ھ�c����ә����??�gY?��#?_�v� ���<���׾]`�<�>$�K>>c������ح��,��>�5�>�[�>OU@>��{?R�_?V�?n��gP� <���l/�*�m�c##<�GX>�T�>x�>��־P�;�.����p�3<���5�*�Ր�<O�K>��="��=.X(>��>�G>�˽�u�$�������>�֠>�/�>�Z�<P}c>��������I?���y�2A����о���x>R�>>>��J?2��O�}� ��+&=�3��>5b�?D��?�Kd?a�B�%���]>6�V>�>R�/<�'>�������� 3>���=��y�����6��;��\>��x>��ǽ�ʾ�PE�2���O�Z�w<�Ͼh��=�¾�&���")�{ɕ�2K�x�ƾ��%��p��#n��(]M���\�q������TB�3	�?pf�?.�>:���������n%>p���z���۟������q��\��3����H���E1�x-F� ����>�yY�AA��(�|���(�L����{?>�3/?�[ƾ�̴�"����g=j%>� �<�6�B���[�����\W?x�9?	O쾆*������>�?{w�>.�%>[$���'��+�>�94?��-?��뼰���6��&����l�?V��?{;?T�*�=h=�K����ֽ"f	?!
?a�>�5���eپUԣ�R�?B�<?��>GX�f��%�����>XS?7�G�3XD>3�>j�>����·O�󝈼����uM(���s> b�<y�����>�>��Ź=[��>�S>�MN��?��b��>�?�_�N���H����d���v�<�?>��1>�i>B>`�(�Y���ω��'�_�L?	��?��S?tk8?^�����ͬ�����=��>"Ӭ>���=\����>���>�h��xr�'�ܘ?�I�?V��?�[Z?��m��dο�	���q��оp�*>_y�=��>z
$>��Ka��P���N���=K�>E<�>�q�>��>
�>�Gv>e����#�qƪ�yь�=�O���n�
no�Q<*��x��5����D���*+�=��=���� �5�"�=���z��=���>('�>MͰ>�i4>��?>�qt��d���|�H���=��:+��e���C�]����l?K�?z��qs��^����>�'X<�:�=��>�m��g,>�˓>Ń�=��>` >��3>X�>��*>V8>��->��+>]�	>:i�>��>��I��(��v�q��^ ��6�yKz? �ǾQ��ӏ��@2��?D�SR3�Ec�=6ɗ�s:v��@���8��F�>,��S��n:�����S�>�B ?���ND->Ru������wf���Z>o�,?3�>�,>��9Nս��ֽR��>y{��A�<X�>�O?-=5?�	L?�(>��"?P��=�l�>z>�V�<��>���>��?�??U?��?F�+>��p����%_�;��]�u�����=��=��S���=*w��҅=�l>G=�Q�=�+���*�۽Q7�;>V?^zB?�?E��>�ܱ��y%��,��?�<>��<�2?V�>�:�>��?�S�>�5�=L����򳾹@����>�>r>J���b��~���h�>_�>�h?��?y����Yݼ��<AZ�=F�i>(q�>�=?E�?3��>N+�>8a뿃����~k�L��x��=g�O��=��I��t�7���2��x��������>���>2�>�ג>W�?��>��>L�>�J�=��!>�4ֽ����i�@�7����=[x�=�=�=潦|���p�c�ӽ�{���%
�,���|?�? G#�����nf�L���$�����>���>���>/��>B��=^Q��;R���>��=B����>&g?���>��6�9��=�D�8qѻ>i�>�V>�q�
M"�?���%��<=��><,?�5�>�a�c�X���n��H��>�U�=q1����?ѿZ?������7��F���T��-�=ھ��k�¾2漨KT�̫m�Y�/�.L"���پԄ��g��>Vv�?̦=i@�:\��X��������¾��<�|��P �>Q>>I�������u��{\�"���f{�z�ƽ\٧>᩾>�.?$�?k�w?<?cu%?�M'��?�$k=¤$?�5"?�'�>�?���>;��>�P�>;�f>D�h>�%ٽ�kn��4Y=��=j-;>�M�=g>�=�+x>N�ٽm۠�s�޽P0ƽ�eU�y��<���=�d�=�W>zC>��?.�<?3�c�(K~��ha�a��UȽK��$>� �=K��4�0>���>��?�Z?x�>��мQ��T��'�ﾭ����1$?*�a?94E?�}�<˫.>�L2�0�����>%�>�>;_��1�����9�==�t�>�^�>�>Ė>�y?O�b?W�"?Mɹ�i*i�jc����@�L>�}J>ZAy>jj�>Y�>���Z����@���KX��DϾֹ��=(�>�&�=Wc�>F�g>���=(:�>��N�}��	���I�¯�=؎}>#�?t��>�%�~�~�
v��I?�롾v����qmо����)>�=>����?�����}���7>=����>�|�?��?5!d?�\C�"��Ew\>��V>K�>�-<�>�'��vl���2>���=	/y�8
����;��\>v�x>��ɽ/�ʾď侃J�����2Z���"�?g�������b¾��xW�����O缁Ѿ�݂���6� #$�v���it������Z��5G���F�?X�?T#)>�s���,�{)�QU��h��=پ�����l���[�c�b�0!Ͼs־�X	�71���6����k*�>�V����H}��H)�W���Mm<>��.?d,ƾ�o��R��H�`=�n%>�w�<Yﾓ�������(��)V?,v9?A��Q��Q޽P>Np?���>_�#>�f��E��A��>s�4?��-?>�μ�����狿M���A>�?&��?��??��I���@�������?u	?���>B ��E1˾�꽪�?��:?㕽>+��V���0J�"f�>3�Z?|�M��_>��>�P�>D�ٽݒ��<�������c����;>�����V�e��U<�A��=唢>�w>��^�59���8�>�;��N�ʳG�J0������<*4?��.>�nj>�\>��(��������,��
]L?���?�oS?�h8?#6��B�좩�QH�=S��>��>��=�k���>���>�����q�����?۩�?��?��Y?l�m��ؿ�ʚ��mӾ-����=���=��$>�E��h=�=
�=f<
	�= ��>��=Q�>��>�5>R�>>V̆��d$��S������F�խ�~�	�i������
ݐ��#�>�������|;��0��G�r���@Z���C���ܾ�UI=��>�l�>G��>*��=Y�W>*�����-���R4�����^�����(���F�����V(��c�
Z�� ��#?%��<���;��>�ޏ���=C�>��}>d)�=�>΀>2T=z�>�Ã>/Ǜ>��>��u>l��>X.�>C���.��r�k�CU�֕�f�S?�[��I��m��O�c�����S>S��>pBK�pnN��X��OӒ��*�>T�*=kؾd�oD�=�$~>�)?�P����>&��ٟ�<]/�;O�5>,�+?��>�η>�#
��/�=�r��?���[�G>_�?�H%?�c_?w�W?���>ͩ�>����>��=���=2>~I.?��7?�{^?��=?*T�=:껽��=�+K=��[��c���_=Fa�<\�ػ�=5�ҽh`�(ms��6��>-�=�8����p=���<��>�@?��?wo�>��g��C���D��0��-��=�L!�d�>��?�qB?͍�>7�>�{���I�<$9��\
���>ܲ2>bs��t���;ff�>K]�>�>?=�"?�A�ɮ�oY>}&�=�H�>��>��?=�>
�s>}E�=-s
���ҿh-�����d��t���4c=7�i�}'ۼ���=i;+�0@!�ܣ ��>�#�>J:�>n�>�J1>��>L��>0��=
�>zx�=?4�c�E=yyͽm�c=�
���S�=/}Ž݅�=!�<�҆�R���B����<¡P��=x�G�?R?��'��b��f�;����������>��>CY�>ճ�>,�=�%��hU��vA�wG��E�>
qh?,��>l�8�_��=8�0��PT:�γ>4��>��>�`�2���U���>�<9��>͔?�O�>��V:[��to�c�
��/�>��\�v�is�?�K?c��DQ�nO�/~8�k�K��i�<���	`,�aۆ���c�@�`��N��O����YK=��>�<�?	�G��җ�dؾ�����=����j�	%,=p�>$NE>Yv%=�����Y�� RB��|>�Ք��$��K_�<=!�=��> r?�?��_?Z8?Mk
?7y�����>�p�>�L%?2!	?��>�?��>'"�>�.�>� �=(�=��!�hƮ���;2��=�x= ��<5��=}f=K��=�{=�>�v�|��}\=>=��"=m��= e=�L>�@�>��K?KB��H���^��0rT�wx����-�]�>��=q�׽��=���>��6?�O5?���>�<��ھ�c����ә����??�gY?��#?_�v� ���<���׾]`�<�>$�K>>c������ح��,��>�5�>�[�>OU@>��{?R�_?V�?n��gP� <���l/�*�m�c##<�GX>�T�>x�>��־P�;�.����p�3<���5�*�Ր�<O�K>��="��=.X(>��>�G>�˽�u�$�������>�֠>�/�>�Z�<P}c>��������I?���y�2A����о���x>R�>>>��J?2��O�}� ��+&=�3��>5b�?D��?�Kd?a�B�%���]>6�V>�>R�/<�'>�������� 3>���=��y�����6��;��\>��x>��ǽ�ʾ�PE�2���O�Z�w<�Ͼh��=�¾�&���")�{ɕ�2K�x�ƾ��%��p��#n��(]M���\�q������TB�3	�?pf�?.�>:���������n%>p���z���۟������q��\��3����H���E1�x-F� ����>�yY�AA��(�|���(�L����{?>�3/?�[ƾ�̴�"����g=j%>� �<�6�B���[�����\W?x�9?	O쾆*������>�?{w�>.�%>[$���'��+�>�94?��-?��뼰���6��&����l�?V��?{;?T�*�=h=�K����ֽ"f	?!
?a�>�5���eپUԣ�R�?B�<?��>GX�f��%�����>XS?7�G�3XD>3�>j�>����·O�󝈼����uM(���s> b�<y�����>�>��Ź=[��>�S>�MN��?��b��>�?�_�N���H����d���v�<�?>��1>�i>B>`�(�Y���ω��'�_�L?	��?��S?tk8?^�����ͬ�����=��>"Ӭ>���=\����>���>�h��xr�'�ܘ?�I�?V��?�[Z?��m��dο�	���q��оp�*>_y�=��>z
$>��Ka��P���N���=K�>E<�>�q�>��>
�>�Gv>e����#�qƪ�yь�=�O���n�
no�Q<*��x��5����D���*+�=��=���� �5�"�=���z��=���>('�>MͰ>�i4>��?>�qt��d���|�H���=��:+��e���C�]����l?K�?z��qs��^����>�'X<�:�=��>�m��g,>�˓>Ń�=��>` >��3>X�>��*>V8>��->��+>]�	>:i�>��>��I��(��v�q��^ ��6�yKz? �ǾQ��ӏ��@2��?D�SR3�Ec�=6ɗ�s:v��@���8��F�>,��S��n:�����S�>�B ?���ND->Ru������wf���Z>o�,?3�>�,>��9Nս��ֽR��>y{��A�<X�>�O?-=5?�	L?�(>��"?P��=�l�>z>�V�<��>���>��?�??U?��?F�+>��p����%_�;��]�u�����=��=��S���=*w��҅=�l>G=�Q�=�+���*�۽Q7�;>V?^zB?�?E��>�ܱ��y%��,��?�<>��<�2?V�>�:�>��?�S�>�5�=L����򳾹@����>�>r>J���b��~���h�>_�>�h?��?y����Yݼ��<AZ�=F�i>(q�>�=?E�?3��>N+�>8a뿃����~k�L��x��=g�O��=��I��t�7���2��x��������>���>2�>�ג>W�?��>��>L�>�J�=��!>�4ֽ����i�@�7����=[x�=�=�=潦|���p�c�ӽ�{���%
�,���|?�? G#�����nf�L���$�����>���>���>/��>B��=^Q��;R���>��=B����>&g?���>��6�9��=�D�8qѻ>i�>�V>�q�
M"�?���%��<=��><,?�5�>�a�c�X���n��H��>�U�=q1����?ѿZ?������7��F���T��-�=ھ��k�¾2漨KT�̫m�Y�/�.L"���پԄ��g��>Vv�?̦=i@�:\��X��������¾��<�|��P �>Q>>I�������u��{\�"���f{�z�ƽ\٧>᩾>�.?$�?k�w?<?cu%?�M'��?�$k=¤$?�5"?�'�>�?���>;��>�P�>;�f>D�h>�%ٽ�kn��4Y=��=j-;>�M�=g>�=�+x>N�ٽm۠�s�޽P0ƽ�eU�y��<���=�d�=�W>zC>��?.�<?3�c�(K~��ha�a��UȽK��$>� �=K��4�0>���>��?�Z?x�>��мQ��T��'�ﾭ����1$?*�a?94E?�}�<˫.>�L2�0�����>%�>�>;_��1�����9�==�t�>�^�>�>Ė>�y?O�b?W�"?Mɹ�i*i�jc����@�L>�}J>ZAy>jj�>Y�>���Z����@���KX��DϾֹ��=(�>�&�=Wc�>F�g>���=(:�>��N�}��	���I�¯�=؎}>#�?t��>�%�~�~�
v��I?�롾v����qmо����)>�=>����?�����}���7>=����>�|�?��?5!d?�\C�"��Ew\>��V>K�>�-<�>�'��vl���2>���=	/y�8
����;��\>v�x>��ɽ/�ʾď侃J�����2Z���"�?g�������b¾��xW�����O缁Ѿ�݂���6� #$�v���it������Z��5G���F�?X�?T#)>�s���,�{)�QU��h��=پ�����l���[�c�b�0!Ͼs־�X	�71���6����k*�>�V����H}��H)�W���Mm<>��.?d,ƾ�o��R��H�`=�n%>�w�<Yﾓ�������(��)V?,v9?A��Q��Q޽P>Np?���>_�#>�f��E��A��>s�4?��-?>�μ�����狿M���A>�?&��?��??��I���@�������?u	?���>B ��E1˾�꽪�?��:?㕽>+��V���0J�"f�>3�Z?|�M��_>��>�P�>D�ٽݒ��<�������c����;>�����V�e��U<�A��=唢>�w>��^�59���8�>�;��N�ʳG�J0������<*4?��.>�nj>�\>��(��������,��
]L?���?�oS?�h8?#6��B�좩�QH�=S��>��>��=�k���>���>�����q�����?۩�?��?��Y?l�m��ؿ�ʚ��mӾ-����=���=��$>�E��h=�=
�=f<
	�= ��>��=Q�>��>�5>R�>>V̆��d$��S������F�խ�~�	�i������
ݐ��#�>�������|;��0��G�r���@Z���C���ܾ�UI=��>�l�>G��>*��=Y�W>*�����-���R4�����^�����(���F�����V(��c�
Z�� ��#?%��<���;��>�ޏ���=C�>��}>d)�=�>΀>2T=z�>�Ã>/Ǜ>��>��u>l��>X.�>C���.��r�k�CU�֕�f�S?�[��I��m��O�c�����S>S��>pBK�pnN��X��OӒ��*�>T�*=kؾd�oD�=�$~>�)?�P����>&��ٟ�<]/�;O�5>,�+?��>�η>�#
��/�=�r��?���[�G>_�?�H%?�c_?w�W?���>ͩ�>����>��=���=2>~I.?��7?�{^?��=?*T�=:껽��=�+K=��[��c���_=Fa�<\�ػ�=5�ҽh`�(ms��6��>-�=�8����p=���<��>�@?��?wo�>��g��C���D��0��-��=�L!�d�>��?�qB?͍�>7�>�{���I�<$9��\
���>ܲ2>bs��t���;ff�>K]�>�>?=�"?�A�ɮ�oY>}&�=�H�>��>��?=�>
�s>}E�=-s
���ҿh-�����d��t���4c=7�i�}'ۼ���=i;+�0@!�ܣ ��>�#�>J:�>n�>�J1>��>L��>0��=
�>zx�=?4�c�E=yyͽm�c=�
���S�=/}Ž݅�=!�<�҆�R���B����<¡P��=x�G�?R?��'��b��f�;����������>��>CY�>ճ�>,�=�%��hU��vA�wG��E�>
qh?,��>l�8�_��=8�0��PT:�γ>4��>��>�`�2���U���>�<9��>͔?�O�>��V:[��to�c�
��/�>��\�v�is�?�K?c��DQ�nO�/~8�k�K��i�<���	`,�aۆ���c�@�`��N��O����YK=��>�<�?	�G��җ�dؾ�����=����j�	%,=p�>$NE>Yv%=�����Y�� RB��|>�Ք��$��K_�<=!�=��> r?�?��_?Z8?Mk
?7y�����>�p�>�L%?2!	?��>�?��>'"�>�.�>� �=(�=��!�hƮ���;2��=�x= ��<5��=}f=K��=�{=�>�v�|��}\=>=��"=m��= e=�L>�@�>��K?KB��H���^��0rT�wx����-�]�>��=q�׽��=���>��6?�O5?���>�<��ھ�c����ә����??�gY?��#?_�v� ���<���׾]`�<�>$�K>>c������ح��,��>�5�>�[�>OU@>��{?R�_?V�?n��gP� <���l/�*�m�c##<�GX>�T�>x�>��־P�;�.����p�3<���5�*�Ր�<O�K>��="��=.X(>��>�G>�˽�u�$�������>�֠>�/�>�Z�<P}c>��������I?���y�2A����о���x>R�>>>��J?2��O�}� ��+&=�3��>5b�?D��?�Kd?a�B�%���]>6�V>�>R�/<�'>�������� 3>���=��y�����6��;��\>��x>��ǽ�ʾ�PE�2���O�Z�w<�Ͼh��=�¾�&���")�{ɕ�2K�x�ƾ��%��p��#n��(]M���\�q������TB�3	�?pf�?.�>:���������n%>p���z���۟������q��\��3����H���E1�x-F� ����>�yY�AA��(�|���(�L����{?>�3/?�[ƾ�̴�"����g=j%>� �<�6�B���[�����\W?x�9?	O쾆*������>�?{w�>.�%>[$���'��+�>�94?��-?��뼰���6��&����l�?V��?{;?T�*�=h=�K����ֽ"f	?!
?a�>�5���eپUԣ�R�?B�<?��>GX�f��%�����>XS?7�G�3XD>3�>j�>����·O�󝈼����uM(���s> b�<y�����>�>��Ź=[��>�S>�MN��?��"��>OA�{�N��H����[��CQ�<�?h���5>�i>�A>(�(�����ω�p*���L?욱?E�S?l8?^�����ᱧ�͘�=��> Ӭ>D��=�����>���>�f�]xr�
�Z�?�J�?���?\Z?��m� 0ʿ*ϓ�6޸�ͶϾ�K�=���={V;>M\���>A�X=Z�Q���c�T��=_�~>��G>���>._U>�6>��/>�߉���%��w���q����J��������U<����M��&�Q�ݾ�d;��꽳E���?���-�ߪ ��w.�Mؠ��6>]^*?�$�>{c<>���=�t3><����̾oLS�����X���b���C��]yS�����W�������녽�-�+}�>W>j>f*�>VW;
�>���>p�:>g�J>/ý>�yT>!i>���>�4�>Φe>X�>�,�=��{>�F�=&��w���v:���Q��;!�C?dr]��]����3�'f߾)����>��?��S>*�'�鸔�C�x���>��F��b�F�˽$ �[�>���>��=��ǻO�n�w��Z�;�=8��>�>b�l�`񏾿'�C٘=,�(?L���k��ȇ>D�;?5pq?��4?���>�X�=nm��B�>�p1<@��>�?��>�m?��G?$�&?�?ַ#=����ݸ�0=;�ս̼�}���7���2����y���<��=II=�=��=oȉ��<�o.=�^�>�&?���>w�>���8UR�ld��T��f�v>c�:>f�a>U�??Ȼ>�[�>_�?�ٹ>��:�����{���3�>�l�>��R�����ݖν�6�=��c>Ͷ]?��0?�i��c�[�S|������>��>C�>[�?b�?�VA>�;��Կo�*��%�hq.�%�J����<2oA�gu��N��+�a���r�<�vl>̵{>��>39G>C�!>�E>.��>�o7>�N,=��=�l�z�u�y2\�5tT;Z�<�
����0��=�2�4��s&����lm�������	?�F+?�Vƽ2iþ��K�ZB��eቾ��>a�%?�3?Οc>N���+���O$�&*���Q��\?�Y{?�q	?�B�ҡ߻�b�j>�r?K�?»�=��*f$�Vb��c��=�y�>0�"?V��>D��#>��	;�����>:�G��;���?�:c?ܾ���-k\�Q�k���)�("f<ae��|$<�h��qA%��DW���"��&,�XD��\�v\�>�,�?u<�<6���k�)���;ߜ�[Q��P��N(t=P?�Ō<�h�� 띾8�Q��_:��Qg����A-�=��a>�A>	Ӳ>$�?��o?Q�?O?:`�=���>�:=)�?��>e�?yI?���>c:u>p�>�	)>�4>4���B��D�Ž�O:�ʩ=	pa>��>�/����Q��)�� >9D�2X�L>߼�/[=��(>ոI>{�>�?N�!?\
�3��Z=�iӽ2"��ԉ$>tT�>�f3>�ؒ�m+���>x��>��?�+�>K� >�匾3_���뾆<o�W�?n�??ޥ?�Ԓ<�W8=�ž˝�g`a=zC�>CA =� |��A�l(��n8��jL>j�>�:�=W�̽瓏?l��?�)~>�s�|�M�gZ������ �Ծ`#�ʘ�>�w�
%�@�i�Bw���}���ķ��K3��	#����B�̷�=�N�=����P�>W��>�&>�l�=]�ؽ�Ͻ �2�W��>|��>�!?f��>]�7=_{u��Ѿ��I?�2��q]�脡���о5i �l�>nj=>/�s�?oD���}������'=��}�>�l�?3��?zZd?��C���Y�\>��U>H�>Y:<aa=�i���ڄ�y4>���=��y��P���;z>]>xx>�Cʽ=wʾ���J D���п�����������Ju����I�z�?��4�^�l��V+��W=��c�u�H�P{�ju=KЋ��� ,����?w�?�|�>My>��6��~P�p�����L�;���k��=m'6�QK��������&3l��f��;;��ٛ>6�V������}�R )������?>�b/?��ľ=Y������
e=%e$>ϙ�<;�v��(:��q
��V?��9?br뾥p��}E�t>؉?�\�>��'>-�V�\�>�O3?��-?t�N)��x-���Ry��z�?�$�?�|>?r�=��T@���
�����?=�?}��>;�m��9����
�1�?�;?*m�>{��%�����<�>&�\?/�M���N>���>���>�:ɽjޒ� �c��G����B�M�;>��»�v
�ٌ_���B�'+�=���>�Gi>��l�gŤ�"��>OA�{�N��H����[��CQ�<�?h���5>�i>�A>(�(�����ω�p*���L?욱?E�S?l8?^�����ᱧ�͘�=��> Ӭ>D��=�����>���>�f�]xr�
�Z�?�J�?���?\Z?��m� 0ʿ*ϓ�6޸�ͶϾ�K�=���={V;>M\���>A�X=Z�Q���c�T��=_�~>��G>���>._U>�6>��/>�߉���%��w���q����J��������U<����M��&�Q�ݾ�d;��꽳E���?���-�ߪ ��w.�Mؠ��6>]^*?�$�>{c<>���=�t3><����̾oLS�����X���b���C��]yS�����W�������녽�-�+}�>W>j>f*�>VW;
�>���>p�:>g�J>/ý>�yT>!i>���>�4�>Φe>X�>�,�=��{>�F�=&��w���v:���Q��;!�C?dr]��]����3�'f߾)����>��?��S>*�'�鸔�C�x���>��F��b�F�˽$ �[�>���>��=��ǻO�n�w��Z�;�=8��>�>b�l�`񏾿'�C٘=,�(?L���k��ȇ>D�;?5pq?��4?���>�X�=nm��B�>�p1<@��>�?��>�m?��G?$�&?�?ַ#=����ݸ�0=;�ս̼�}���7���2����y���<��=II=�=��=oȉ��<�o.=�^�>�&?���>w�>���8UR�ld��T��f�v>c�:>f�a>U�??Ȼ>�[�>_�?�ٹ>��:�����{���3�>�l�>��R�����ݖν�6�=��c>Ͷ]?��0?�i��c�[�S|������>��>C�>[�?b�?�VA>�;��Կo�*��%�hq.�%�J����<2oA�gu��N��+�a���r�<�vl>̵{>��>39G>C�!>�E>.��>�o7>�N,=��=�l�z�u�y2\�5tT;Z�<�
����0��=�2�4��s&����lm�������	?�F+?�Vƽ2iþ��K�ZB��eቾ��>a�%?�3?Οc>N���+���O$�&*���Q��\?�Y{?�q	?�B�ҡ߻�b�j>�r?K�?»�=��*f$�Vb��c��=�y�>0�"?V��>D��#>��	;�����>:�G��;���?�:c?ܾ���-k\�Q�k���)�("f<ae��|$<�h��qA%��DW���"��&,�XD��\�v\�>�,�?u<�<6���k�)���;ߜ�[Q��P��N(t=P?�Ō<�h�� 띾8�Q��_:��Qg����A-�=��a>�A>	Ӳ>$�?��o?Q�?O?:`�=���>�:=)�?��>e�?yI?���>c:u>p�>�	)>�4>4���B��D�Ž�O:�ʩ=	pa>��>�/����Q��)�� >9D�2X�L>߼�/[=��(>ոI>{�>�?N�!?\
�3��Z=�iӽ2"��ԉ$>tT�>�f3>�ؒ�m+���>x��>��?�+�>K� >�匾3_���뾆<o�W�?n�??ޥ?�Ԓ<�W8=�ž˝�g`a=zC�>CA =� |��A�l(��n8��jL>j�>�:�=W�̽瓏?l��?�)~>�s�|�M�gZ������ �Ծ`#�ʘ�>�w�
%�@�i�Bw���}���ķ��K3��	#����B�̷�=�N�=����P�>W��>�&>�l�=]�ؽ�Ͻ �2�W��>|��>�!?f��>]�7=_{u��Ѿ��I?�2��q]�脡���о5i �l�>nj=>/�s�?oD���}������'=��}�>�l�?3��?zZd?��C���Y�\>��U>H�>Y:<aa=�i���ڄ�y4>���=��y��P���;z>]>xx>�Cʽ=wʾ���J D���п�����������Ju����I�z�?��4�^�l��V+��W=��c�u�H�P{�ju=KЋ��� ,����?w�?�|�>My>��6��~P�p�����L�;���k��=m'6�QK��������&3l��f��;;��ٛ>6�V������}�R )������?>�b/?��ľ=Y������
e=%e$>ϙ�<;�v��(:��q
��V?��9?br뾥p��}E�t>؉?�\�>��'>-�V�\�>�O3?��-?t�N)��x-���Ry��z�?�$�?�|>?r�=��T@���
�����?=�?}��>;�m��9����
�1�?�;?*m�>{��%�����<�>&�\?/�M���N>���>���>�:ɽjޒ� �c��G����B�M�;>��»�v
�ٌ_���B�'+�=���>�Gi>��l�gŤ�"��>OA�{�N��H����[��CQ�<�?h���5>�i>�A>(�(�����ω�p*���L?욱?E�S?l8?^�����ᱧ�͘�=��> Ӭ>D��=�����>���>�f�]xr�
�Z�?�J�?���?\Z?��m� 0ʿ*ϓ�6޸�ͶϾ�K�=���={V;>M\���>A�X=Z�Q���c�T��=_�~>��G>���>._U>�6>��/>�߉���%��w���q����J��������U<����M��&�Q�ݾ�d;��꽳E���?���-�ߪ ��w.�Mؠ��6>]^*?�$�>{c<>���=�t3><����̾oLS�����X���b���C��]yS�����W�������녽�-�+}�>W>j>f*�>VW;
�>���>p�:>g�J>/ý>�yT>!i>���>�4�>Φe>X�>�,�=��{>�F�=&��w���v:���Q��;!�C?dr]��]����3�'f߾)����>��?��S>*�'�鸔�C�x���>��F��b�F�˽$ �[�>���>��=��ǻO�n�w��Z�;�=8��>�>b�l�`񏾿'�C٘=,�(?L���k��ȇ>D�;?5pq?��4?���>�X�=nm��B�>�p1<@��>�?��>�m?��G?$�&?�?ַ#=����ݸ�0=;�ս̼�}���7���2����y���<��=II=�=��=oȉ��<�o.=�^�>�&?���>w�>���8UR�ld��T��f�v>c�:>f�a>U�??Ȼ>�[�>_�?�ٹ>��:�����{���3�>�l�>��R�����ݖν�6�=��c>Ͷ]?��0?�i��c�[�S|������>��>C�>[�?b�?�VA>�;��Կo�*��%�hq.�%�J����<2oA�gu��N��+�a���r�<�vl>̵{>��>39G>C�!>�E>.��>�o7>�N,=��=�l�z�u�y2\�5tT;Z�<�
����0��=�2�4��s&����lm�������	?�F+?�Vƽ2iþ��K�ZB��eቾ��>a�%?�3?Οc>N���+���O$�&*���Q��\?�Y{?�q	?�B�ҡ߻�b�j>�r?K�?»�=��*f$�Vb��c��=�y�>0�"?V��>D��#>��	;�����>:�G��;���?�:c?ܾ���-k\�Q�k���)�("f<ae��|$<�h��qA%��DW���"��&,�XD��\�v\�>�,�?u<�<6���k�)���;ߜ�[Q��P��N(t=P?�Ō<�h�� 띾8�Q��_:��Qg����A-�=��a>�A>	Ӳ>$�?��o?Q�?O?:`�=���>�:=)�?��>e�?yI?���>c:u>p�>�	)>�4>4���B��D�Ž�O:�ʩ=	pa>��>�/����Q��)�� >9D�2X�L>߼�/[=��(>ոI>{�>�?N�!?\
�3��Z=�iӽ2"��ԉ$>tT�>�f3>�ؒ�m+���>x��>��?�+�>K� >�匾3_���뾆<o�W�?n�??ޥ?�Ԓ<�W8=�ž˝�g`a=zC�>CA =� |��A�l(��n8��jL>j�>�:�=W�̽瓏?l��?�)~>�s�|�M�gZ������ �Ծ`#�ʘ�>�w�
%�@�i�Bw���}���ķ��K3��	#����B�̷�=�N�=����P�>W��>�&>�l�=]�ؽ�Ͻ �2�W��>|��>�!?f��>]�7=_{u��Ѿ��I?�2��q]�脡���о5i �l�>nj=>/�s�?oD���}������'=��}�>�l�?3��?zZd?��C���Y�\>��U>H�>Y:<aa=�i���ڄ�y4>���=��y��P���;z>]>xx>�Cʽ=wʾ���J D���п�����������Ju����I�z�?��4�^�l��V+��W=��c�u�H�P{�ju=KЋ��� ,����?w�?�|�>My>��6��~P�p�����L�;���k��=m'6�QK��������&3l��f��;;��ٛ>6�V������}�R )������?>�b/?��ľ=Y������
e=%e$>ϙ�<;�v��(:��q
��V?��9?br뾥p��}E�t>؉?�\�>��'>-�V�\�>�O3?��-?t�N)��x-���Ry��z�?�$�?�|>?r�=��T@���
�����?=�?}��>;�m��9����
�1�?�;?*m�>{��%�����<�>&�\?/�M���N>���>���>�:ɽjޒ� �c��G����B�M�;>��»�v
�ٌ_���B�'+�=���>�Gi>��l�gŤ�S��>�쾃(H�#G�����42�8��;���>���6>T>,�>d-�����/ϊ�5��SLE?n�?�V?�>7?1��q��B���M=>j�>"��>Lv�=<H�
��>b�>�.���r��w���?l��?Eu�?HU?V{e�����Ϸy�l�L��(T�C�~>H�=�9F>����Y�=ēl;��<�n�<��=���>�8e>��w>��N>�-<>�>�7���������ѫ����@�{J���6����yd;gK���:�@��럾��9��2���s�C����W��9�"� �� ����>��>g���1��o#��۾��h�Y���}ԾI�־]\%��� � ������Vľf�E�m<
�^�!=F�����>�ۏ���=Me�>�$�<����u��=lv�>!��>��i�=�9>Gƣ>���>�T>�kQ=_,��ۂ>�H>s�� ̊��T=�X|�l�\;�8*?G5��>�J�%A<��i�M�}�g	�>�e?h<{>� !�Z.��R���O��>=TU=Ԑ�(��
���О>�E?^;J>Z�=���P=�4��Ay�@9=��S>�13>ZՔ=�]>� 7o�O�w=V�?����>g��>Ú-?�o?�P?wx�>C�X��-�3??'�>�d�>��>of�>��)?��]?$"L?�}>�>����",>`�D>I����H�M���E=v����xӽ:�<Ⱥ�=rG�4�ɺv���D������>�=n�=?e�>��"?V��>��>u9���)�CiX�?����`c>�)�<_��>I&>H�?��?��>�5>��c����kn���>��>�E��	x���"�"��>%��>�c?�X?��*w����Ľ?�<>�?��-?�<Q?iR�>�G:<h �-��Vjӿ�$���!�)��A���@�;L�<���M����8��-�w������<	t\>>�>�up>��D>�>R3>�R�>�OG>�̈́=k�=]9�;�e;`�E��M=9�DG<��P��l���AƼ��������l�I���>��M�bټ�	?�?l���Ye��`t��3���	����}�>�7�>@�>p��>�-�=�|���W��nC���W����>	�a?�?�B/��-�=GR��2<��>Ѡ�>!�>RfC�݉�٥��z<��>x�?�Ş>�7���Z�?�l��t	��>é9<[`�p:�?�c[?����.���b�}fC��!�Q*�<>,����Z��������):/��4���� �$h�dެ=1l�>��?|\���w<Тþ$����w�Ft�C=��=0��>z�>�3��v�6
��Ƹ��qL��b��z>C�>�Ƚ>� ?�k?� `?��?%�?��ܽ���>h�F=o��>���>m?��	?.��>�|>AL�>�]�=F��)��'�}����<�W���t�=s�>x�>������=���<`M=�f� �T�짨�Q��;(��<��="W=#��=��
?�@G?.=о�W����h=��g=��`>s�B>MY�>��P>@V�yJ.�I�\>��>/];?,�?RJ�>�ž+��ܴ����:��� ?G95?5	?,��=N8>����J�˾8ѐ<B�>��M>�%<��.�됾�#�r���>#��>Ma_>v)=%aT?�n(?n��>J����'���i����=əͽ�'C>�,�>�=콶�`&N��:��d�c���'�/�Z>TA��?
�;����>�ɩ>Q��=�o���"t��{<�Ⱦ�K߽eV
��C?C{�>��>���=��<+����g�R�I?h���8=�Oˠ�uо�����>#k=>8���h?Ud
���}�[ڥ���<����>�q�?���?3
d?b D�EY��]>�MV>��>.3)<�W?��������I�3>z��=�x�����Y�;�}\>kx>߷ʽ.�ʾ����jF�:���G@��=�G���>{��w�� ���P��X��L<���s�ʽ9���*Rf��8�������1Ͼ�����O�i8?��0?�h�=�2���O���(� e�ж�@�e����<ҕƾ������оAO �o���y/�9L�����?�>��]��ˏ�'ez��.*����U3>a
,?����̱��&�fr�=pa>�`<<|������Wi����
��IX?�{8?+��y��.�齳�>w�?iT�>�&>�'����뽨��>��2?�1*?+��������׊�J���7X�?_'�?R�??�M��T@��	����J? 
?��>Kj���ѾL��N�?w�9?���>�����������>��Z?�|K�r`>���>I�>ğ佫a��Q�0��Õ���X�K�5>5�Ļi��9�h�q@���=Q�>O�v>�^_����k�>����N�TtH�9��̱�9��<�? ��><�h>�>/�(�aŌ�����b&��tL?/O�?��R?�;8?�U��y;�.;�����=���>m�>�G�=��
�/P�>�?�>���x�q�ϑ�Fi?e�?a�?�Z?��l�bVȿʌ�䔏��j����<O�=��9>�I��<,�=�>�<��
����<��=p��>I�\>;LS>h�>�\�=�M>�܆�G:"�H���	����^�\4>����(R����$�n��	��[���~��������,/]����`���ܽ���z�����>��@>ɼ4>�ǫ>��,>ϝؽ��>�]wԽ0��:}����$��}���:�Y%n�>����%B��(���=�.׾��>���ǉ�����>��=04=P�T>j�#�A>�&��h�<0�	>��=Z#>$�
>m׆>��=(���\l>�Η��藿���8�¾��T�z+=?{N>�w��}�6�_$��a>=j3�>�g^=	������rM�A�Ӊ�>�$�bt�	��<��z> 6�>�L>�i>��;�fr=_R��]�<�D<>��2=�`�>��<����@Y��ࡎ>�H�>n�*�T.�>\+�>�5?��U?�[?����>�>+�Q>I(�>/7���Q��s�><?��?xI\?m)?��=ygT<��u<�-�=���X	��iW��<�<g�[���5=	J>-U;X��=o������E(�<��l<X'+=��=K�>�#?%x�>��>/����^���e�vO��JF>ꋽ�O�>2�>�?�V?s�L>z�=��s�����_6�bN�>�]�>7-z�K۔���=�I�>�~�>u�X?�<0?�l۽C�g���<;��L���>]��>�2?p��>iէ>,6������̿-�!�:�,����8��<�_Խ��\�5E*=N�*���O�֖�<�YZ>]|h>�Ov><�b>�f>	A>BZ�>]�_>��=�=���;ڃ¼s�ý���<�����<{Y.�19=�4�: 1��j��^<*�u~�<�༟z�Ѯ?�?���D�b��yY����Z���ٿ>G��>�>�:�>�Զ=����CR���8�
�+��=�>��a?H�?��3
>
4��2<��>�-�>_' >��$�`�/�?���6�<��>|�?��>��:��\�q�n�~�X&�>":���w��bȅ?eic?�H�.c�5�wYS�NFԾmy�=�
�q�u*8�E���A�K�&�j~��滾���?�;�?
����_��K�A�Qɏ�LB���'������Wm�/7?s�>�*�=a��=��y���-�������B�����;>C��>�j+?C�!?X�U?�)?p�?e���U��>ⵟ=9b�>EP�>%�?e�"?�?>�M>ip!>]�����=�������8w�=�(:K�=��=#{Y>�����=�#>�|e�[a�<]ZI�RɎ;$��="�B=��4=��=+`>I8?:�C?�2ؽ��>8�F>;2</ݼ��Q>z+n=� ;� ���!<��>��-?�
�>[]�>3�V>��ɾ`����˾�=�_@?TH%?u��>��X�w*o><����EL�
Xb>4Z������̾ۗھ����g(�\�Z>ћ�>&�¼d>��|?T7C??� ?����v+��"v���*��t�w6��u�>��>���=�ھ��3���n�CO_�@�2��W���A����<���=H�>�o3>�=�>B�<!��@�ƽ��<� ��T(�>���>k.	?�'Q>J�`=d>���"���:?�͝�2�
����A�޾B=z� (�=�>>�Fӽ�P?��M�b�����,�K��>��?���?�a?Y�4���/�>7J�>m7>>`�=�b��3��<
�e>�J�=d}[�<b����0R>o�>�Jg���Ǿ��a�p��ح���+�^6��AM����
��J��s�����5�?»��۾�ڟ������ ��-%�{2���̾����a��H�"?A�>?���=�h��~D��}A�-3� p��Js��#��O���^��I!C�����۩�� �?�2����X�$>C�8��p���Z�������HG=�.?�y����o���!��==x*5>6F�����`H���닿�4��<?2_%?kZ�}\�_��� >�D&?Mn
?5w>ط��������>�A%?�Z�>����^7���5����Ͻڂ�?�վ?��Q?��R��S[���쾣�� ?|`�>J��>a���*������<��
?��;?�Ѿ>A��?sl�9���K�>� I?iQc��	'>��>l�>8ȶ��yX�Dt����*m5=f�>Tz�����͘����L�>�2�>�=�>*�!�독�:Y�>`��%O���H�)��������<�8?���>�i>�>��(������Ή�r�2�L?[}�?S?�\8?�������E���dא=��>�ʬ>:�=~�ͱ�>���>��n5r��D��@?�)�?R��?�%Z?�um�H��d���eo)���&�V�K>	�>Y#D>�-�����=��μ�e>�;��=R+�>��k>F�>�>X\o>uag>�����#�x����2��,�:�l���66�!u������d��̶�
������ۦ�tW�����1���R���S۽2����_>a�>I�>/� >TqE=h�M=s�;�X�HWy�š޾ʸ�>%��!�|�ԾI������kƵ�q���p�����?E	{>@PZ>&��>T�<��>��f>�0��yQ>ϜX>��=K�?>�(�>u�>��0>��>�u=���=�-_>狁�(3��G�J��U���J����>�ޕ����O�"����ڗ̾5=>
�>-�;'0�Si����x����>S���B�������~�Y��>"]�>�џ=����+��t�/��ؼ�=j+:>od>��)�P�{����DD�=I1?�ȹ���g=U�>>4?�?�cU?���>��?m$�7��>)P�>p>�>���>{�>J�1?��U?�D?�0?�t>�H�3�ڽ���=�ԣ=�W�� ��`���(T�������`=��EF<ݺ&=l��<)=*�ڼ�h�=�ns=��>�t"?�>��>�F���;��X��@��v��Ɖ���� ?��>��3?�v?&?nx=o�(���O���!�>�=�6�	��e�����?�9�>x1~?�tR?0�ѽ_����c>��$>I��>���>��d?�U?��>fy�>#��mӿ�$�D�!���P�݈;v�<���M��U�7!�-�V���ș�<#�\>B�>��p>�E>��>�<3>�R�>�HG>�ф=)�=E;�;ގ;'�E�"�M=�
�-DG<d�P�.����$Ƽ
�������I���>�[:�}8ټ��?�k?��)�H2����f�!���X�� ��>�K�>lZ�>H��>���=}e�e�U�q�A���G�[Y�>�dh?-@�>n�8�2�=�,���:��>`�>�8>g�a����Ϙ�^��<f��>0�?��>u���;[��fo���
�T�>�V(= 	�R�?�`?���)��� �nNH�a����="�꽔^[��i��=�"��7�]������[v��=��>߼�?y1u�#��=p>�������D��Y�����R=aCw=g��>�F>��1�|���X��3Ҿl1J�T��<�Y�>-�=���>��?W�?��T?��$?�&?=##=|U&?1v�=T7�>WA�>��?ω?�?�X�>��>�M>Y�#=��˽Rt���'��8=��>sX->0�5>���<N(�=@Ⱦ=J[=D*&����|G/���W��G<༮=�>Y[�=߯?�Q"?-`ӽ�/C���"�.3���<>�NP>$���p�k�uW�;�J]>��>��.?��>�Dw=-�پl��~��^��=��?��3?�A�>��T;�:�=���F����O�=��P> �m�鉾���5��&\ ��w�>�Ӑ>��=���=��?�?8��>�|��C:�˲l�:�23���<�S�>�>l�@�u���|A�O�w��c�KJG���R�z�ͽ�=xG>_3>���=��>9�y>�i�=ߐʼS��.{r�`iѼ��>zH�>��!?��?>�.������u����I?ߜ���i�L�jrоEO���>�<>8�v�?N����}�����G=�Ë�>5��?��?�>d?��C�P/���\>�KV>��>�/<��>�
 �5���n�3>��=]y�����;G]>�Ey>��ɽ��ʾ�4���H�Zĵ�gN���?�\����=��c��_���(����x�x�=� ۾ʬ�r%���ǽ�Zþ��u�پ��B�,$�7?l��?�������4��?�"t
�Q�yp��@=�=qS¾|�罜�E��ݾ�ﾆR'��������4��(�>)3H�'N���$��"*���=��v>@ #?�N¾@���1 ��=S	>���<NZ�ǌ�p~���F�.{F?��8?o�Ӿ���������=4�?'E�>��>ZЧ������L�>�V;?�y.?��i�ύ�v��B�<}�?��?1�??f�O���A�
�����0?��?d��>����s�̾�h�L?@�9?P��>P��b���3�� �>+�[?�=N��Qb>���>�N�>I�ｦ�����%�)��뙅�w�9>#H	���EYh��>���=�	�>��x>��\�������>˾�U��T�C�	�q<��Y@�����>}@;�*>/�p>��=����艿�k���e8��]>?�
�?�$Y?��4?�
�3cپ؃��d�= 2�>P��>-4�=%���W�>U�>�3뾧�j�S
�98?BN�?�8�?��]?��m�A�oS��%���C�Ⱦ�2->��h=�h>�o��@�'��2�=����p@>"e�>�>�9�>�Rk>��V>>�:>�ނ�/������ul��NZ9������4���ҡ��s\�*�2в��펾�!q�q/��S�"��i��E4��=N�����=1w
?&�>�Xn>;=I>�D>+������H��������-�@$�����ž��=�2C����]����P�;�!�#�?e�=�S�<F8�>�����=��>�'�=�v�=��\>��=H��=pd�=㧉>|�=ah>��=��{>7�=�g��Wn��8�:�d�S��M;�A? �e�����4U1�=4ݾ�3���G�>:?��N>��%��󔿡iy�ٳ�>�6[�~0_�	���h9T��O�>���> P�={ᆼ�e%��t�ҩ��=�~�>
>����!��������=�>{{��,>��>�T?U�U?T�E?¡�>y�>�M�<S�>eQ�=��A>�m�>��>��#?Mw[?��;?qi�>�w>z�0�h��<���=�B:�`�`�Kޛ�_#>+��	��<!����TF<�w=����'h=��o=��==��M���K�>q�>?�T�>+�>U�<�qDH���J�h�P�ʚ=W�%�н>���>�Q�>F�>��>�k�=������_�#l�>��+>C:��p�J��"�>C�A>}P`?��?�T�y	/�w&M<P��=f*	?}�)?��+?���>�U=4]�Ȝ��Dڿ)<�&>+�fi<խ<�!N�<�sP�����%�\��J#�[j�={�>�+�>t`�>Ն >P[>��L>y^�>�_>:>+q�=�B|=�g=�ꋽ�*��V|<4�=Q�X�1�b=Eǯ�tֽ׬��2^��殮�76��q3���??X�)?���E�,�ɽ��l�ɾ��辝�>ʲ�>��8?�m>�4��	��It���D�2����j�>��w?9~?��[��ؼp�:=��>�)�>���xa�>�������BᇾS����%?��>^\�>�����'�qw���?���>��:�1��,��?AT?>S���þ�R�H	ƾ�jѾ2���h�,6Ľ#i�2:!��4R�0e����5�@r�(��=��?���?��ؾ�ｌ���u������.�����&=�y�=��>�5�>�Η=�_�=\�U<��U`��QB���>~S+>9k5=Ƚ?$3?X�x?T)�>k\7?�`>_�>�-���!?\��>8��>�/:?i�(?D��>�?i�f>�P���z46���6���:Ύ�=M�=`�5>"��>�zB>������۵�X�S �=N�X�I=K
p<�%>ur>�� ?tc?�="w{=0�2��S��g
Z>���T>��)�����<k��>n�>���>�5?�0�>�o>�����OL��sؾF�X=�?G$?I�?��
=_�W>X��������=|g�>?:�<�^�����R��W�=�dn>�|�> �>~�>¾j?���>U?�+6���A�+�8��a��ֽ�>۰򽂐�>�u�=���$3��a�He9���2�eՇ���Ho�=�HX> �<�1>�w=qM�=�(�=,t��zs�S£>��=r\	>�|�>!�%?C�=>'��>i��tT��I?����Nj�d�sо�M���>��<>����?z��$�}�|��YH=�͋�>Έ�?���?
?d?�C�f(���\>:OV>��>m
/<��>�!�����g�3>_�=~y�����,�;o]>�Ey>��ɽO�ʾ�3��H�H8����D�F���ѵ�N�����<�e�M��=/���J�(7ྻˎ�ȷ�9y ��庽�彽����d��������?�C?��v>�+=��P�/{�����
>z�c��Wz�|_�����y��{������p��ӂ3���-�)���2�>���<X���7��ʆA�\�=�(����>=lh���K$,���=#�=��e��A����ᝠ�y􋾄�v?R�?}�_��3@������@+�i�r?G9�>E���ӗ�� z�O��>2��=D#:?o9>?dB�x���)�a�?i�? �6? J�=�wl�[�V�<����;V?�� >�X>�Nw=\d�#�F��'���H?�>�������`�-���:?�?�Nǽz�u>���>kq>{�<I^��,���n}_���>ؒ�>o�;)�����)�Ow��g�>`�>���>y��=�gо:Y�>`��%O���H�)��������<�8?���>�i>�>��(������Ή�r�2�L?[}�?S?�\8?�������E���dא=��>�ʬ>:�=~�ͱ�>���>��n5r��D��@?�)�?R��?�%Z?�um�H��d���eo)���&�V�K>	�>Y#D>�-�����=��μ�e>�;��=R+�>��k>F�>�>X\o>uag>�����#�x����2��,�:�l���66�!u������d��̶�
������ۦ�tW�����1���R���S۽2����_>a�>I�>/� >TqE=h�M=s�;�X�HWy�š޾ʸ�>%��!�|�ԾI������kƵ�q���p�����?E	{>@PZ>&��>T�<��>��f>�0��yQ>ϜX>��=K�?>�(�>u�>��0>��>�u=���=�-_>狁�(3��G�J��U���J����>�ޕ����O�"����ڗ̾5=>
�>-�;'0�Si����x����>S���B�������~�Y��>"]�>�џ=����+��t�/��ؼ�=j+:>od>��)�P�{����DD�=I1?�ȹ���g=U�>>4?�?�cU?���>��?m$�7��>)P�>p>�>���>{�>J�1?��U?�D?�0?�t>�H�3�ڽ���=�ԣ=�W�� ��`���(T�������`=��EF<ݺ&=l��<)=*�ڼ�h�=�ns=��>�t"?�>��>�F���;��X��@��v��Ɖ���� ?��>��3?�v?&?nx=o�(���O���!�>�=�6�	��e�����?�9�>x1~?�tR?0�ѽ_����c>��$>I��>���>��d?�U?��>fy�>#��mӿ�$�D�!���P�݈;v�<���M��U�7!�-�V���ș�<#�\>B�>��p>�E>��>�<3>�R�>�HG>�ф=)�=E;�;ގ;'�E�"�M=�
�-DG<d�P�.����$Ƽ
�������I���>�[:�}8ټ��?�k?��)�H2����f�!���X�� ��>�K�>lZ�>H��>���=}e�e�U�q�A���G�[Y�>�dh?-@�>n�8�2�=�,���:��>`�>�8>g�a����Ϙ�^��<f��>0�?��>u���;[��fo���
�T�>�V(= 	�R�?�`?���)��� �nNH�a����="�꽔^[��i��=�"��7�]������[v��=��>߼�?y1u�#��=p>�������D��Y�����R=aCw=g��>�F>��1�|���X��3Ҿl1J�T��<�Y�>-�=���>��?W�?��T?��$?�&?=##=|U&?1v�=T7�>WA�>��?ω?�?�X�>��>�M>Y�#=��˽Rt���'��8=��>sX->0�5>���<N(�=@Ⱦ=J[=D*&����|G/���W��G<༮=�>Y[�=߯?�Q"?-`ӽ�/C���"�.3���<>�NP>$���p�k�uW�;�J]>��>��.?��>�Dw=-�پl��~��^��=��?��3?�A�>��T;�:�=���F����O�=��P> �m�鉾���5��&\ ��w�>�Ӑ>��=���=��?�?8��>�|��C:�˲l�:�23���<�S�>�>l�@�u���|A�O�w��c�KJG���R�z�ͽ�=xG>_3>���=��>9�y>�i�=ߐʼS��.{r�`iѼ��>zH�>��!?��?>�.������u����I?ߜ���i�L�jrоEO���>�<>8�v�?N����}�����G=�Ë�>5��?��?�>d?��C�P/���\>�KV>��>�/<��>�
 �5���n�3>��=]y�����;G]>�Ey>��ɽ��ʾ�4���H�Zĵ�gN���?�\����=��c��_���(����x�x�=� ۾ʬ�r%���ǽ�Zþ��u�پ��B�,$�7?l��?�������4��?�"t
�Q�yp��@=�=qS¾|�罜�E��ݾ�ﾆR'��������4��(�>)3H�'N���$��"*���=��v>@ #?�N¾@���1 ��=S	>���<NZ�ǌ�p~���F�.{F?��8?o�Ӿ���������=4�?'E�>��>ZЧ������L�>�V;?�y.?��i�ύ�v��B�<}�?��?1�??f�O���A�
�����0?��?d��>����s�̾�h�L?@�9?P��>P��b���3�� �>+�[?�=N��Qb>���>�N�>I�ｦ�����%�)��뙅�w�9>#H	���EYh��>���=�	�>��x>��\�������>˾�U��T�C�	�q<��Y@�����>}@;�*>/�p>��=����艿�k���e8��]>?�
�?�$Y?��4?�
�3cپ؃��d�= 2�>P��>-4�=%���W�>U�>�3뾧�j�S
�98?BN�?�8�?��]?��m�A�oS��%���C�Ⱦ�2->��h=�h>�o��@�'��2�=����p@>"e�>�>�9�>�Rk>��V>>�:>�ނ�/������ul��NZ9������4���ҡ��s\�*�2в��펾�!q�q/��S�"��i��E4��=N�����=1w
?&�>�Xn>;=I>�D>+������H��������-�@$�����ž��=�2C����]����P�;�!�#�?e�=�S�<F8�>�����=��>�'�=�v�=��\>��=H��=pd�=㧉>|�=ah>��=��{>7�=�g��Wn��8�:�d�S��M;�A? �e�����4U1�=4ݾ�3���G�>:?��N>��%��󔿡iy�ٳ�>�6[�~0_�	���h9T��O�>���> P�={ᆼ�e%��t�ҩ��=�~�>
>����!��������=�>{{��,>��>�T?U�U?T�E?¡�>y�>�M�<S�>eQ�=��A>�m�>��>��#?Mw[?��;?qi�>�w>z�0�h��<���=�B:�`�`�Kޛ�_#>+��	��<!����TF<�w=����'h=��o=��==��M���K�>q�>?�T�>+�>U�<�qDH���J�h�P�ʚ=W�%�н>���>�Q�>F�>��>�k�=������_�#l�>��+>C:��p�J��"�>C�A>}P`?��?�T�y	/�w&M<P��=f*	?}�)?��+?���>�U=4]�Ȝ��Dڿ)<�&>+�fi<խ<�!N�<�sP�����%�\��J#�[j�={�>�+�>t`�>Ն >P[>��L>y^�>�_>:>+q�=�B|=�g=�ꋽ�*��V|<4�=Q�X�1�b=Eǯ�tֽ׬��2^��殮�76��q3���??X�)?���E�,�ɽ��l�ɾ��辝�>ʲ�>��8?�m>�4��	��It���D�2����j�>��w?9~?��[��ؼp�:=��>�)�>���xa�>�������BᇾS����%?��>^\�>�����'�qw���?���>��:�1��,��?AT?>S���þ�R�H	ƾ�jѾ2���h�,6Ľ#i�2:!��4R�0e����5�@r�(��=��?���?��ؾ�ｌ���u������.�����&=�y�=��>�5�>�Η=�_�=\�U<��U`��QB���>~S+>9k5=Ƚ?$3?X�x?T)�>k\7?�`>_�>�-���!?\��>8��>�/:?i�(?D��>�?i�f>�P���z46���6���:Ύ�=M�=`�5>"��>�zB>������۵�X�S �=N�X�I=K
p<�%>ur>�� ?tc?�="w{=0�2��S��g
Z>���T>��)�����<k��>n�>���>�5?�0�>�o>�����OL��sؾF�X=�?G$?I�?��
=_�W>X��������=|g�>?:�<�^�����R��W�=�dn>�|�> �>~�>¾j?���>U?�+6���A�+�8��a��ֽ�>۰򽂐�>�u�=���$3��a�He9���2�eՇ���Ho�=�HX> �<�1>�w=qM�=�(�=,t��zs�S£>��=r\	>�|�>!�%?C�=>'��>i��tT��I?����Nj�d�sо�M���>��<>����?z��$�}�|��YH=�͋�>Έ�?���?
?d?�C�f(���\>:OV>��>m
/<��>�!�����g�3>_�=~y�����,�;o]>�Ey>��ɽO�ʾ�3��H�H8����D�F���ѵ�N�����<�e�M��=/���J�(7ྻˎ�ȷ�9y ��庽�彽����d��������?�C?��v>�+=��P�/{�����
>z�c��Wz�|_�����y��{������p��ӂ3���-�)���2�>���<X���7��ʆA�\�=�(����>=lh���K$,���=#�=��e��A����ᝠ�y􋾄�v?R�?}�_��3@������@+�i�r?G9�>E���ӗ�� z�O��>2��=D#:?o9>?dB�x���)�a�?i�? �6? J�=�wl�[�V�<����;V?�� >�X>�Nw=\d�#�F��'���H?�>�������`�-���:?�?�Nǽz�u>���>kq>{�<I^��,���n}_���>ؒ�>o�;)�����)�Ow��g�>`�>���>y��=�gо]��>A�l�N�ͪH����3���L�<��?)���5>�i>A>�(�����ω��+�.�L?���?g�S?�k8?�]�����9���㙐={��>�Ҭ>�=���*�>���>�f辒xr��ę?�J�?n��?�[Z?5�m����K���6ZվJ���f>ō>�c>XK*=_�����dF1>�}>S�>4�?�¡>�Ŭ>mv�>|��>�S�=�%~��"�F��,����:�M���7�!c�"*%�(�e��۾����$ʥ�-����ҽ� �=);��-ɼvA�;'�ɾ�+g=�?���>t+?�/�>Nw>��B��j�Y�3�j���X�!��	�&�Ҿ����i�G��}��C��������=!�꾟�'?�f�;�*�=��>�&轱�>f_�>�l�=?�=���=� >�7>���<���>�G�=�)>k0�=�|>A�=�ل�JI����:�1�P���;��B?�Z�[k����2�O�� `���ӄ>e�?��Q>�0'�̈́���Ax�8��>dA��/c�[�Ͻ%�(�/n�>�W�>�J�=��g����Y@u����� �=��>�>��g��M���*�N	�=T�>H����-�=�m>"�!?X�h?�^;?0�=��>��@>�Y�>4>ɉ_>�j]>�>E�?s�??:�6?YP�>ګ�=x��~��<=E>���]�f�䭖���Ƽ~:���<��N�U.�=�r�=��3�6Y0=�	�=	�5����<HV�=�
?��H?\�>U>�=����
�A.$��8¾�XM<��D;x�0>�{�>`�>-�>(�>�[>��1<�����#���>�IT>�W�Ӄ����S��b�>x�>ps�?Gi?��@?�t(Žy��=�>?�#7?� H?�?��>h=½E������N�eɾ�cK�t��>�"�>l�=�_���1��h>�5��/��>&��>���>S�>HR�>'&>��>��>$��=��������9����;*��<4஼7���������B��f�;�B����<ϴC���7�Z�	�t!=G?x ?$j���-�>/վ�*���3��h�>�[�>џ?��"?𙷽�z,��G\��e��D����>�7+?a�?s�� >��5xܽ�9V>�?:b>����S��z��$N�	W=>2?q0�>B�ݽ?2X�FB`�&����>9>f�	�-t�?��K?�:�r����g�["�"���̑.�@�=�9Ƚ��þd�
�V�R��Ǿ./%��K�V��=%z?���?������E��k�sA����ß���5W>S�B>��?�"=>�۰����Ѷm�{�<�64˾�Gýq��>�<�>���>�J?I!s?�'s?�T�>�nG?^�=�h#?YGd� �>�?��'?��?�c?oV�>���>�e�>p`�8y�w�����=�OJ>���>Ġi>���=���=�ݥ=���=�"1=����L ��O�=��	��~�s�����;�4>�?�\8?�&���Ŏ��_�����P>К>d�>mټ�/�������=�t?9@?j7?���>ܓB�I�#��LȾN-����>�5b?B�>Ś��RC>�����4h���o���>7�H>ݸ��]�e�����\�I��>Q4�>�4q> ,�>[�|?��&?��?��=Q��8)e���|��O��9��>~y>�;=q�K�1�n!�AHx�h�Z���X�\���/6&���=y�>o:U<�H>q� =��>��7��g�x)μ��>>�p���">ş�>;��>@[�>��>�׾�)�N�I?Vt���c����Nkо�.���>��<>|��!�?4���}�����1=���>%��?���?:d?�'D�_�L�\>RHV>[>`.<P�>�\X�A��/�3>b��=�?y����C`�;]�\>�\y>�Vɽz�ʾ�侞"H��(���L��cx����N�O�@ĕ�Ce��7���6�R�������K�ē'��*��1@��g���������;��Gʐ?!}^?5ܧ>����SD#�lGѾ���L߁�:]��N���9ɇ�W/r�#z��Q�ʾ�ݾ���O�2�"�O� ��V��>�\<�Y��Á���a��%>␽r<�>����
�#¿�I.�����=:�=�I�7�~���t̡�ǫ�((�?*o%?P伾Q���+��n{>*�?�?2��>�:��[�|�|��R0%? d?���$qH��W��wCr����?�"�?3�J?�k�<��*�C^�0�q�؛)?y�>+��>l+��V�����Z�>�k?�#��4#�?n����L���>���?�@��7>OB�>*�>h`>�\���+$=�[ؾ�5���9�<a�ν��D=:���1r��H�>7��>�h?>��������>����D�9��j�)�!��>��,����0�>�Ψ�~�)>���>x<V�@�+��ʡ���y�=�	?�?��s?uo)?z$ �����k?�E8>���>��>��>>��t=e�>�.?xr���U������3?�E�?TH�?��R?f">�s^ѿ�������Ҿa�>j��=�~>���u�Q>�>lƽE���Gl�=8G�>�ay>�w�>��>PR�>_�=�܆�S�%�i@������.k��� �A���wh���[n潼s�L��n3���v�=J6�<�{ �@@ͼ�H���E/�����Z),>�x?�U�>*/�>
ug>0>>�֝����&܍�:��o�	���9�޾��ľ|�d��G
��,���t��}"��i[�u��>���<��A>P��>�
$<��&>Oz�>��"=�آ=��
>���=ĸ:>�Y.>v�]>��>�?+><>έy>��=�_�����9�bKO�,,�;��C?g�_��)��¼3���߾LO��T{�>r?�T>�-'��S��k�x�(��>,F��!`�+�ʽ���Nl�>ix�>-6�=��ʻ����z�7O�1g�=�>Z�>j����6�����T��=��?4����{P�>ΙH?#�v?bv?�g�>�'?e�����=* ��D,��݈=���>�OU?E�Q?W"3?�		?C=�=�n��a<RD!;��6���w����N"�=���>�>��'=���?j��sĻ'�u=�==�`�>�,>�� ?��;?I��>�X�>@[�Tc5���3��)����q=#н��>���>l�?��>o��>g�>�j��������&*�>��>�T���d�8��� �d>ԏ >�6?O�%?�oU��p.��>tn>�q�>�?�t	?���>��k>ߨ��iO��{ҿ��v�x�V�
��=�ަ>e4H��U�>����Y
?����Nx���p�X>hO?{�$>��>�N�>ȝS��?�>��c=��>��=���<<�>��5��hT>�<��r�>=�<H =AV�<�^#��s�8,�=8Z,�������� ?h�?#�
�����>q
�ͅ4���� ?��*?�|?��S? r> f&�� c��zT�=ֻ��=�H?4~_?������Y=v�<9R�>�`c>,V>���=�~̽8��־�	ļI�>�2�>�/\>q�q��[2���B��J��8�=E�<��E �>Ġ?�}.?X7��!��rG��t���:�pj>K��/��>
��ذQ�p�c�v�Q���1�#i�=�kN>��?��?��t�S���ｿ�{�������>)W��ŏ�>=q�>1)��J����t���I�W- �H���� ?t��>|[�>ƍ?�1?9�3?F��>W�!?��۾Q�(>�U�=�?>��I?�Q?�/_?J��>��>36>�g�̠ؾ�~��Z��j�d�𯚽��<�V�=��j>)�]>�v>�=e�d<G�vA�>�= g>Η�=��<���=��=e�?c�?��'<b;�=���=]U��~�O>�Y�;2>��a�J�G��=D��>a?(4$?:�>��=X���<����پ����q�>�!?�| ? #3>I6�>������}��]��9g��J6���Ծ���H����w�k��>�p�>I�,>��>b��?u6?��>wn����p� 	y�:�P���:�9��<���>� �=@<�=��w�W���m���e�"��~��=[�̽z:�=���<m!��u��>ũ>8�>D�s��h2�c���]�>�=M9�>�?���>諵>o[�>2v��6��rkI?ʬ��\E�nW����˾"��.�>WfD>��q�?�(	��}�b�����;�`��>.��?
�?�d?
r=����w�\>�Z>u%>l�<�/?���1�f��XV2>ø�=��u�J�#:$HX>�v>��Ͻ�u̾y���G��	��{`�sp�C�׾��f�G���o���Z
�z���X��_���&���z�O�����o��S���*b�L4f�����K�?[׀?�[E>��+�Ya1�����ᾝY]<2����=����݀��Q���2���Uj#��3����/ξ�o�>K�=�˾��X뀿�?-��N���>�S+?���i⮾"��P�=��>/���s�\Ì�^N�����g[?�|6?Mt�e��)��Q>�-
?�{�>��+>�y���C߽�ޟ>��*?ԕ%? ����������1�qH�?�?B�??�JN�"fA�<[�M��ԅ?^?���>(��c}̾l���
?�D9?h��>Յ�1l��2�����>��[?��M�S�a>T\�>�]�>�0�Sk��5O$��蒾eK��Bq9>��߻�J���h��<�Z�=��>�x>R\�����,��>!�����H��f�@h	�\Ds�[�� >"?ࡾ[�>mG�>�M.>;�'7��[���/����/&?Rg�?�Zs?+�)?8�f���f�Ž��=�4`>LR�>V'>��ӽ���>Sl?�淾�o�� Ǿ#�+?�]�?!J�?�6O?�Yj�+@ӿ�Y�����(�ɾb�>�7�==lI>���Ӂ>��=U��iT���+>�[�>��>f	�>my�>�p�>&�>6��h�%������ы�-�B��>�q ������̽��Y��`�)h�?�N�� 0��qԽ���/�=���X�,�dq��0��9P?(��>
>>�ƛ>G�8>B���xS���I?��XT�@վ6_�������[���V����оV����-���>��-�u�3>�z�>B�C���=�1>e.�=�j,>�ʍ>;��>ۋb>�܉>+�W>���<��?>D蓻�w>�#w=����fG�y�6�x6F���<��C?��Y��뛾E�2���9)���'�>��	?�X>F�%��K��6�v�H��>ݐ^���i�:�Խ�%���>���>��=�R���?���hv��S��9�=OT�>�z	>��8�I=�����l4�=5~�>	�ľ���b{�=dfY?:7c?=�|?��>Z��>ė>��>�B���ل�=��>Cu%?�?�r?��+?,��>1]�=����*�߽Z���s���Yf	�mߖ��ks=�/�=Y�t=2/v�-B�=67�=��=f�Ǻ��z=E��;,A�>0�>6?��d?æ�>ї=x2-��h��'z�Ԥ����=��>�N	?�>^z-?W��>��>�ML<�Ħ�7�Ӿ���ԗ>��`>t�$�r�X��<�<�Ű>���>�X?א?L	�������>�!�=�(?x??��3?�X?9	�=�j��O	�=�˿+zn�v�>�zC,�=������>�~$�> �=��{}�=��>��>Ӊ>P�>�N�>a5K>8i�$>�>���=��>2=*>Nh���>�}��n,K=��Y�vX�M�=�A���=��ؼ�.+�=�r��җ��4��A�$?��2?Zp�+ݾ"լ��@�&=�2�+?�3?<]J?|�?W�= �;�E�|���q�M0� ����%�?(\a?i�����=N���>>? �>�>[���5˾�ѾP���&=��>�02>�Y�N��ǖ�v��N�>'�������?�+\?a�X��
j������8�sA��I�<��8<�¾�`�� ���G������<N�@�۾����H?[q�?���EWԽ%@��� ���b��m�>��>_޴=?�^>������$�G�C�QD�຾���>��?_�y>#Ʃ>�?��0?�%w?IL?5�1?=�d������Pʾ�*��;%�>o��>Z�?���>煙>1d�>5=������rg��>�q>�W����=q��<��>�m>�����0�=|ŗ=�����9ɽ�}�x��=`��=�轼��=A��=�?-�3?:��S=��D�!(�<���=oß������+�rH��7�>T�=9?�y?��>�0�>��߀!��4Ⱦ�N��v�>��P?*�>G�>�ϳ>�9پkM�։q�D���I�=L���߹����پ�T�2�>� >�0�=`�>��?�u?l�?;�
��d��t���%�
<~�%�N=��5>��=m��;D9�0��(��:;i�����"�=N�����=6]>���%NC�6=|��p=н��:{�<+�G>�x�=MP?#�>��A?���>��>bU����B�qOI?=ѡ�K����N˾�����>2jC>�����?�����~�C(��m<����>h�?Z�?7Uc?!A���HY>X�N>��>�<w=����r�y��-:>��=ˤs�X��:�0<_|^>��y>ľ���žɅ��9��!�����M�<�̽t���=3���g��Jϼ�����{�bӾ�����N<,[^�k�p>8��B򻾅�B�sE�?$/a?��?)">o p������.��� �� _Ҿp���W�����ھ1
Ͼ�*¾��c�d�L�2�5��� �>ޔ����t��x�%�?�u��������:(?O����%��yL�=Q�=�l(=�4���Z3�Q��|{��)��=�q?4^4?J����?!��2���.f>p�?h(�>P\�>���������>� 3?I� ?	UY;�d������t=R��?D�?��??n�>��A�e�w���� ?Zm?�K�>r�����žq�����	?'�3?{�>7q�������K��>�]?UHM�Dz]>IU�>��>H�ٽz����e)�����	���8>Y����6c���9���=��>"kv>�d�@ா�C�>M-m�Z�Q�ɇ��� ����Y��)?߁��z��>z��>ټU>{�b��9������w��i��>D��?@zy?3�"?J�վT�{s�7ʖ>f�=f��>��=��%=z�?9�$?�/\��U@��0�R?N?�Y�?Iv�?�3<?�m�׿���������о�nE>��=�� >�?+�xK>?�=?�>�v޻V��=慍>?ň>t,�>N�T>�E�>�k^>ކ��S&��ج�Hn����)�e������N��Hξk#��⮾����E���p����,m��]��J���Ԅ�?޽G�Ҿ�|V���1?���>�ǅ=!�>ߕy=e�վ�����kľ����'�=�����|ھ���=�#��|�ľ�h��9�;��K�>Sm��K�>~�?�#C>C�r>�3�>�>V��N�=��>
�j>��>0%�>i�=�j>��I=�Dy>��=~r�������9���S��=��sA?7�[�ZY����2��t۾"���"��>��	?�rU>��&�a�����x����>T�O���]�#�ӽ5����>Gn�>�w�=G'������y�����Ч=5�>֠>�r�׵��y���=H��>)ү�ί��Z>0?�!j?��s?���>��>b!�<��=�1-��������>h��>�k�>g�H?��F?KQ�>�c:=oI�l� ;������v�w�ý�P��'w>$�6>��#=����e���<�%�g�=5@=xM�=�����k�=F��={�?�G?0�>]�> r���c�h�_��=���>���uн>A�?F?�%�>9M?��=��o�+�徱k��5�>dc4>`v6��l�/�=CDp>��
>��P?E�	?�j>'�V�Э���l>;?o"%?��?��>7��=(~8����ҿ�lU�<�T�� ���>j<^��3.8>��=;L>��h�1���8>6��>�b�>@܇>���=$g">(u�>͡=>j�z>��8>��h��>�d�]��<55�Oٿ��V;��]r�d�p=䅎��yT��\
����<xe.�"�_= Q#?&8<?����g>	�,A̾�G�+���?�<?fX?�P1?�>�>Ba4���v�^�V����1�5= ��?--*?<��H>/	��!��>���>�A>� �=������¾������{G�>� ?�TJ>��$�i���&��D+�y��=���ͶZ�*��?��??��G��ǂ��0�g�-��_-��?s>�׾42���:���W��@�j�3I�����_e2>}�? ��?Ђ���:����[(���И���̾?40�y�>K�>���>Y������^q0�d]��oԾ�ݨ=��>�c]>g�>��?wxH?o�T?3`�>xo/?��:�!ۻ�� S����>Ǘ�>��#?�_�>�ͱ>_��>{���9ؾ�M���h�E��dpĽ��&=��>��2>�>1>$�+=5Z�=��	>��5�����_4�ʖ�;aN�=w�>�3M>��`>Ƶ?ouB?�,���g�F�b>8�,�)�/��͊�U�O�������<��y=���>A0?u�P?T4	>�\�>��>�D�ʾ�	��;�>�!)?�[?��>�o
?>s�:֯�=鴽v�5>_��!���:��f/쾨�8<�>���>p">£>��?���>y��>�(�ڪ^������66�
����(8��׼>�;#?�]o<�!��s��=t�EM���-�M���x�B���;")(>�!>�S=��=V�b=�:ڽ�Oּ�Z�ND��� �=�� ?]�?v.5?��>�o�=��辪FB�w�I?�����m��⠾�Hо9��$>D?=>��"�?[����}����c6=���>�|�?���?Ed?C�����\>�DV>E�>�-<\�>�7�������3>�:�=��y�B���ݛ;�]>�3y>t>ʽ��ʾ�/�DH�5V����p��f�Ѹ}��&��o��̾<�</���E/�� �'��{���u������R<��n��k��\c��Y�?��?h��>�/.>��>�נ�9���������v�� ���������1��Y������9�U�#F�(J�p�>v�q���p�^w���M�	<ݽ�t�3?�<���
O��*��z�=dC����u��n9�`������Ř<m�o?$�/?�	��~g� �ܾ�.>.? ��>�>�N���L���>s�?&o�>$�>����+�}��Ȍ��O�?�0�?��>?q�G��
A���*�� ?a�?���>�K����ɾ����+?:/6??x�>�����-m�*��>��Y?��M��aZ>��>,ǖ>?R��뚕�C�+�����K���66>;�����r�`�+0�[h�=E��>�Rp>��`��w�����>����N���J�f-�ŋ"�R�r<|3?�)��
>�p>kL>�)��:��H����Z�>J?ֱ?�\T?]�7?����~�쾯7����=��>�3�>���=��6��>���>����qp���?tv�?j2�?�X?	�l�-iӿ�����&������4Q>��>�'�>;����Q�=� +=�k�=��=���=�6�>9�>��>��s>��>=�->���;:$��B��x���ݱ����������ù�
ڋ�9���L��j8`�l����򽄅�m!R�wԩ�`����k?��>KY>�y�>�!>	�����ܾ\�Ѿ������h��A肾�^���Q5��u�Z����ξ�P <֮����>�j��զO�y��>��ʭf>l�>�pX=s� ��M>w�>�.�>]HC=:�>�y>��>���=s.9>�����Ou��uj���A����D�u�E?
w��B�����=���9�Z�Q�>^��>���>/�����8m�P��>{b��3b�Ff	��7��H�}>��>��>��m<2�\��"��2���0>���>��=CF�=�2���*��:>f��>���ʛ�=A"�>u?2��?T�G?r�h>R��>�ho=��	>���=�>Y�>5\&>�r3?UO?�g	?r��>�	>�q3>��==㜾Ģ��$�=���=�%����=nd����=���=s�z���=u$�>G�̽�$���/ >=�?�Z??�jE>1�>�U�a5X���g�9$��"'�>�z�<X>�C�>:4�>��>�N?Od=�����Ѿ���>�|\>~�8�3�X�<)8>�k>��=F(?�?��>��(�K��DX>� ?@?DN�>f��>e_>����	�e:ο2�!���=/}�=e�=D�=��}>c�-��(��aFc���g>�-�>�l>pi�>wo�>�be>�>?�>��[>��<�o5>]\+��t��f�Y=�^">:���M�(��0"���\�����B�P��h=������!?��D?�Yh��0��`վ��4�)��?��>
?S�4?Ҩ>��-���w���h���4�@���َ?a�Y?P�����=hݞ��ח<?��>ם>ԙR>��<i�Խ>���\ǅ>�>�%�>�
�>�h]>��4۾a�ƾ��&>�1X=�$n����?g`T?D5�����+����*�8��>z����Ӿ��<�Y(�m�T�VKD�(3��;��e4>��?��?�r��{��)�w��7��ʽ����l��>z�>��>3��4uA�F�P�M3.�
��g�t>FK
?0Y>�w�>I�	?��0?_'�?�O)?xM?&�3���=g���/p>��5>���>X2�>��?��>L_�>���I-����ɽ3����n=ʐ��$}�=�c>�k>7�2>H��=��Q=/����޽a��|+=�)t<�j�<`[�<#�l>��3>�?p5?����������v>9�4���<����b��ʟ�%�X:fZE�3/��Y�+?��Y?)�F>��=�����7��L��{':����>�?^�
?j��>X��>J.��:ξ�iսW�t>&q�����ʍ����Ծ�
=�n�>溥>�w(��l�>"s?iq�>q?�����H�˽e���2�폼�U���>�?�������'S�h�R���3�Mh�<P�:�Z����*�<�vE>�`I=�w�=@��=���
��?I���x��o�����>sY�>ykL?R��>$�R��V��U,�M�I?���#k�w堾�^оs����>��<>���?�����}�h	���A=���>���?���?N>d?�C��(�^�\>�IV>��>IZ/<ݒ>�����k����3>k�=�y����#I�;��\>�9y>uɽs�ʾ�.侤_H�H̼���c�����Cj&������X������Z\=�Vݻ0�p�g�i���S�sA����(��7��ҽ��ľ/Ej����?!�e?���>���=�lb�
Ѿ;�ᾃ'����N{�ځ�?<�Q;����䜾Ď꾸'_���6�x4
��7�>h�������s{��|0�%dԽ!��=�$?�q��9`W�p�/��#>^Q�=\��W��w{��"���PO_���h?��4?�>�����#��*S>	?h�>���>f����V���>6?*�?�N=<�����?K�<�0�?���?�;A??փ��9�.)�1J��v�>m��>�?y�MO����=b�?}�? �l>��~���k��?��m?�lH��><>�9�>�[�>���9����<8�>��N����8�=%�⼬���	J>�����>�>�,�><��I쪾��>��޾��H�6BL�cD
��"+��:Z�?�o�=�>��U>�I>(����1�������E?2J�?Q�S?4@7?���b>���i˽.��=x�>�ݨ>���=����h�>�:�>��޾��q�4�����?�6�?��?z�[?�m��̷ֿ��;���Uھ̆S>}�=h�c>�1�����=��=N<>��>�U(�;���>��>e]�>��D>⹘>ڧ�>+P���&�)p���1���2�f��������_������D���ݮ����Y�V��L��*�~�:�ľ�/]����=����h#����><|�>(x�>��i>��>�!���4�BD��[�=�L$��{ؾ�U�� Ӿ�?5���c�Ⴞ?��G��<�-�����>T7;0;�n*?Ѥ�<�~�>��>���=�zֽ[>}֧>u�>�>៳>�Y�=!v�>��>Ԁw>��=.��������:��T��׉98zC?5�Y�sЗ�7G1�E�۾�������>�?�OT>��'�(���Vw���>hN�<kZ�_1ǽ�G��a�>yd�> n�=����̼[~��|�}g�=n�>Y
>c[���������ҍ=�s�>��˾=����a�>��F?��?�u?}�>��$?-�k��f��l��w ^;=�>M��=�H!?��?M�?���=��=dL��>0�~CZ��J��������;�=�>K��=J�6o�O=�>�3=>#l�=�m��bs�=�M�<�5?Q�D?�%�>�̘>�Y�mHR��[p�
{��>�����>'|�>��?p��>�[?��O=���������B�>ׯ�>�%�Зs���!>U��>��0<�F?l[,?	d�>&��i�D�{>�)?AU?�h�>�y�>�Z>�c������οV�/�ES�yQ�׃><���+>��.��p��=�z>��G��T����>޶>�΄>���=�9E>��>���>Df�=T]<>��=$c����O<e�����=�_�=F>�D�<�R,>� \=�=�� �r�c]	�y� =k���y�^*?^?���=��A������K�5��'�?���>NK7?�YV>`+?��0�&l��ˈ�xE��ڼG�?�/?����q�#>�'5��V#�/_�>D}>���="������㷾qB>�}�>�9�>�A�>�&�=�������Q����@>��<π��h�?x�>?�_�0⥾\<!����?8���>�;���.��BH>��^�x)5���X�8��$��N�>�U?�b�?2~�T�3�YU��?3��Ziv�:�w�nKܽ�J���=�Ce>ɚ�w����{A��2M��Q��q*�=&��>֤*>��L>{�?T�P?.�j?�H?�o+?'~�4�>�.i�%>.�>� �>d9 ?��>ec�>��>�o��(���Ž��B��!�=cm�<��E�mO=2�> �|>)���_� X���h��/�ϼ@��W6���/�<ec�=�>�cE>$�?b�7?9�(=�T�xf>g��<�Ѽ�1�ȣ=�j<�(+,��n�YI�>a/?>P?げ>4;>�	��)W�<���Ĵн!�>�??�?Y&�>K'(?愭�:���(����>�B]>����%�ק��=�?a�>�j=�ٱ>ۅ}?��?׺>������a��4{�~.���Ҽ�����9>o��>d��<�#�����U�=#Z��OC�1�<�nR�����R:G�H��>�T�>Ʉ!<�Y�>��)=NSt�g��=G��\ʱ>���>5>0?'��>B�	>���,�:�vI?����X��W��*`;Z��l>�&B>.T���?Q�e�}�����Q�<�fe�>/X�?��?��c?T�C����,rY>6�M>�|>� <):����2����6>���=|(y�N��ʐ�;�Q]>��x>��Ľ��ǾT�⾟�>��ſ�n�v�C�oĞ�7�;���cﺾ|,˽>ړ�&�^=�.�;k������ˌ����8�Խ&l���;Ⱦ"E�;L��?]{n?��?���=}M;�H���%[սIL��586=N��O���������ھ ����˾�q^�G�-��־ɕ�>σI�����[~�S�,������b.>�.?�SǾjӨ�ex�-Չ=��>��=�����f��Κ������(Y?�#9?�8ᾍp��2�
�J�!>�U	?��>�p+>���љ�͑>V5?�)?{<ϼ�L��oΊ��U�Q��?9ż?��@?x���!:��X��6)����>�?=��>_Q��Υ��&����?X#1?s��>p�
�������U ? >[?��O��jQ>�&�>��>.-ڽ4Ƈ�QGV�$��{WмK�>�����.�?tB���?���=�?�>�vw>�B��{[��Ұ�>m�[���E��Y�wA
��c����սDM�>�ݽ���>>��ǽi�S��݋�U�������W06?��?A�G?��-?a����������f>LRb>�Z>�=y��=H5�>��>2���I��̾�� ?���?_�?��h?Y�T�5ڿ/Q���SϾ�����> �=�p�=D��[�<Ǖ �
g���;���=���>�Z�>���>�.>AH->�x�=i[����!�G�������>�W�2��55�����6&�㘃�����q��D����n��`U��P��Ò���H��?������s;(?�H�>�?�y�=F�F>�ǫ� IJ�����%�W��s��V�� ����վ3j�������vȾ;#Y��ѫ��_߾�s�>�"���B>�>�>��C==_� ��p�=v������=W�=;=�g<>2G>���>���;�=,>T>ˬ�=�����4��!;�#{V�'�+<	D?��`�ӎ��O{3�ݾ7���{N�>�q?
�Q>;&��r��%�v����>�,3��Mf��xҽ�����><"�>�ݼ=?W�x��n�o��� �=��>�f	>�/��7	�����,�=7N�>���Q`=ÂX>52-?:�p?0�3?�Y�=,��>�I5>�ͤ>}�1>�C�>���>b�>|#?��D?��?D��>g�=�M��DBF<����I����?���4�
)b�$r�;U���Ժ�W�=��>���=�#>@�>h;�bh�x��O��>Q�>? ��>�,�>�$��@4��@�|�	�-�>j�ս(��>Y��>��?6�>Ű�>d?->r^���p��뾮�>��Y><�W�i7p��=]�>�
i>N?��!?��ٽ��T����=^��=�A�>�?E4?;8�>��!>�w�����̿=k'��jF�t����+=�U
=ͬ�؊���e�Vvs��J)��W�ճ1>�&�>v�r>|�=>ڂ��:Ǐ�|_�>��>��">CX>>{�=�*8>
`�=��=xت�=�=��A��H">v���.6)��x���t=�ь��S�<����,Q?�;?�������*~:�[Yg�F��ʗ+?�?�)?�L�>R.徻9���k��Q���A�=df�?��	?�o佋�P��Q=v��=A�$>�Z�>\�;>h�/>�3*�]����c>�Z�>y:?a�?����eG���X�B��h�>[8>���ž?~;?�"����J
D��J��k,�� ?Y��������*�N��:+���#���>���_�@���/?R[�?60�g��T;پ�ױ��E)�V��(��>Ҿ��w�?����!�����Gr���Ҿ�6�:�ʹ>6\?�彈��>��=j<�>�U?�aO?S�)?��H�t*-?څF�%�6?�?�#k?�d?�:_?��A?9*4?_)�����Ԇ��뻇�Ӓ�<�B������=��=Pr�<C)�=�>�R��"�9/K=��u=���=���=>�>�wG>sq?��-?��ֽI��;��f<5��� ��<,��=�Z(>���p�F�J,�<hl[>(� ?�$?8�>U=q���ׅ���Q �n��=[�?��+?�l ?��4=��=WMؾ])|�f=h8>#��<m�p��6���}8����>D��>���=[�>�ue?n%?�]?z�����
�]�$��f'��A����8G�>28>�?�=Z)��1�.�-a��~��U���>8���]&>L-(>(�	>b��>ѧ?>�?�=N+����A������k�=A���;�>���>�.?5
?s3>S��KQ�0�J?�>���m�y��ܾϾ�n�/J >��7>���Q�?��Nр�+K��8�>���>_t�?L��?J�f?�h>�h� �F+R>UeS>�>&>�n<IM�j%C��rg��I=>5�=�*r�	�����<�oS>$~�>�K��U�ʾ�q޾`�b��f���Dg��>Nѱ�yE����'�F˱�&�q>�!����b�!��Bu����q4~��P��cE��A޲�����NY�?q�:?:�?��=+�(�+���{@�`��>�;���<(J�N�c���U��U��s=�N����U��0�3#��>�1�.�������HB��Q%�@��>��8?��ھ�"�����z��=��=kN�������}������]�e?= D?s����
���=�娏=��>��>|�2>_聾���VG�>��>?H�?q�=p䊿^������<���?�n�?�P?��M��h&��վe�c��7r>V��><,?Ǡ���Fp��Ar=��>���>iX�>Z�)��������0�>��r?]�w�*��=��>dw?2�?�g�R�sJ�=�`������>Pġ��^����K:��$�{n>3��>&�>�,���
'�,-�>������ �y���'�Pz���1�=:�?�J��b��>Ek�>g��h% �W���~���ᾼ4�G?޲�?Љl?��`?�پx�*����D4�<Pi�>i�>Q
�>�b�>��1?��S���8��k��nۈ>���?9�@���?�)��ӿ�x����Ծ��Ԛ"<1��s>��3��4V<o����zr��4����	>c�>^ى>��>�1>l�=��<>����"�'��u���Μ��UP��J ��l�B��J�)�*l��	0-�FZv�W�c���?�m	����9V������#���G�T�^>�?�$?ma�>U�,=\8">6�ٽ�i+���u�߂�����U�/C�3d���{��M���q�¾�\��8��Q�����>.��ç?>1Q�>��=_��>VM�>S�t=v�=ҟ�=8U>\�>��=��>�
$>�p>c��>O�>���=+�Y��EJ8������n���K?���b�(�4��H����eq>Q?�*7>+e.����O�m��%�>��|�G�ӕ��tϽGj>�G�>�E=;*%�6w,=�_��	�"�H>!�>�C�=1�=}X��#F5��B�=��>'�r�3��=R�3>5?��l?�aB?���=^�?�=[Ke>�8ý�Q�>1�>u�>�
7?)�L?$,?���>�r�=�h�ϔ���X2=~#"��&o��*7�k~�)Q�=�S�=4�<	$�=*�p=�b������C�=F����͛�����tc	?ؠI?M��>�K�>�e:�.md��|d�mN=7�"=�u#=�?�?���>#�>��>x��;��a�Í��<a���Y�>��=�!E��u[�+⎽���=�w�>3L;?Ob?5��=����`�=Qʉ>��>�?@:?fǽ>���<G��]���W�п�?>��1t������f��x
d��F
��:��N�����vp�X�X=x�>��}>�X�>%�f>���>5���V�>QT'>�.>-��=�q�F@<�Y�;퓃=D>���=��w������,O��%;r�����~ӽg�q�����llJ?�}
?�d���&����/����N��W?kf�=eU?�-?� .>�[¾Z�i�V����r�<�?���?�PN?�&P�6���{h��*��s�-?�޵>�|0>�G��"u��(���yh��P*?���>��!?=C������Z�h�{�Ծ��>q�{< �;�t�?�\?��{��9��=t��]R����ݖ>���¾D�W��nr��s� �H�ze�[$�h�<G ?e��?�T;u�<.��5&�����������Y>�{�=�j?��n=�W�4ھ�s�����Ǌe�uq�>��.?��=�3�>�=Z��>|Bc?�mH?f�9?$+=��-?!����>�C�=7�L?��C?|�?�}?,#?::�>*���~���o�VPX=�	y����;�e�=�� >���;�D>��=]�&�=@B�v�y=�: >�>���= �=\�D>��>�?��#?6z��R>RP�G�;r����o�<]�=
��>���=9�>���>M �>�e"?v�>/�.�ۡ��"��}��9�=�k?W a?���>�د>�p>�l���S��y���'��hԾ��Ɓ��y�NL½�D�>Gޒ>하���>O�?m��>�z?搞�Y�G�*=n�7�ƾbE����(n?�t?)��ik�EA��t4��Pzm�W�2� Z=�M��ڪ=q��m��q�>�/�'c��̩>wk;t����N ��k>�Zf>���>�2B?�U�>%> n��g-���I?󍡾�i��4qо$��M�>�=>�գ?�����}����L=�en�>u��?���?�Dd?(�C�j���\>�V>��>w�0<%�>�����L����3>���=�y�����۠�;�]>8.y>��ɽ��ʾ8(�>xH�?\���u���<�Yо;mо�K��U,��l�� ½�����;��IZ��,Ծ��/�\�꽐oG�$�������}�?7NT?�?���== !��AJ��eD���x=��ԾK����?^��U�_���k�Ծ����+�����^�6��ww�>�[X��+��}�F�(��	���?>{k/?<wƾ]�����2n=M%>���<���J���}����T
���W?_�9?��<���3!ཁ�>T�?cX�>��#>,��W�_�>N$4?��-?��Լ*Ɏ��5��?O��6�?u��?ߜl?5��j>����V��>x��>�?�]�>'�0���4>aս�r?? 7�>��>V����q���P����>�N�?�����?>ӳ�>t�7?�c�d�H�����:�'��<	�>fJ=��ĽZ	J���ͽQR�>;Q�>��f�������[�"?d;�oy�3�N��܆�h�H��F:>��X?�u8�)�>E5>x��>e�N�v�m�YR��L��f�i?cP�?�}?�?��۾B�˾��Ҽ���>r�t>�ٴ<@�z��u�����>Х3>jTپ�����"Ⱦ��?���?��?��q?�h�lѿM���,Gܾ�TѾc��=�H>���<�9��ތ�Vk�*M<��p��#>�O�>�>�\h>-2>6�=�=�2��F�"�����X���R�B�+��IK��	q�~�7��≾�x��o˙�;J���<��,�{|�o$���B�+焽!;����=\#?�˫>��n>��<��=�A]�� ��rx�8����� �J)ƾ����\��Z�g�H�����A�Ӽ���oT?%�-�d�>�&?N�T� h?>��k>�N><���Ď�>�����r;�G>,�>=��=�@�=ypI>�>���=������r�����v^��+j?(�ؾ!򔽃r��,"�6�_�'�>G�?6�>��:���x���>������0�}D^���^I�>�#�>�#�=z->~�6�F�꾹�ս�A�>���>�7>���=���6�b�μ��P�>���@r>�'5>��'?�}t?��7?���=	)�>��L>V��>��>��6>��o>���>{?�=?\R(?.��>;��=u�p��4�=�Ȳ=���^��������&�����(ݐ=�����rͼĂ�<=߻�N	�)��<��?�1?[�>���>�Y�P>c�"Z��� �^��G��=�^?�G:>�?�RB>�D�>�K�;�!Ҿ�V ��;��>s'>��|��Xh��A���Ո>*>�J�?���>��Q�с�=��a�bz7>.0?E?��*?�m?o�M<�Eξ���������$�Y8@���v�[�<��ƾ����l.9��E¾����륾t(Ӻ�\�=��>Rk�>���=�>�=񓻼�%�>��=��@>��<.�<�%��L!P>�6=�$�=��
�t���d=����+�v=}\<�d;�>�=�h�����ak<?�ת>�=*�!��L���������M�>�o�>�ZQ?��I>{y>�~;���2��^�оf?@��?��@?��M�E�9>y�=è�>��=8)�>4V�>;���:�<\�۽AB&>���>�H?=��>O8ݼBe����v�A��a�>d�A=<La����?�X?��.��B�G�Ҍp���_�."�=�	��t%>E"�G~��b�WJ�`�G����#>�)3?�׶?����?�%>�M��F����e�3���v��=G��>s ?$��"�>��"�{*7����c���-=2�?�,�<�\0?�P>��1?�uk?�bH?8�&?e]�SQ=? о�4?�6U=?�a3?�i?;�#?a<	?�J�>6j8��  �!X>�HK��-2����&=�N">>�
>K����=�剽�X6=��-�0�%��#{�꥝;��=�U�=�A>e�=�S?P}+?���Ь6>B����K�����OQ�r�=�}=v<�KU��b��>���>?���>Mi���,�t'�lF ���>D�4?f�H?�2?�����=z�ܾ�`��F�7妼]�=ϴ�=C�k��������>���>rE>h2�>%�w?},?�5/?vC���!�lX���)�ŸN�W��;�ڐ>
H�>D��=Q)Ծ&s&��da�2%i��`/�������F0�=0�=�4�=GV>��=��=���=t�E�:v���랼Y^��͂�>��>�S?f��>���=�ݾ.��7
S?�����������Ң��e���=Cab>���t�?O3?�)ok�+���*D�ٍ�>�!�?��?�lz?ũ轓6��%6>aOr>�>b�����g�jd!�ƽ<�Y>�^6>I��+���r�`<�H>�b>BHڽW�Ͼ�!վ�e�Dy��j拿f|A>w�/��J�&���%  ���}4콶0�����]M�=R-����^<y��=U"�����V춾�
���j�?�C?���>D!=[	�Bݾ"Gƾ��H=7�ԧz�x��\(�=:O�7۾��ľ�	���)��$(��о*��>Z�:��L\�2�X���*�gU��p�>�I?%m���m��'�g*�=B��=�;��:@C�@㟿�}��T(Ž;�?�pY?`���V�,���P�>�#?�  ?!��>�sվ�'��4?E?y�$?�>n���rġ���>Z��?4͸?��O?���ź1�gQr����ɬ?ù
?^�>%�5��`�xy��(?�0?Qu�>���놿s�"�C�>~s?`C��x��>��>��>�����㽹,���Ͼ��������YP=?����Խd`�>	�>�>�(=����/&?Td���^��#��8�˾�������>r?����,=�]>ex�>��@�.M��6�'D���Ѐ?��?T�a?K�8?�S��d�Z�f���>��?�F�=)�>�������>�1���P���*���K?���?�b�?�L�?�^J��_ӿ��)�Ծ�*����=_v�=G41>1��nB����=���d]�S�=��>4؍>Rm>W�F>���=�==�Є�8G#��]���县YR�&f%�t�~ۈ�>�+��m��	��W���
ٽgPݽr[�<kJK��+v�ڤ��ꊾt>->pH?��>ՙ�>��=XH.>Ė��m�"��G���߾��f��;����	Ձ�#Lb�s�^��qu���������9�>I���k�=���>����->�>���=ߝ>'�>4�>��`>L?>4�h>՜t>�@T>Z��=��{>29�=����
���v:�J�Q�c^�;��C?��]��Q��/�3��߾������>:}?�.S>��'��Ô�Y�x�W��>^H�k$b�Ş˽!�_�>$��>�C�=�Ż&��px����R�=Ǜ�>��
>�m��揾�iY�=�:�>�
������~F>��0?[z?�^7?��6>�?���=�ȥ>}p�9��>B��>z�>��+?��7?i�+?���>���=w�:�vWf=�P�=�rN�$o���X��� ˼���%�ϼsq��e��=���=Hf���1*>K��=�)��UA�IjB=��>�<??s��>w��>K{���UM�H�V���ཁa=g��==��>�6�>��>+~�>�-�>߽&=��%�a��-�����>}�L>j�r��C��XY�<�B>U>��`?v~-?��Ѽ�82��$>�g�=}
�>�� ?Y�?���>��=-�	�co�����yA5��Z!�jLý����l��ˉ��ߔ��⃝�}�<�b�ϔ�>���>�9�>l�]=��ջVb��i�>�p�=ܒ>G��<���<�#=\���{��o�'=�t�<��A�r�>^���s�>���G�s�2�$�ݻ--??>��>���4N�=8���S*�V_�<씈>�W�>��m?�]>���\�ؾ�C#��5��֨�*Q�>�p?��K?����R>�hJ>�&�>���<���>lI'>�wp��ʭ�x%ͼ?�=)�>24#?�z�>��#>��N������8��;�>"���3X�?X�=?��X��L��e59�_�v�RX�e�>J&���2�G��^���[��7L��l�"I��<9)���>(&�?)���)�����z���ޗ2���=����=���>� �>��Խ.I྄��ξ�2D�i�=��	?�D��e�?�^��k�>�sk?��A?�&?"$�>�o+?5:�T�>����@]?�5?@K?{�,?�v�>|Z>����콦�,��{<���G]�<�D>���=��L=l6>l�<��=��/�<�J�ب��^�<'�=�>�=j9�=LS>%�	?��.??oֽ�?�=�B�<µ����=�jm<���=![;���s����<�ŋ>V� ?	�'?���>J�;�o�Ҿ�˻��X
>( ?-;?е�>�|�<tϡ=g�Ǿ�L����<F��=�����>��s��򯈾Z߻Ő�>A��>a��'�>�]?L�?���>]Ͼ�M�Ã��U��X^�G�>2�+?�)?B0A��+̾��,�Ai��oaO�F�r�<$=>c�.��x�<a >��I=l��>��x�>�����F�����a�h��#��0X>�M�>�͏�@�Z>JTA>e�%�׺	��p?D�����1���W�$���н� 4>2�>���7�>3y�IJ��&��8�f���M>7F�?�G�?�-�?c-��a����5>�04>Ն�>g�=d����t==����d�>��>]b��=�Y��=��?p�)>����h���ʾP�=�ݵ�p����=�þ��ƾ����,~�� Ⱦl/������U8,�:"��P׾�:S>�ϼ=�����k�{�i
��V�?g��>�?y�G>�3���L�TSӾ =���2�~D����+��Iľo}Ӿ���Z����;���)��
"�>���g逿	�|�(�k��zj>�2?�ϾC�g�]���)=z�=U)�th�'���Վ�rO��Wa?�!J?]�𾴒(��o���=8d?���>a�>��9�R�t��>�-? D8?	�`<�%�����Y|�=ȯ�?�ж?��E?��3��)7��|ξ]�-�?�y?nO�>�1V�mL���ި���?�3?�Ҧ>4A����ZD!���> �b?��n����>'��>br�>�P��e�g�ɽ	����ýlN;=�>=Q�na���;�=�	>.ĝ>��8>���:���>��N�sI�Ŝ����e_<!�?Ut��
>4)h>h�>r�)�t���׉������I?=��?�HT?t{8?����T�KD��y��=���>0}�>s��=\��ɟ�>=��>W�辿;r�̼�n�?��?1>�?2�X?�"n�_�ѿឿUF۾��ƾq+~=��=Q�>?ϽO�,>ϔG�
�۽C���o�>�>Mb�>�ހ>�>	�>
�v>z���*�ʯ��V���0o�/D��K�:�־�P&����%�����~쾎*f=�����aV�����/Ͻq����|��'�=$�#?@�>xў>Kj.>��{=U䎾^���N7�1׾�/ܾvq������J�;찾Ag6�M���#а�;O��b�
?Șܺ�A�=k��>P)f�a8>?�>p��=��(>s�T>�a">i%J>�_>t�I>��->/8>���=��?(�>��c�������v�p�M�e�Q��?`w��y�����ξ�۾�pþ{�	?zF?.l=�]1�������O��>�B�GKq���=��s<Ξ\>E~
?�="� �CJ�,�ؾ���Я#>D.>�<F=�>pt�=^Z:��h��@g�>�g���!���)�>�c?B}�?�<:?Q3�=��+?fP@����>��?��?�/�<=�>�~3?�cF?-�S?u|?���<�Zj��Z�<(�����A�1����罕�>KP=����:��;N�\�����IJ=ae�=R<5#���3����?D�K?V�>�է��;޾��j�#�.�w(r=ĀT�,�>;�>,F?�2>�~ ?�	�>g� ��-޾���i�>1?��>8���гh���C���(>���>�*�?�IF?ă��%%�=����`R>��'?��k?��|?��?�炽����������ѿ$*�����	n�	����ky�H*־�6=�!%<?Mw�xI��3��=J,>* >?�u> ��>K��>���>�R�>�xF>t�>��=L��=9�w����I��=���;L�=�����x=kW(��䦽��|�5�M�) ��Y��}�;, ?}?۞?�`?K�M	a�U��{����3�>c�>d��>P��>��=�����Q��=��W;����>lf?��>��;��[�=�n7�u�;<E0�>��>��>gj���~ۛ�AJ�<t��>��?,؟>���j[�MFk�h�z��>1]V=����?9�?R&�>�0���վ�����z��
O���>Rl=�/U"?��^�y덿����+����[����k�<�%?�p�?9�W������
�oUe�$b&�D6��8s��0�>H��>�}f>G��n��"M���W
�' �}�Ҽ;��>M{�=�w�>;ٌ>\�R?�*s?��I?=2>?S�=%�-?(¾�N�>��>;25?���>��?��>Ț�>�-�>�S>����ϓ�-�˼�V���d>y6>bCY=��^��2�<G,`��V�uw�=��;>C����0=������<�C�=�:>a2?@�L?�ד�q�H=��𼝋���q>*�>6�4=P�>>o>z� ��+�=�
?H�?�4�>�0;��~���
��W��9>�8#?Ŷg?'�'?��>_$=T���w��͖>H�|>��2�۔ܽ�����#��-�2��>�?��A>{q>�\{?��L?��?xҽ�=�&�l�h�$���/��C�=]��>-�>���<Ϝ��FI<�ˑs���V���4��g#�U�X��E�<�� >���=w�>,)�=�>_~�=��}�R_b�L��=�U�=F�>�D�>��?�o>���=�2���E����I?�/���x�Z����<о�C�>�2=>?���?^�
�v�}������=����>�?د�?c6d?��C�h�E�\>V>	�>s�/<��=��,����4>Ű�=�@y�1#���[�;��\>h�x>[Nɽr�ʾ���6H�a�����Z�<��-Ͼ�X��3̾D�ľ�zG���� ��'���uu���W&��eD���/�`h��A���u�늑?2'�?�7�>��:�/��D��I۾���<�����pn��T ��=������ݾ�' �	�5��^;�#vK��j�Rp�>ռW��⑿��|��0)����>�>>S�.?�ƾUr��݄�Y�o=v#>-.�<�3����Ě����vW?�9?/뾪����u�
>?�?a�>Aq&>����C��̓>u3?{�,?My��������X\��p?�?v��?C�@?u�D�itC���Df�B?��?Y��>���4�˾�`ν�
?�E8?��>%������Ê�*�>��Y?~�P��a>���>��>zw�`"���@;�7��B�9��@>�y�����%h��7���=�ʠ>7�p>�O�J9�����>�<�N�N�U�H����>����<��?!��2>�i>A6>O�(����HЉ�q3���L?���?��S?gk8?�X���������^��=��>�ˬ>�ί=<����>T��>�j�)xr���o�?pH�?��?F\Z?��m�׿o!��s��4��<��=�>�R:>�@p�\�>@jS=ꑄ����=B��>�ы>c�M>��~>��>l�}>,8H>$��A�&����V���>�K�Y�������*L��ᒾsh-�j+��v%�����zνM���4B�����;����~p�#�=�S@?�-?卽^'�>��=�6��}��;�p;L��r�O$޾�7�ǡо�N����%8����j�x����x����>�=�Y>�s?�>��=<�>�1P=�ws��aD>�n�>�~I>���=���>��^>��<>��(=��>痨=�B���{��R5���X���C<�F? Y������0� پj���2�>��?q�X>�#��䓿Å|��{�>7�=�;Oq��)ӽ�]鼗ې>�Q�>�1�=ݐ�<�pټ�y�����c�=x�r>�
>�*J<ȋ�[m����=\u�>�J۾�V��S� >F<1?ʱ�?s
�?��>к?$���&��>!<�>�?@��>��>A~/? Z:?�t/?��>���=��{�S#J>bb+>՝��v;�G�W�,�7�$�9$�=�� �_W}=/D��( �ov��l�<9��<��=aB>�??rG?I�>�]P>�����n>�c� ��c>���h�ݻ�J?$f?�n�>��J?pR?��<�cE< y�/EA���>Ml�>v�c��7f�W��=��A>c��>p@J?��5?�&=TFc�k3���=��>Q{??�V?"��>�i>��Ͼ����׿�%�P�"�+Q���:<�Q��1�Q��>���9����ڦ�d]�>*%>���>��>@d�>s�>2� ��$�>�fK>]]:>9w����)8�=�����	=y17���=��)>�lY�c:'�8l��� 但�̽IT���ｾ=�=��)?;�9?���oϾ��=x�;�J��gr�>`�>!''?L6�����Q�բZ��c�3n'���=�y�?�7T?mW��c>���������>c��=�= h|<
�=`״=}��ӱ�>�B?�h>�#�=�����6��[����_>~`=LB���V�?
kw?�h^�}F2�4��<���#�Z���e�:{�=C�g��۾��V��s�%پ��#����d��=8�	?	�?G��>E��7gU�)6���|N��[����U�r��u�>>ż�>۾[���;�<�4���#ڝ>���>�Y�=cœ>��>�?�hj?	�/?�+?<�u���(?S�<�?�X�>�S?66?��?c��>*�>�6�=��U����;쥾Z-޻��K=B�=�2(>�8#>��<)Ì=8�;8�<Ǡ<~,=L��s�����A=r4>��;>a&>X�?Z1?�z�����a�>Y�;�&��>��>���>������YM=�G>-�?��Z?z.+?Ю�>9��0i+�1}ﾻ8'�9�>�~?r��>��t>�L�=��
�\�k�jሽ/�>>���N�s��jҾ0ޭ�f��=�gM>�s�>�n�>�;�>�O?��?�f#?�x+��Q���o�����N���K�`��k�>A��>�&:��ӾA���T~��*Z�v�5���=�)������(�> 1}>f����9n>O >)�<F�9�,��`�=��y>˶�>g�?9b?=�z>rQ>�\���$�O�I?塠�X�� r���Ͼ.���>�=>{� �"u?ݍ
���}�Uݥ�f�<����>Jv�?���?��c?ME���\>�U>�>�-<��?��N�Yd��(�3>��=��y�qA��c�;��[>Sx>�A˽��ʾ�X㾕xF�G溿�E^����k�%��Ǆ��ϾR�����3[��O�����^�Ыk��\R�E��%��S�,��3��٦�����?k?kp�>�F8>��G����?>�/�����Ͼ�踽��E�Je������dK���'��qb�O�P��bѾ:͛>�WY��?��}�|���(�h����E?>�2/?Yƾ�´���L8f=O%>�U�<�Mﾦ������W�
��hW?��9?�?�$-��$�Z�>��?zs�>ڠ%>����콈�>s.4?}�-?N]�_���6������c�?���?ɾ??3�:��SA�J�	������>�C?��>����.��fK
� F?�n3?���>J&�B��\f���>�k^?r�L�q�^>4��>�s�>sn�\ؒ���)�Zl��j?Q��i9>���;�����\�B�kV�=�n�>Ps>5�h�m������>���v�N��H����@����<z�?�L�/�>��g>-�>a�(��+��Fቿ\��V�L?l�?��S?~C8?^��rx�ҷ��؃�=9�>L��>gx�=�-�{Ԟ>^K�>����q���ֈ?"/�?I��?z2Z?ܔm�s�ؿĝ�
J��`�Ծ�p�=�~�=c�m>�Q��.�=J��=F�<Jnc��S>rs�>�.�>�w�>�)>��">�'!>�m��%,�Q���(���A�b������u��f�׾��Ⱦ9&6�K���t��s9���S���Ͻ~;�Ą[��W�0�`���>O2<?9��>d����<>��$��w���D���,��>Z���8�Ss��[��L{վ�؀�2��s!��m�Y2��$��)?}VE>��a>A�>��i��>�?Xg��P��K�d>�>���>�>%�!>��
>��]>\]=>Y��>���>������������3���=rk?L.��3�R6�KR�� �=��,�>N!L?���>n0.�!���f�����>�>�a��x{<ӺܻR��>�v?����$�=G�վ��2�i��I��>��Q>���>%�>����N��ƭ�KP�>�\�����T�>�B?ݒ?%Z�?���>��^?z��>y,?q��>�V�>�9�>/e�>lkV?X�?Ê�?��?3ݔ=�١��� ��B����$����w����O=ZX�=�6>z�q=�Ι;/��������>h��=�>{�`=�x8> X	?��&?�)&?ՙ�>�	Q=���(��BP�ӧ���>޶I>I6?G�?Ҹ�>�P�>&S=�Fɽ����Ʊ���>��=>�X��e�鱕���><��>,80?�('?����k�?ѣ>�4Q�kz�>R{&?;�U?1�>B�i>&6y�����!ҿ^��{�=�o�L�	��ι=�㍽�w�<�Q��ٷ��U����"S>?�>RM�>���>X��>���>Vf>�0�>�A�>��3=���=ee��&¼�j �H��=��򽚰���ۇ<�D+<�F�=�8=U��o�ҽ��=�8=E�л��?�6?��.����Ap��u�:�Y�#����>'��>���>�E���b�=�=B��ߝ����,w5����=(!?ФJ?~����u�=�7��e���?�{�>�b���(s������=�J��!�>K�.?�(=�Q�=�V��L�6���#5>H-o<T�:���?a�u?D���?~羰EE�ИF�Д�?RE�1�/>( �WXM�����!p�/���8�,{
���B<�?�? �/C9>��n��m���J�K�u��s�=B;�k�>�Y�=�{� �6�$W��FP�#g����M>>.?I�>[->`h?��6?b�a?�0?�0"?w���-�>wN�=���>ٵ>,f?�A?m��>|5�>o��>��>�IO��������bK����<P�=j�>f0�>阀=��=q8ּ�C�=����|t��N���ŧf��a�<��=w5>(u�=ES"?=U?�J{��}�Of=�� m>$]��>�[���Uӽ��=,=f>S��>�J?�?�ἆh"��J��0��Z���V[?��g?�(�>�q�y��;��:��犾/o<>Щ�>ccս�΅��|���j�
;��g$>���>ϒ�>dƞ>&\?%�?��=����&��q����T�¾�7�>E%ʽ���=Y�
��P��`��,���d�e�&�e[>���ͪ,�>/�>D�=Ud�=��>Պ�= }�>t��te�<?�;��E�!��>�� ?�%�>��o>��'>d�ƾ��b�I?P����j�頾�jоT+���>��<>�����?�����}��	��eE=�p��>���?��?uAd?@�C��%���\>HV>��>k0<͐>���������3>��=J�y�����D�;_�\>BMy>�ɽR�ʾ4�A}H��q����J��A	�AA��v��h���d���9'���2��vw�i��<�x�8�#��1W�D���ř���۽)C��V_��e��?�	�?&S�>m�3=�FK��Z��7&�F����~@=<�`��V��������'�G���Zc�'BN�u���A�>u>T�y��|�=�'��S��$)8>�.?�}ƾ�ű����b=p�>�D<IJ��#���^���W?��8?t}�wK���N׽�>�?^��>>3%>~��8A/�>�4?X�.?����D=����������?<�?� ??�;��@�Ȣ
��T	����>l�?W�>:c��{��(���	?�J3?��>���j�������>1�\?�uK�$�Y><��>��>y���َ��k��^��4$��
>>��|���b�<+��O�=X��>�x>ǩc�������>�K�h�N�Q�H����G���6�<t�?ȃ�F>6i>�,>�(�����Љ�����L?ȗ�?�S?�k8?}R�����b������=���>gҬ>*��=������>���>�f�yr�S���?�G�?Z��?WZ?��m���ٿ�t������Ҿ�>���=��=!���oT>0C>Ǵ=J�ԽާK>�J�>[k>nu4>��z>_��>��L>�x����_}��7V���E2��/�L; ���Q��������=YP%���ݾ�Ñ�]!�=����������9�a���Ⱦ���<�b�>�v?���><�?>~�=�E��^y���j���6�Gi���4��π������@u�"�c��%k�@\����)#���?|}>�sH>_�?<䋼Yd�=�%i>D�=��&>���=Aw>eN�>@�>��G>q_�<Uk�=�o>�b�>�i�>�f���	H�|�ܾ3�=3��?G��7������@G�-�ƾ���>z�%?c9J=]�T��:��f��	�d>��F�g�Y�d����rF;9�V>>ܷ>	��<	�'��5`���d�R֒�?���o�=��>ʑ�=�Au��SE�����$:>N������؆�>��?��?�E?��-��?���>�[?᳽��>���>���>P9O?75F?��a?p,?Z&>04N�+�=0{�=�A�>7=}��=
J;=��Q��p>$�>8ｽ�m=�[H�~����'W>@'-;��c=�B�=�~?��D?N��>-Q�=J`��z�W���D�l�^>p�+����۰>�$?�{>��>�v�>�GQ��%���'�_{;��>��o>�B��Kzm�!��=�*X>�F%?B�y?w��>��Ē��U&=7W�>�,,?��a?�aP?6a�=(.	=�g侸����ӿ�a-�4�龳�νu+7=ߞ��j�7��N�=�1>~Y�n�y���>{��>Gb�=("�>��m> >u�:>���>�$>��=ŀ�=B'���<=<�q�]X�<�2�$E�<]�Y�N�B�D9C=[On�e���-�b=߃=����s�F��5?g�?a͘�=5}��P��}�	��&����>!g�>�B�>w�>z�= ���W�$H�j[t�?�>��]?���>�u�hr�=@+��>���+�>��{>�>�e�<(�A���m���8��>�?�q�>�ϖ��$[�l�w����[�>)ļ���4:_?��}?h2;��4Y��q�QQ6��+ܾ�NP>�
9=��B-�M�X���i�-푾�+�� Ɂ��~6>ښ?w��?*�j�ؾ%?�������z��^�viǽ�?��>e  ������վk<^�������=�w=��=3�>%?'�?��d?�?Z`?�#�d��>�����>�K�>�.?���>F�>�m>hj>ЄZ>��<
E�ؓ�x�7S��w�=D>i��=��G���`=K��=|��=��m���	��K�%S齐=�P`�%4>f�B>��?�X=?�,<
�/�p��~t���ݹ=��$>e�D����G�о*'ϼ�+�<D��>\4?��<>vTu�����G�-��^V��^�L?�sI?v�?>�I���U��5=���=6�<G��=�[��$�ξ�7�����=v�>k��>��>s�w>Iim?��?��>���=l]&��я�Yj+��lZ�Z�$�@�#>��>Dn0��/�jT�|���
R�Z�J��?�=��r���;w�=Ԑ�=M�=��=>AJ�=ҋZ=kn�<�F����<4�}�["�>ᩐ>,Y�>���=��A>o*콨W⾹�I?���yi��栾rо����>o�<> ���?��4�}�����F=�x��>��?@��?Q>d?{�C��!���\>�NV>@�>�/<S�>����n����3>��=�vy�����Q�;� ]>�Hy>�ɽQ�ʾo2�N�H���˿��d��٭��j�55�������%��/]�֌�=�D�^
��F�'4"�����^᜾~��K��<{���?����?�5?��=#rs>�-�����U{��R��=�i�<O�������炓<A^��Գ���r��b����0�T74�k���K�>g�X�W,����|���(����	�>>&U/?čƾ�������l=�$>(y�<��5��������{�W7W?߾9?�/쾃%��	c�-O>�?:>�>~%>|㓾8�:�>��3?�o-?�-�7���� ���䗼�`�?���?~{A?\C��?�o4�4׽���> f�>ګ�>�h���Ⱦ�Խ?�s?�>��
ၿY�1��%�>I�L?��J��mG> ��>�#�>z󼽲����4�ޏ��b�m�2>Z��R�Mt�� E�o�=2��>��S>W����e�>7����N�v�H��e�jU�끙<%�?�=󾎫>�h>=�>��(�y������
��M?KM�?�R?�$8?���e��m=����=���>Im�>-��=����>	��>�5�jr�:A�Dq?���?|��?��Z?��l�+�ӿ����H���������=4�Y<Y�>>bJX��B>��>�ϥ�=O�=��9>q�>C1{>/�>��=,n]>t�_>�-����"�pA��Hɒ�
yB�((�G���M�0�e5���;q����곾?y����ϤM�.����{��Y)��+d�T�.�	�=�f_?�F#?�i��B��=�|�=����,1��N��d����J� 9r�M���bT����K��9��ϕr�mN�BK?��?>$��>�|�>.�=֒>ʤ=ʋ�=L㻏0�>Cs�>Pb�=�A=Bs�>��>^��>���=�;�>L�>^��W����A�@,K�m����{?¤پ����Pp��Cν�(��Nk<>=&G?�\�>{D�؈�������e>hg����8�
`B���S�Cւ> ��>��)=��V��*���q�!Z��|>�e=���>��>������`���W�>鮧��G����<�g?��?}nm?�Ï>��+?�
#>��S>.˗���>��>��>�+?lp[?|�R?�6?�F:!������;<O>��%�O㮽ۗܽ�&��3>57�=�@i=22=�&�=#�=G�><۫L��$��L϶=X��= ?͆u?�j>���:!-���.�<rU��@���>� ��Ӣ�>7�L?��>Ø�>D��>�ռ8���﮾��߾䡂>�P">kd�Y��r*N=��6?�DB?�Ty?���>
V�=�ɾ����=��>a8,?b�U?��'?b>��i���d)��^,���Ŀ��x��_�����=fl�$B�=�>�����7>Mh�>3c^��?�=wP>8f<>1x>>��>|N�>hq>,;>a�#> Q����<�y½�5Ľ���O��=ZjԽL>ҽ����:�����5Y;�L=$Iy����8?)?�q*?�R;(H�W��{-����|?G�V>"�)?��>�=ED��M���aj�������=JHY?��?��P�U�1>Q���J���@�>Y.�>IZ�=64	=���H�	=�K�!?��$?�O�>:��=�%b�ܢk��`��_�f>��>�*�ڵ�?��}?8�T���(%� �T���P�0�e>${�=� ؾW5���5�Ml��^�"�F��r������b?ų?12����۽P�������������V>��>�u�>/iL=���ml��Z?��f:��'����=[�&?<�>��L>�u�>#?�g?�)?��? �ȼq],?�b�=&O	?RZ�>_7?��?��?Ǫ�>���>J�e>SӤ=7-彂k���U�<�;�<3 :=�O�=+��=4�I�`���0����=��=�����=�=�q�<k�����<�05>��?ҟ]?��٪V�\��<m����w}���M>�.=��Ͼ���1�>~C�>9K�>�P? �?��(���5��A���GW=��T?�_T?O%?F�A�T���xU���z>�zڽU��>�T=B櫽#y������uT��q�>�>�=J>y'j>��d?�|[?�U(?����D��fu�ߗi�dۈ�@D3��??>��;mv�����M�O��[���쁿d�i��"��\�3����z0�>�*B>���ڒ>��>^h=4aӽp��_�"����i�>�T?�:?MB�>�->���8M9��MI?��dz��G����˾}޼!>c�C>���^6?��	�ce|�>ݤ�>����>��?��?b?��G��G�)P>��I>�X>�;�; $�����iK��?*>%F�=��}����n�\�i,R>�w>3ν��þ~ھ`Y�o���iqH��0���'��z��ھ��Ѿ��5�ho������䊾�oy�fn���6���ɽ�����"��Ȋ���6ߕ?��?*H>�2���-C���.��F�G5\<H�ž3��9ǽ��3���뾅ٶ��׾E���3I��q��Y��Gٜ>�GV��n|���(��r��H�:>G�/?��ƾ����,��Yl=�� >�<�<~_�K+��"󚿡O	�גW?��9?��fi��c8��m>ha?��>��%>�<�������L�>F5?�.?�ռI���"��&���	�?�]�?0@?�N��A���G��6�?q"?"_�>����#̾`���d�?د9?w-�>~���l��M(��>B~[?��M�҃b>���>p��>���Ⓘ����i���6��:>Wv&������g��;�&��=�z�>A�x>�}^����%��>h�Ҿ�^I�k)����_�`����=?���"He>wO>i�>]IF�H���8}���PM��4?>@�?N�[?�o:?d��Щ�� ��L�@>>��>P�]>�<���>���>�ڤ�8af�.�d�	?���?���?�]?��J�Z�ۿ����u��^�ܾNM>@پ=8<�>]E��-5=������W=C�LA'�|h�>�*�>c�>[�m>�P�>He>cr���!� ���j싿<,(��{��&��6�އ�e�������Ѧ��ݾ��὆�^����I��]�Խ��� �g�>J.>?�U?;qս4=D>�l�=1������&���c���f1��Z%���n�!��GL����b�,O��W�4����"D�>"<�b>V�>�����6>��>u��n^^=�/>��=ɹ2>T�=�8>�q=�lw>��=�Ã>��=�>��-h��Hk+�ܘ/�./�<߶O?��Z�򹿾�$5��־[z��鼅>)??�J|>o|��Ė��������>�{>�Ig�k� ��1���s�>z��>� >�4=TP��.��x?@�|%T=��> �N>���:/_���潧�:�4�>)[�����>v�,?:��?1�h?�F�=��'?�U>�e?f��;�}v>��>U��>@PY?GK^?X�E?E�?M��=u2/���;�#�;X=�	�!�L��)��t�Z�E��<hR�<gG�1H�<���=�]+��w�=2;��F=��>h�>��P?��>~>�M�
�;L����]7�<_�0���>���>�K?W�>���>ULc>{O�=���������>�\
>��p����y5��җ>z??r��?/�?�Q���x��j�8�F_¼���>�-?��E?ޮ�>�2;�W|�S��adֿ��O�~&�q��=$��=#nf>43���,��ؠ��FU>B�4��b����>6�>��>ؕ4>���>u`�>���>y�%>b�=�D�=������ˠI��u;���U~I=����%>5>$y�=�������#JQ�%��)Ʋ���@?$�>�6���S,=�x۽�>d�k����&C?6'?jL?�Y>��>8I�/����e�]	����>\t?5y@?������=�ˆ���۾�?���>`S{=��ת�|��������F4?��p?���>T���H[/�E�E(�d��=�&>+����?��_?h�7�����z�"��9&��~���)�x�< �������O	��kR�"O��^6��ۄ�ohi>Av#?�x�?�������=�p�����7�[��꘽i��=M�>8i�>���>�\���!1��K��>+���4�e
�>G/?�D�p�>n��>��#?��m?x5;?��:?�]��ۄ?f�Ƚ
��>��Q>jH?�/?�?5V�>{:�>�m>#�t��r�����:���=M�9>�9>[�
>��\<�_+=��<7�=��۽�07�� �=X:s=N=�z@>c�?>,r�>=��>��D?gj�����$3>6�X=�g�=�L�>�m�>K�}�\���/6=!b�>�>��D?�6�>��>�,����I���#�s���C!?e�K?|��>��=�>S>�b3�K�<[\X>��k>�"����V����u��*�\9>E3�>s1�=q�p>�cf?ˁa?�#?w`��ۉ	��3d�*�B�~�־<>�p�>��Y=�a=�4��I0�*YW��O���\��_𽚹f��qA�n_>�>ei���4�>��[>�(I��bԼ*A���=x��
M=)��>T �>Z3�>�ؽ���S�$���I?v����h����oо�1���>��<>��!�?#���}��	��F=����>M��?���?�<d?��C��.�9�\>�JV>>�0/<��>��������g�3>o�=pvy�������;�]>�By>Q�ɽ�ʾ�,�q|H������K��_8�݌��n�z�!@Ⱦ�B��@L��OT�/���щ��g������v�=��:���=��u���!5�e�?��?��>	f<Fd��$;���-��Ģ=)�	��� ����T���hӾ3��{��AA������7�$�����>��W�����.{���(��m��8Q<>+/?�Wľ8'����z�e=��>�U�<U��ޯ��ܗ�����/�W?�A:?������=�>΁	?`��>g`+>�ʏ���ܽO�>�<5?��+?���گ��w���:����?.��?)�O?����,K��1��jh��>^2�>��?\&���Lb�w����`F?s�:?��p>��������}�F�>o�D?�K�����>�|�>ӆ�>�(۽k��H�5�v�������+s9=�4�=���������;��>��> �P><U��ܪ�����>V����H�?}C����Ȉ&�dC�<���> ��{%:>1��>��#>#("��s��Uы��a��P?p_�?�VT?>5?���q��)������=r��> ��>cV�=�,��~�>��>4P�׌i�Q6���X?�	�?�,�?0�V?H�l�JzԿ�ĝ����`O߾"�>8�m>�Ps>n!Խ!��<w�	������ s�NJ�>�=>>��l>$B|>ϒ>��;>�<���W,�,���딿��*���~�ω��,j)��M���*O���뾓����{��d�Ŗ�J����ͷ��3&�kL�����<�}?J?�_R>f�G>��=~I(�.	��FG�{QҾ��7���P��۾� �2���s;~��Ͼ������9�ɾ^-�>�z\��[>B�(?=�E<���=�N>Hʚ>A->gE
>��<���< �P>�S3<�ܟ>�5�>��==A�>�1�>�׏��>��aھ�q2�Ka��I�?���=T���o/�"ķ��kc�rG	�]�$?TV�x[�����À�떖>�2���W��lZ>����s><��>}<E�0v5>�Q>?g����<�P2����>qK�=r]���l�0�ѽ�h�>|?��%
=/RI����>�9?��1?�OQ�8ur>�I�>˃�>Q�>�:�>��>� >��@?p&)?�QH?��?���<�߬�^�^<���+-�����I��RJ�ŷB=����i�3=�=�F|>rW���ļ��<Z��=z6Q����=�  ?A?d�2>��>���Fy��Id��8>�Uջ�#b����>G;>��?-4>ؠ�>6�=����c�	�ǯF�O�>ٲ>U�w�ë���N�>�3N>^����Jk?�I?����ϰ��(�=�7=��>��?N�?D��>ݽ=�t�<��	��޿��H���8�qI�<w��<�w��2��B#��(��rUž.־3���ً���+>%�=6�d<r��<l^,>���>�M>D`K=0�>�Xo<� ����2�/�4>�P=��>���=@9�<�)a�z��=op������	��Z��W�=T$?N��>��c�:�-�L��ѽ� ,��>�2�>_xL?��"?�D�>򬢾`���g���?�C� ?���?�i"?�.F�y�����;���I�>�ш>�C�>%����V̾yH�=Ɯ>�o�>�&?'�>l�z���о]���~�����>+�<z5�u�?jj?��M�Jž7'���&�� ���ؼ�ᇾ�iE���+��F��)��&��E��fR��^m?H/�?�[����=��оI�ȿ�]Y���=��M�=}��n�>�L���욼�;�M
��熾3�k���h��f��h=e>�F�>�n=?|6?Da?� "?��?9��6��>_Ɏ>���>#�>� &?���>@�>�q�>�J�>�>cu�=	ĉ��fb��B��g��-�7�Rq�=P,=-�>D͡>sC�=W\Ͻ�9��^2������<D>��;��6��r�<1��=��?�C)?r�Z��)>h�-�w肾DЮ=��j=ru�=��������L�=�r	?P/?؉�>�$�=�S���i��+����=*D?�~>?	:�>�g�>z��>:!�)J����=��=��.�����������=���>2�&>�_p>Fj> �}?�m>?JH#?٭��h1�pax�j&'��DI������Q�>8V�>�
�=�۾�4�Պt��~`���2��O���E��,�<�q�=��">��4>3~�=��">�J�<�d��<iϽy<����n�>ih�>C?LV>|�=�����A�I?�O���R�%���Ѿe(��T>�=>���d:?V��{�}�8���=����>��?_f�?J�b?uC�D��� ]>˩[>K>�g<��8�+H��ꋽ�0>y*�=r{��蕾ʧ&:E�W>Wt>����n�ɾN��N�8��Ѿ�9U��T����|�������Q��Ծ�˽ З���ξH��cqa��6Ѿ�.>�2>�žL���߾D��x7x?,�c?�.�>�L>&��<s��I־GK���<W��[��qͳ��*->(�=�q[�:p>��Y�:8:�$G侁#�YÜ>��Q�4I����z��&�ٸ���/>�!1?}����o������j=�<">	�j<7p�E܋��K��{��	4U?r�8?u����v˽�>�m?v��>�H>���@wؽ?�>Y[0?YB+?�=��x���V��o�R��Ȼ?��?j�@?W��T0�?�&�:�<���>��?WY�>��L�� ���+}'?5�*?1i�>�����R�(��y�?��s?��&M8>W��>ўh>y���u����۽XA��5������>���=��g�O�����ᗆ�T?�>SF>��6������W�>�$��vN�>�9��/�x�_���3>vF�>�[�@Y�=~��>��4>��,��q��(���℞�V?N?��?z]?	6?�"ƾg�ھ�r��u=~F�>��>��>S��7>N�c>����Z������>ie�?���?-u?g�L��PϿ����T˾�>Ǿ��:>[�=��^>�Lɽ�5�=�=�j=6+b���=��>ͅ�>�#�>1�>>��A>�Z+>t����X+���c�F3-�8i�	����_�O��F�0���۽��ݾ!����;�<�����=�1�1p���R��%�u>� ?}�?i�>�B=AG;>6����A,�s$�q���t)�}<���G��s@�J^�&� ���ξP<��"�н,���W
?�=>�==��>)��<[pK>��>]3>���=��>c�����=��>B^�>��>>p:�>j�p=�{)>���>�`��2������P���
���?g=�8J�@}����4�%�Y�> �>��=m�v�೘��Е�,k>`� >vT�������="�O>�շ>s��<ɠ�=馼7�kO:K���wOJ>���>D�(���D�=v��;_>2��>/B���P>L��><G?z3j?%�?d�C��Q�>~�=3�K>��>Q�>`U�="��Tۘ>D6??�?n��>	=Z����*'=��>�Ɂ�B���ݡ� �&��i��!*�=8��=Rp">�d���>�̠�ȴ3����W=h<�V���v�>�-?�f�>�@�>�D��E�8�����)|�.'S�p�/>8<�>��>;�>Ҍ�>���>9w�>j,�����jmپ�Y�>���=˙{� 3����#�L�>���>�bZ?�?ҒN�'�2:h�>��>惲>d?��?�y�>q��>�:>z

���׿.|��T2�޹�=�_>>�Y=�{9�g���Z�>t�����8�о*}>��?���>=[xg=a��=0�>Mh�=��W>7��=�F���<��Y=�H<�3�w�=�y�C��`9��<N��;�M=W*=�]X=���=�&?T�>�6d�T�Q�G^��쐾�￾>\	=���>U�n>?,��>R��C���U�H�о.y?]a?��?�´�c)=C�r��ޏ�	�>c+=�P���-@>�C��9��݋>(6?{�?-�!>b��<��/�~Zm�!u��8��>9��<�Y��[�?�?�?��+�yЈ�3�׾��2����(l>�D��6�������	��_��5��O־1���ݏ�$�?	ѥ?�t쾌���Ҿ_W���y�0
�p��=ͫ�=z��>$p	>T���>%��Ѯ"�C�žL䴾ΤA�x�	><�>�t�>�_5?3��>5v??�0?��+?�u`�=0�>z5>&��>^ �>�|�>�>ؠ�>��?�C�>�18>.�>M�|�7�|���D>�L�=4�`��k\>�>+>��=�W>�>N��=�"�7�j<�`���Ľ`FG=|�:b=\�Z��<���>9�9?{'O���I�c_*���W��;>S7Y>���gU��ظr����v��>�>8?J�>���>��=Jx��{��8��+=�"B?:�J?�k?8|p=;>��1������A,>�=>��=LK��G�����RD>*��>���=��/>��>�it?D\7?'?�.���'*���a�[.4����=`��>L��>�5�=�Ӿ��.���j��DT��+�vD5�ßC�PU$;]}�=�#�=>*8>�>� 8>���<b�׽\����j����(��`�>Jԥ>�d�>8�m>��=�d��]q��w�I?�����j������tо��|�>��<>����?F����}����I=��~�>~��?���?�@d?r�C�5(�;�\>CV>��>��0<W�>�n��]���a�3>t��=ݙy�����;
]>~My>��ɽ��ʾ�/�ϻH��ſ���J�=��4�&�龁1��R��}t��_�_�	��>C\Ծ��ᾈ�+�Nꀾ)G�>Y�;��Ǿ���AپSҋ?$+?;��>_n >g����	�������<�����Mɾ��
�FI���]�'�k�����+�"�R/9���<���K��g�>�HH�����z����*��vk�Pc>� 2?`�վ@��y����=��=>#
a=���}ꄿ䊔�DH���U?Y36?�y�7�����*>�?s��>k8=>�����(�|q>�0?�4.?n���Ì�$덿x1<�ƺ?���?"�H?-�弘4H�N:���->��>�P>3l�>.��=��󾞮�=��%?*�?��=A��Chs��>x�i�:?jor?;dh��V8=zp�>�΄>�(>��V����������=�[> Zk�<nž�:B����>���>��>�CF�Z���j��>���~}N��pH����Ժ�떏<��?(r��>J�h>�>�{(��������b�l�L?F��?JS?bk8?�����I�N�����=#
�>�\�>t �=��	�솟>��>��bur��+�EW?`�?٭�?�?Z?�Nm�Q�Ϳ������ZȾ�I�=}��=�F>?�@�7-�=�<)������;{�#>��r>T9>��r>�p>�F4>�(>@p����&�sL�������i8�D���"�$Un�ƈ���b�QB��񫾞35��?��l��7s#�����5���¾g�繅A?�r�>M�v>x~`>J�>X�#��ȩ��Oh�x��� ��L׾<�����ӾN����� ����(�ܼ�����
?߉�=�<�>�>4��Z �=�l�>'>�f>��B>	=�y>�>�'Q>NF>s-p>��>�T�>��=w�����5�&�V.O� [�= pO?-M���qz���"��¿�1G���[�>r?�A]>R|��.��Z�g�u]�>3yA�j ��4���=p��>���>��=c�$u��Vt��k,�:�>ǰ�>�?>ĩx=�)_�$���u�=���>�־�=�E���?ᇁ?�$?�!>L��>�?W�>�6��$�<��>3S!?��?x�?�O?��S?&T�=�0����<�j�=�[@�)���F�ؽ�
ý[G��v>���x�3=�Vf=��(�l�S��Pc�.�ͽ�Իp��=8��>��7?�J�>(B�>#&���@�t���Ƕ=po��i��;T(�>�>>��='�>\�>|�<9���jR��	�޾���>~��=9����ȕ�� >��>�h�>�Nr?q��>����}���>��V>�p�>LQF?W?F?_�
?�	�>�i���	��Iʿ����<�狼<QQ�=�����ڑ���>������S����>B{?=��h=���>�5�>|��>㽖=j��>d]=Y�=4t><�����=9_'����=�K�=wbt<�40���<�E�=<��Քa��#=���=�=*�n���?Vh?CS)�ŋ�Q@f����g��Bh�>ia�>��>�Z�>�7�=���L�U�3>A���H���>�;h?A-�>89�;�=p-�lI�: �>�4�>�>��b�a�_���֚<��>;�?<�>9c�cH[�<do�r�
��W�>��IB}����?UW�?��n������"�fj4�B���+ҷ>-�-�񷛾.��0F�K(Q���־ð&�N���Y���?��?�=龪/��xI���Y˿#�������hh��#S�0"�>Q�=�'��ɺ��	��j�F��h�����g%3���->�-�>l�?`�
?޲i?��?�?�ٕ����>�ҫ����>��>�	?j�?ѯ?�4�>�w�>���=�=Z�Z�� ��GR�>��B=e���ҳ%>���=�7�=�o�>�>'�ƼJ���p������<	��=ft2���<��=�P�=�?k�+??ܾ�i��>k�����>���<2�����1�����$3>NEt>�'<?�I@?s�?\�v>�K��m�o����t8+=m�?�-;?`�?n�=|�8��i�?���N�=�=������`Ȱ��~�=�M�>���>�>���>�q?��>in�>��0�7bu�n�}�Zv'�"h��I���E4�>�9?&��p��~ -��n���\z��B\�?ƾ��X�O?0��T�=|�=a�>^@O>�ݥ>�+�(�=*��<���W�9?�<+��>�ò>':A>Q�n>j��@E<��I?����0p�����Xо�+�}>g7=>+E�!�?����}����(=�_��>�|�?���?�-d?K�C�����\>�U>�>{b1<�`>�1Y�J����{3> ��=Hcy�y㕾#�;r]>�y>�ɽ�ʾ(�pH�:EĿ�s��L��B���&��(�,�?���W >�>���g����2*��9>����|����1��F5���ξ�]�?��=?�w�>����/W�3�پ�+��O c>a���t#�l��=R\߽�!���_������߾rH���̾�g����>|Y��8����|�*�(�����:M?>�8/?�hƾhִ�ґ��Zg=�d%>&�<�;�$���*������BW?5�9?AC�+���p�6�>�?�a�>w�%>l$��$��=�>�=4?ؖ-?�Y����4���/���h�?���?L�??��J�ƇB���	�x'��?H/?���>c6��D�ƾ� ��Z
?��7?���>�� ��X��p����>�-\?#�N��a>;L�>m+�>�8��̑�8��x���Q�0���<>4#*���w^��(?��=�=>��>?Uq>�(\�C�����>5�龆�N�2H�������k�<Y�?���>�f>��
>�;)��E��|̉�� �҉K?C-�?��R?Ā8?{������j8��t�=�ä>���>�=�=Px��0�> 	�>��Ws���!�?���?�X�?�sZ?Il�>Gӿ��!��������=%�=��>>��޽�ɭ=��K=�ɘ�)Z=�n�>���>o>D;x>w�T>ϛ<>��.>r�����#��ʤ�4ْ��[B�� ���wg��{	��y�����ȴ���L�������<Г�y�G�^���T>�SVھ����x�)?i��>�S~>i۸>�=Q����>��0���Rj�Е�B\��<۾�����ྩ+��ս����Yͷ=`���q?I��=�R���>i�����=�_�>�=��>\*>41�=��M>��b>0\>b5}>ƒ�>v�p��>�2�>�v��Q���뾇n#���P����?�U�>�IO�c5h�J^A���3�����?��>U�-�/����}��b�>Aؖ���н>Ľ�<U�=�3��L�>kO=u�<�,:�Pe��L1�=#i;=C4�>O�2>yc�:��}�ƾ@���>��5��:==xi&>	�f?$O�?��D?$2�'��=���>X�>���>Dm�>�?(g�>V*?�U�?��I?0E1?���G-m�7#D>�?�=��+����=��y��(����>j�=��L����<�h)>��A�������=U��=ƽV=Kc¼�?a2?��f>P�>���)['��.��NB��U��6Q=�?ĦB=B-?A@?���>��F�^򽠰��o����$�>�l����}������t�=D�>Mq�>��w?�J�>no���9o=��">��]��%�>�qL?474?�P�>�A�>�\> 
�S=ڿ�x*��B�����l�I'>�h����Ft�=���I���ng�>�O=! ->��)>��*>���>�"�>L��>�f�=��=b��=dk���<w=x� ;K7/�Ԗ���K>0O�,���Ѭ=h�q�B|��B�ݽ2�������j�<<?� ?F����AH�O�\����������^�>���>��>��>.��<҂�|/V��?�a><�r��>R�]?�4�>�>��W>����6���>Қ�>h�=�']�����⠾-�A=�s�>��?yҠ>&�潏�_�t`����<V�>�x�<��#��ʐ?_G^?�[3�/�P�1�-�{q&����Y=�=��F�������O�}�>��-о�L �А�c���
?H�?�[�
׎�z������pP"�E*��Ƽ���/��>�
�驾���I�{ެ�2���1<<���>_��=@	�>�z?��?�q?��?��?0NT���>K�>Km�>���>� ?��?7�
?���>��>R��=q�*=�H�����.�={!~��-�=E
>�,>h����f=ֺ�=�!<�;$���(<�Pȼ�ƪ����=�:�=�>z4u=I?[�?u���N��=����m��Ҥ>3�=ᶓ>:Y���c���B���t<�p?��>��?�O�=����G���cF��p�D?� `?���>�s>�Ǽb
"����n�@>��>������+=�(o�Fs#�q
`��B�>|ɢ>=�>�<s>D'z?��@?#CK?τ��^(�Jr��xH�.F��v�Ż��>�EY>)�#>�\����q��t���I�Z�?�`�r�_:�dJs=�V=.��<��t>%%�=}��<P�=��a������{>�����>�)�>��?�=Ǌ��E��ʾu�I?m���5������оT�&���>o�@>�|��y?G�� F~�7����=�9��>��?D��?X�c?�C�����$a>��Q>C�>�a�<S�A�� �%D��o6>�F�=pdx��b��0;ZY\>�A|>_�ͽ��ɾ?�?GG�X����mt��Lc>Az�>X���|G�&E�VbU��3B�e��=�歾���,��vW�T���B�۾����]�½{���P��?�!w?EU>�
�<,-�)���8�
�_.�=|ʾ��|��P�����i-׾)�������/��g�\�KrA�!�<���>��W�w�����z��(�񳥼;�A>x�/?��ž��s�==ȥ>�4F<��ub��%���B�	�3zU?:?R�澨F��p�پ>��?VJ�>z�/>�r��y��C�>�`2?�r)?oX�����l����v��
�?.��?�B@?z�*���I����Z�B��	?�?���>�*��O�����9V�?�)/?���>هξ�A{���)�?t3e?�Ft�_�6>��>�(}>P�ֻ��1���<�Z��nc���=���<&�:���M�8�=w�>0F�>�rY�����\��>!$���N���H�������<c�?*���>@&i>+�>��(�/��yˉ��7� �L?���?ktS?�_8?�+���ﾽY���=%��>��>$}�=Z��C��>���>&h�s}r���j�?5�?V��?�SZ?��m�%~ʿ4,���v��W��.4�=`<>�b>].ؽ5J>��=�zP=v�ȼ>N��>F�F>� E>��E>]�F>��Z>Gg���(�z稿�&��C�<�������c��#���?b�m���ǅ������6T��A���T=�DU��D���F���� >�L?9��>�.�>�(>"�.>󌂾�B���d��C���s�;�����Ѿ�[��r 4���q��]���ӽ�� �P?vr=jX> ��>�c���=�<�>�w�=|#>�3>�>��O>�I->�K/>ܑ>��V>�c>��>Ub�>����б_�o�4��P�`���}�q?�3�Mfc��iJ���پ�$8��n��Z�	?�nB=ӅU�:���=�����>nf����!�"G;��ZŽ �>Ԥ�>��Ľ.�0���=Xž��=�>h"�>���=���o�
 ^�$����>�sA���>�)>��b?(x?H?����>f�>�?�ŧ>k��>�f>\}2>&P??o�R?7�R?~m(?�t	��M��1w>U�S>>�7���=;���פ�@��b�����yr<H�<w�=��>َ�>�
<c?-���=�'?�2?���>>9?H跾4F����<NZ<ߗy�S=6p�>�o=�T�>���>O��=� �=F�?�����ā¾��>~,�=����Փ���x�=�[�>�P?��M?��?O��X�=���=_�->�H\>��?�2-?�??��>b@�=c�Sÿk��49E��.F��ϗ>��;> $����>�%-=?@�-��=2�H>���>��>���=��>�V>A�>Ļ�>T�d=v}�=t��=j�+�9<�8��=��]=,ͪ=����F�*<D��g��<�3��,�<���� ���=g�?]�?�)�;-	8���;�䞾������Z>�u3>�+�>O�?�9�>�Ͼ�hT��XM����?O�u?��?�f�Bgz=�ń<����4�>z��>`N>�ҼmV>�ȥ��0=�ǹ>d�?c�>�[@��]O�cd��7��>�D?=�����?=�f?'?2�����S$��85�������h>j��B���M��$����N������8�eP��đ�<�?v�?��Ͼ��>�fž	%��7.b��<������G���?��)�� ܾ����;��<�P����1D�@�~��">E�>�?qk�>?�W?Z= ?;��>C�����?d��=?�?��?5�?��?;�?t|�>���>�B>�=_ܽ,���j�4=m=�Q&=J�=�
2>�̘=0�A���=��*=�%��a潛\a<
��<O�����=���=]{�=5�?��%?�6)�0�2=����cD��f>&y�<�ܹ�7{U=M�Z��Ŭ�� >���>I��>���>�1�=eʾ �۾���Õ��l?��=?x�?#N#>ڑu����7;��C>U�=��F��=��J ھ|˾a0��?Ѣ>�N�>�D�>�T�>0^t?%�o?�q?�1�m0H�q�1�]����=�[=6�ɼ�����Ck��2�����w�~��%I���\�m���!<8Ҋ>i��=��K>f�=&�W=oO�9�B"�T����>�e,="��>��>��>��>�f ��S����ɾ��I?Zx���m�LҠ��jо) �V�>x3=>F/���?��P�}����ZU=�vy�>�x�?��?�/d?
�C���5]>�
V>�>�3<y>�&�������3>(��=�ry�w���5�;�\>xpy>*�ɽj�ʾ�"��WI��Ҵ�lLb�g
�F���`}��Uڔ����j�
�A����������5���O�ax�"��h½���䷂�Y�K�.:�?���?�� >�E=�7B�^�4�������t�����Н����P�\m��cҾ���)��a8�u ��6*�Ȗ�>��O����3y�Y�(�Kɼ/�T>j�,?��ʾ���x���H=�h.>�=o�쾵���hs��u���U?��6?�%�%y����J|1>+?���>��>Qn��8��&��>g04?�y1?Az���������6�.<�;�?�N�?`k@?�-<�W�D�io�f��� ?��?���>�/��T���k립?��<?�r�>3���f�����nC�>0�Y?P�%�V>���>���>����7r���D�64���y��v3>�@q<yn��b�d3�MR�=w�>ب�>�O�jF�����>�?꾓�N���H�y�����t��<Ǉ?=��;>�i>�6>�(�����Љ� ,���L?���?��S?�j8?�V�� �ȧ�ޥ�=
��>h̬>5��=o����>{��>�c�Zwr����?�H�?��?\Z?��m���޿ ����;��ƾ���=R�=K>�3ڽ�7�=�E=���<4p�����<�|>��X>�ߘ>��>십>QhR>����jv+�@-�������~:�b�����C�v���
�G���,�%���̾9꼾�｣<�s�� �����bFU��,��/���s?�b�>�.>�|?����">��ھ�G��P/���M�\�1��R���ݫ�;�p���ɾԞ<���a=c�Ծ�F�>U�=Vm>���>�U�=;�n>�UO>Ö>,��=��	��h�=�i�;�Y)��Nm>�p�=U.�>Շ�>"��>P��=���zр�y
�0U�k�]��75?2�D�`��h�7��ž<����X�>m?N�>��"�ʾ���u����>��{��:��=�Ͻ��=7�>�e�>Q�C=�*=a�׼*��ڸ��=쏗>��3>�t=�͂���ѽ�6=�@�>Q���ݽ	R�<g��>!�"?
KF?f�c>�;�>h�T>���>���=1o>�dd>�%�>�jI?��a?�}5?	G?��<���������k߽=�n�r�������m>D�ݽ�^����9�\/"�5��[d�g�f��3=}ۗ�X��<�?>߲?��"?��>��>]�J�FZU��?'�AN5�/0��0m�=dd7?#��>)�?B"�>ɟ�>��>��=Uپk�����>�ڒ>glx��0n�d��>Q�>n
">��F?��I?/3��ɉ�ta+='b�>_?"�?�R�?�d�>٧�=�&��nM��ڿ��#�e�.�?.ϽDʼ�xQ=�\{�pWD�5!���7
����Y(?=2`E>��>�!�>�<>��g>F@>C�>W�B>Z�">bh�=	9�;B�=�M
���?>�c�<!Gf=�p�$G�=��3=oy�B��F�:�ٶ1���g�[�0�֊	?i�4?@Ļ|;��1ھ4j+��gG�X��>B�-?��F?L�=�ℾ2SP��熿[m��2͛�����'�?��R?��W�=�}��Z����x�>uѝ>a��=��@�;U���'�=ʦ?~\�>0/k>���=�W�����|�D�U>j=U���F�?��A?��Q���|���%�=�����H����>����� �ç�<�S�1\o�������B�3c��P�>�~ ?>��?�U��!9�o^���N��d�⾌/=�b^>�Y�>*�H>w������iy���ξ���=}�>T�,>=�>�P�>M�[?W�7?�>?>?���p�&?�����>�F?&�2?�==?CJ=?�ͻt��>fv�D��;z�X� �1���)���F�c�{���=��E�r}=H/<�ar�=-s�=�Q�=� =pK껐��=�F=s��=ZE�>k�[=;d?ܺ?H��Sv�=�?w%>�i�%>=$7��+��Z��K轂�V> � ?Z/?ۏ??Щ2>����E�pf�ӧ�l>)?{Q]?2X�=���<	?8w���`"��.*U>a�:��~���D���F��M�Q��>د�=
�{>y{�>]�Z?��(?���>��q���T���~�[S��>G��X>od�>T�>�5��e&��OM� ���m�:�#WT�A�=T�ѩ�@>�"y>b�6>�	��>��e�`���u�@>���> Ă=�M�>��?�2?�=�7�=�Ӿ���E?�����l�jV���̾I�V�"�A>�mJ>(��[�?w���U�t�����G.���>��?[��?��a?ʁ�,����3>b�,>es�=�S�<�I:�-V�I	S=��G>��>��{��y���������=�9>:!����⾠��䧻<�BʿN���O�=2����;�Oɼwݞ���;>CQ�;��` �f�`�8����`p��6��P�+��J��6
n�s|�EȜ?��s?�W?KP	>U�.��o�6�`�0��됾@��������X=
�Y�Ⱦ#y�����g�T��/)�`s:����>�Y�w@��R�|���(�����Gu?>�4/?9_ƾ_ɴ����g=CX%>�l�<�?��������%
��aW?�9?�K��(��c*��>��?�r�>��%>�#���*�q&�>�84?��-?�$켂���9��D����l�? �?��??�N���A�>��3v��?rK?{�>勾Ug̾a��1$?_�9?�ͼ>R��+#�������>�Z?�O�Xv`>ȝ�>�>��������r��
���^��58>��ʻ?�a,g�G�=�P �=��>��|>�_�����S�=���pn�0un�4]E�9tѾ�:>�!?N���_p����>��I�����?��Ӡ�A(��sd?���?N@P? ��>f����оT͐�A]��&(>_^�>4%�=����>P��>]p��H�e���پ�X�>y[�? �?��9?,sj��uʿ�4���Tþ�h��go�=R�m=��\>�����h=C8�<27�<xGļ��*>��>�<>��>�ă>X�w>@�X>�����
"�:��-���2�]���)�$��CJ���y�� �<���⽾y�,�̩M�)��K6;��ս-�s�u����l>/�4?��'?{\,>Z��>7KW>Դ���w������9�h�7�j_�(Ҁ�I#��������������J�J�ƽ;q�����>����pT=���>̒�=���=��>�t���l.=ܑ4>×>4�U>�LN>��>�>�=��>�.=��>�>����o��gؾ�p'�ra`��"? y��	b�/8�Q^ᾫԖ��¸>�q"?��=��{f��i��v�>�5��������5�>��>��>%�E�U��<ubm<oG����ᗽ�]�>�>Db�V�>���0�S�T>�o�>B�Ծ�3= �.="  ?�i?�7Q?�[�>*e�>x�>�	?ѽ.>s?��{=%�t>�Z?�gz?f�V?#&/?0�<��ɾ�����/�z��.�g;�jF����=����=�>I�>K�>ߊ+=�֑<:M:GUE>�ʟ=���;�{�>YE?+L�>�>�>�}j����K�P�!�0o�=<_P=ZN�>��">�*?<�>��>Ի�>��u�%��1�(��<�>�l>��@�}��K>a��;faӽ�.7?��)?ŪҼ��������:�=�S�>�t?}?�d�>߷�!
>�g	�ѿ
�*��*��h�� *���E>����hh���=w���7��*>����C��>X��>wć>�h�>d�>�>8a	>8l=�m�=r��<L����<0�=���BQ���:=Ž�;�Q��cs<x\�5-��mh�� =vN?@?(P�<�Yb=²�#W޾`���� >�`�>�u�>7 ?#��=p��M�I���7��91��?��E?���>�=��W=Z�w=�|6=�C�>3p�>)n>���Tg�����~}���>�(?�+>��Y�`�B�m�x�,��G��>_=�Ჽ9~�?�46?�N�)]¾@J�z� ��9�Ȱ)>|��)N��Qأ����k>��	���
퐾��=�\t�>Ƭ�?��o�ؕ;>3̓����)`��n���5��=� �F ?��m�������*�(��đ�	��M��x\ͼg5�=��>�?�z?
RP?D�?Ϥ�>n�@���?L�=+d�>B��>{z?�+
?Y^?6��>}K>�")<|8������J��b��<b=�<�Ǯ=5N%>lX>\m=��K=u�r=$��<b�Q��<��������=��=�Y�=�3>;?PR?a�8�K>L��>E�#9Z=`����~�F>�c�=i� ��J>�'���e%?��#?gN(>f����v�pe־乪��ۺ��'?�}6?�l�=V��/_�>ޅi�䒨�47V>S�|>��(>3��sU�4wϾ0R�Qt�>�r�>�.O>�1V>�{b?Ie@?H?ڛ���Z�L��pU��<��i���y��>�Q>����4��G��N�_��p�ӳ��o���F'��74>�->���=�OC>ð�>�o)>3�'�F��>y<���[��0��>�}�>/^#?@�}>T�g;�6��V�d�I?����7��^����jϾ�9!��>#�>>-��e�?���F}�?���=����>;��?P��?v#d?��?�����X>$Q>Cn>�e< �:�'�p�}���0>Z��=g�y��������;D�Y>NNq>��˽͊Ⱦ��$�9��a��z���ۗA��b*�d�Ⱦ�羰>�����>�qľ����-����̯���9��L�d�̍�s�I�IՀ=%y�,]�?;5o?~5>%�����OоX�ﾗ�>$b����:"��]��;�O ��u�hv/�s`W�8�Y�Zv:>�ľډ�����%��lb;/�e>�L?o����0?��>6ϖ=Ώ�=r�Ѿ�ǆ��o���¼��Q?�JK?��t����½}\�=��?�~�>^6>��ƾǙ���>��G?��'?�s�={h��`������?���?(�I?9"��lR�����N'=`H ?l�>]�>��~��1���I˽P1?o�?ռ�>tӾ-Ƈ�y��0��>�m9?t�1��>�d�>�^�>L�?�W������;�P�"ލ�C��=��b=���l@���|�M��;���>�Q>b
y���¾��>�A�I�N���H�{���v�͈�<T�?Hp��R>|�h>W�>_�(�����É������L?C��?��S?hW8?pp��$�~�����=Ѧ>	��>�Ѯ=}���>���>/B辩,r�}��?�G�?,��?EZ?ǖm���ӿ�6��ޤ;�۾`u=?��=���>h������=�Ճ��ڒ��:�<�\6=��>�T>�K>fK>(|v>E�>ٙ����&����{���]E���'�׾࠽�۾L�����o׾�� �J�-���C���箾�n���d�<�;�����=�?�\�>��>g��>r�|>�A��Jɾ�ꌾ��ҾB��*)�:z�"��u2������c�N�p�J=���'?�E>�Ⱥ<L%?d��<�+{>�;�9�<|���>�=e(=�h�>�m_=�Ž��#>��b>��~>�=N��m���� 8�*VI�/ݕ:�*A?@�Z�󉔾lf1�^0߾m���M=�>e�?h+T>q1%��ʓ�6:x����>��B��b�!ͽ��
��=�>���>ݎ�=^���K!���s������=?\�>5�>u˙�k*�����T�=2��>�(����þ$Ko��L=?;>P?##?"��>4k>�	K>�>5�پ�R�>!	<�T�>. ]?4�L?�t?��A?B��_χ��bu��=<TʽNe�:���1
�;�"�=ԯv� h����=_��=H|�<�^=�~�=�&�X?T��8P��?��>?�)�>�2�>N��A��T"l��I��dD;>�5�>�J�>���>�@"?2;|>�<�>��o>*]����Jc��;��>�@�>�mf��s��b%)�,�4>��[>�H:?��>?��=T~>�J���%����>���>l]?��G?�B�>8~������	�Z�&�P7��KϾ�k���L>�W2>��4<��l��N2=<RC�99=���=�σ=,�V>�m]�3�F>:�>w��> 6[>�]�=�=�C8�Á���:�g�I����;.�>{X�=�]>�l>#W���|�`I<֓�)8�1I��?�?�PۻuΚ�t^�u��aX���w�>�S�>�?E�#?X��ص��������y��)?�hQ?X#?!��t��),q��p��@�>�f�>��J>\i�=�[��kA��D�!�;�>�?U��>~���h�f���i�+S����>�<�ｭ^�?��>?��(�uS��?�G������|�*��>�m���Ͻ��Ƚ�J��Y=��T,�m9W�O2��/�xB?h!�?<��Y5��^L�X��n4��Թ��������z+?��P>J_>����i��v�־F��Cյ=����lj>���>�~T?}YX?�l�><"?c�>~�&lF?z慨����N?��=e�
?u�&?m@:���<c�K��:6��l߽\�.��Ύ=K����>�٤=��=u���z�=�\>).
>��=�%��$(��{>�.G>���=�7<;ɵ�=�~?J�;?�S���m<��=��ʽ�^O=�j���[>��=&�j��=�K9x�?�y?��|>�=*>����i �L;��r�;��?�?�3>nʠ:æ>�����ɽ}ϼM�='"�������f˙���Խj=D>m�o>���>x�m>�wm?k,?��?^O��:�8��e�r�P�w7a����S5���p�>���=�K'�6�/�?�e���O�6p�����?�*���s�rR�>�g>�G>$��>h�>����kr=vEE<d����}5>�|>^D�>�?�O>��}��UӾX��)"A?9������E�h�R���߽i�9>�p�>�E=`P?�L�=�����j����/�?�?1��?s�c?��컝?���6>Z�>i�=����'"I�O~��2��=hA�=��>��V�̅�a�5=�[�>\2>���ӽ��K�a�P=�l���`f�-+T�l�⣾N㾞\����˝�C����D�@����Z�������̾��*���Q��S��_^��Uˌ?4.�?C=�>Tw�=�6׾y�������XN>)Õ�6ȶ����FG���,�������4���
����Z"쾍|�>��Y��L���x{� �'��ͅ��?>|E.?
ƾ�W��t��.m=��>�ޒ<U��z���kD���.�}�V?�9?K��8�����۽Ѷ>�?��>7'>֪��������>L3?-{,?w��35��큌���Ƽ(*�?���?6�I?���;�e�����Ж�>^�?���>2�>=×��W�I�m�x�??��1?3\?[���O�v��޾Ǵ>�>��#�հs<���>�?�x����>U�=�-��޽T.�=��<Rɽ�A���$<�0&���/>C+F>��&�r,�����>�A���N���H������O�<��?'��6>Fi> A>��(�����ω�~+�D�L?���?Z�S?;l8?�]��������k��=/��>�Ѭ>@��=�����>���>�e辯wr���v�?�J�?��?�[Z?ڙm��%ɿ�h��qk߾�[��Y�J���Y=���>|P�n�+>�C=׬�=���[�<�٨>�.t>� �>��>�2�=�H>�t��C�'��A���#���+y��.���|b��
��p�ݾF��X��ü�~B=p �<���Ӿ�4��\ؾ���[/?���>�d�>���>F-q>���?��=����������l�?����{����{��<���X�Pj�=M��!�?��/=ф�<���>��N�9�>a��=V��=U�1=x�f>^��>���=�:�=�6�=_���i>��=��;�tG��%蜿�M���^O��=��0W>3�&?��<-B��r���PC�I�"�KV�>]qO?�6	?d�ྪy����<��>��Z�GMQ�|	�o�R>P��>���>��z<�9ҽ
�9��}y��3�z���*�=�y>n�=K!%���!�vz.�*��>������=B+�>8u)?�y?��>?~���:#�>ȝ>]�>Ԣ�=�j>$�>Z�>�5?��@?~9?�C�>Ky=��S��
�=�ʔ=s�,����ɼD��;J2���=S�I�l+���h*=&� =׏�;�gw<A���7v=��>N+?1�)?���>3uY>O.q�{�i���U���=��p>�F>�u�>^)?�?�-~>��e>Oy�=w붾���}����>8U�>��v��[����b>|> �<_y�?�/T?D����2Y��3^>]�>Cz�>�.?قJ?�μ#�9>���I�#�ο"�'�[~,��L�>�;)*�=����X=ԉ=��?��K��������C>zf�>F�>�ۆ>+&>+�>S�>���>�<W>�@�=bq>��>��L[Q=7�5�]��3i��DL�����|��Џ?�Jڻ��ɽ.���1����?�?�����؍���|��H�i�ľU.�>�g�>>��>���>(�=T���)�V�_�B��d���>Ca?�!�>�C��>=��}��4�=|7�>�{�>7|J>�ɽ��-��ݟ����{ʸ>�9?Q2v>��(��Be���c�|7�DΩ>��[=�����?iZ2?a��ဓ�˱,�v��OQ���>ǇP�F��I�ɽ�W�םS�{+����b�î>xO?�:�?��Ⱦsf
<�"��f8��=�r��Ū����<���>>?�q�>�t�=�������'�����`+D�"��>ѷx>�?��>G�^?MsS?�F?�:!?�q��D?�/��:Ů>���>r?�??�%?Z��>o�?��^>[�����4�0��=���:$ݽ�z�=��{>�̽e�.>��|=1Ϝ=�?�aٽ<y"ٽ�-===7>��J>��=�{�>�,?#(?�Y]����+�>N0�:�f����>yI4=���������#>��t>3�?�?ڡ>#�H�ȍ�u7D���� ��Y�?�\?z��>()>p�i>���p������=��j>��;+%x�� L�s�ξ�Á���>T�>��>bK�>�Fb?�3?z�>侅�G�W��f��Q����D�:ʗ>�հ>=/?�֪=v
�'�E�?�����B��f%�cc�<v��Y`�g.>�(>�xA=%�e=�T>�t="�1�`��ai�<ѷѽ�m>�O�>�a>P�,=+u�=�W�%�ľ��I?r����j�R1sо�J���>��<>����?H��:�}�����G=�ˍ�>S��?3��?�>d?;�C��)���\><MV>��>|*/<�>�����J�3>��=l|y����E)�;�]>`Ey>�ɽ��ʾ%2�H�UT����X��ν��Ͼw�s�ߟ��\x�}�R�FF��3�mؾՎ��1��[.���1��r1�]�Z���怾���?`�v?%�=>3�:<�M�=�Uʾ�,�=GL��r�%�ʾ�=A��K����ݾ�ѯ������3�^�$�&��ݛ>��X� ��+�|�o�(�!����/>>K/?�Wƾ'������4j=X�%>�:�<yR�x���/�����
��W?�9?B��C���k�ݽsL>з?9��>�$>�e���v���>��3?)a-?Bp��<��hJ��$����W�?%��?C?�#'�/�?����z����I?��?��>�M�Ҿ�8���G?.87?7�>(����~���$�?�D?�cW���N>�A�>"��>+ڽ?(����/:�N�����2OF>�`�;Ѐ�<�A��a���=@�>�t�> �]��c��ƕ>q����T��N�.�׽��=�Z�>B ιУ=�W>wO)>���鋿�ً��0нf?V?zA�?�3M?\g7?|��`'�Z����#+=_�>�>`�-=,~2�T0�>���>��о]�`��<�գ�>?��?�?�?9P?�u��>̿K^��.E��?R��M�=-��=a�W>�go�v��=.j�<Ƚ�;�_��/"�=Iޖ>|4q>E�_>��>��A>��j>���[D+�U���4��{�M�[9����V�)�b��O���t��7���u׾C�����WCC���R�z�$�=@8�B�˾��I�n��>�~�>��>�?X�.>u��������Z�����S�7�Ǿ���h��G�`?{�sb�����<f$��'?t��}*
>)�>Ƽ���>�i->
q��$���Ä=���>]�>&��>��k>�<׽��=�+���r�>s�=>�5~�g ������|P���;�'?�	���v�+�2���mPھ�)�>e�
?�p�=��&�p���z�����>��!j��V���h��=�.�>6�>r���Č=���ѧ���z0�@�=�!�>��O>|��=U����/����=�d�>��q{��;6=R?��Q?�G?�n�>r��>j;�=O*�>aR�=ء�>_ʃ>]��>8u�>9�;?��^?�$4?�I�=�Ѿ1���ְ�!l2�XƯ=���m��=�5t=v>B0ʽy��;*�>�+���`V�sh"�/	�=,�޽B����� ?J,G?g�>��a>hT�,�V�iA'��l)<�`;=�Jq�'��>x
�>��>�3�>	�?��<JZýɉH�=,J���>�EU>ǆ�|��� ��=r�=SH>��s?�Z?�����ֽi�$>��!���>@s?�ɴ>J��>x��>N�����\P�ȴ[�F<B����TQ�Ul�>w@��>>�̃��ҋ�ה�;KW>��<T���Ƣ>�Q?鰬>��Z>B'�>�b�>K�
� ��=oI��p��=��n=�n+�g?��i�Ĝ=O�>at�=����h����)>�n	>J�v=�i��aM?�??k4��^��z�f�����u�����> ��>h��>�s�>BЪ=������M��?:���C���>r�m?h�?f�9�:Q�=�(��ࣞ��F�>u+�>,
>?W@��^�̤���m�;`��>ӑ?��>k�&�A�Z��Tj����r�>�f#=u����Hx?27?���a¾H5��R���%��p6>�]��8b得��R���H�o��*�R������\��b?F��?���&Y=k�þp��� ���[��-F�G�>��??�5?3p��x��:��8ľ�ґ�����W�>�	�>2q�>��"?�1?�NI?h��>}��>�nѾ��0?�B=�y�>���>:.=�2?��!?�R"?zRL>����W|�G�V�4*"��g8=+���d�iw�=�6�=�mt��N�=�u$�`��=��=(�>6f|>}rb=�|�9->�KM=i�7>#�?Y�"?�v:=���=��A>bs�
	�=򈺽A3m>��=���h��=F2���M(?H�A?P|�>w
�=�ܱ��Ѿh`�-�/���D?��V?
^�=��ļt	�>�1��®q>�^̽�Z>UG����g�u���@�q>�L">��>{5�>�N>�O?��?,�?��Խ�9-�����H�C��5���?pT�>;4�>��':�!N��p��o�[py���U��z�__�ϖ�W�V>e~:>�qy>��f>b�>bК<��O����b"��V�s(^�~�`>I	?)��=�2">�w��@l�d�I?�`��Y2�S����gо�1 ��,>��<>����?�n���}�|���'=���>�?z��?=.d?V�C�vo��\>w�V>�1>,�(<}>�B�UH���e4>���=ˍy��(����;e&\>��x>�cȽT�ʾk��(H�����bz������˾?��� ��=,�ֽX>�[a�Zx9�&�i�Rʺ��c��ȾYG�CS���W6�mv��5�?�cx?9i�> �:=�H��Ʈ�t���s�=���9\g<��Ⱦ������̚��\�*�)�X+d�q=3���� ��>��X�2����|��(�AA����@>�J/?��ž����#��l=��%>�M�<�+�p~���h���t�ܞW?0�9?�E�p������>P�?���>�x'>N��K��E�>f�3?�7-?���x���=���|��3\�?3��?L�<?������(��'���%����>�.?�n?��?��M���;Nv??r4?�@�>�����r��[���!?��?*�;��a�=գ>�2f>�Qѽ-JO�x��g�%��=c��>�'���m�r�%�ʗ���f齴�>9�>�a���r��o�>���_%�J!����#�ž�KڽH ?]�ƾ���>5�~=YK:=�o6������T���ҽ�P:??@�?�I?:?�h����$�E�*2����=���>���>l�!�`">.X�>+q"��	~�Ν�_NG?`��?�t�?��\?Ak��'ο�����ٮ�LU��)B>��>�DZ>Ĕ���l>���=a�;�S=_{B>���>-*�>�u>��<>��:>d�6>r&����(��ğ�``���0�^�WS�O�j�(�R�Q����� ��H�����U���0�$	3��X����<����[��=�*<?o�>.u>6>0a>,p��(�
�+����ӅA�]ƭ�AW��c�������?a��ؾb3�j���>+��u�>x)��T�=���>�ҕ���l>}͇<�wb>~�=A~�=�ּ=~�x>i�=6>�8x>�U�>�)~>F�>��>ŋ��U邿f+J��[Z���o�dzD?Bi&�y0ɾ(k�}��Y�@0�>u�'?���>d�����M%P�i��>k�� ���r��:�нL��>$��>�l��[t=!�������@�\�>"��>��>�I-=Z����yC��_�=m�>C�߾�=!�t>�?�~s?�6?g, >Җ>
�>8R|>;J�=��o>y(> �u>/W?��A?��1?1��>1^�=|L���_�ذ7�e,ܽ�#-�u�콈�<fmU=��0=fU;���=2ĵ=��=�}<�t<�M�\j=��A='��>m�0?��>b�>'���� U�/6>�����j�=�"�8Ӝ>\�>Q��>l��>��>�q>��=sؒ�x;ڀ�>j>->'�y�z������>�Ŋ>6�[?v?Y������#��E=q�>�(%?>�A?O��>~�=����&�>f�Xm��$<��>�tA>�'�>���;Bq�=}�$���� �<�rb>�`�>?d�>��7>Fe�>��>���>��s>��=Fj�=��� �&��pg�W�<�Mi=À���ؽ!������Ъ����Ľ�M���'�;�X��M��"�1?ٔ?J+����=17��b)���CɾHM�>x5>f6?�?zj�����8��UT�$�����>U�v?n�?�Fk�6g>����<��m%? �=[G:�w��<+%�=XL�5�>���>=?Oc�>�q��c�[����������>sU��$�N�>��?)^,?ȱھ`�^�3Q�w�I��� ��h�>��F�,�ͼͥ۾�o,��'Y���Bl�l������==?�Ԗ?���{�p>6�{v��Zm�����8�>�d>�t�>�=J�]f��������I���L���>��?��,=;GM> ?�Ą>�e�?��Z?��A?�9�;P�3?<{��I�> �?��b?��)?�?eom>�UV>��>����s��B���U�<�,����=�L0>��%>ɑ�=���<T�w=~<�*׽�M���=�1�=.��=f->��>�#>��?�(?�꾐�9>Z���ᅠ��/5>���=�O=Aپ�3�b�;9C�� �> 
/?�#?�&�>N���˷���޾� ��?Gy�?�3�>�����>z���];޷^>%F��=Vx>;T<�2-����i@ɾ���>n��>�b-��"y>7��?Ի?��?].>�x���kZ��%�~��>/:#�+:?��>��*>�s澀>�i��� ���8�>o,>�U���>����>.��=_hp>�DH>���>U�=�����]c���V���j>:��>�J<>�]�>Cڇ>���<��̾�-�7�H?K�I�c	!��7������uL�	�>��>UZp��
�>�a6�&���ˠ�6� ��>�I�?1g�?��K?����V����9>���$;ؽ՘D�W�=�A���Cu��	z>�{c�8�
���ľ�;�F�>�4�>\��=�T����޾�Br=8����kC��NS=�ҾY��L〾������x�.^���g��4;����X걽?�=>8_��7��Rо�Aؾ�<��-�?K��?A�>�Nݼ�l8��(���*��7�3��[��ĥ���\%=^�о�jɾ��ᾳ0�,�L��a�TFJ�鿛>d�Y�@��I�|�u�(�-���?>5/?PcƾR̴�	��`�g=�_%><�;�ή��{������aW?&�9?�P�-+���὏�>^�?Gq�>��%>�'��2�x(�>�84?�-?�m�����9�������l�?4�?��??��M��A�������?<�
?���>:��˾���3�
?§9?��>f��]��~���G�>�[?��N��xc>���>ٖ>� ��o���'*����^'d�)j7>��ۻ(�h���=�(��=�ߟ>nu>��]�ؓ��{��>�0��y�.��;�2���I����Ž��?ل��;p>�Y�>@d	>�$8�Wێ�F���|����O?���?�9D?�LA?"�������c��=!�>
�`>d��=2o�<4�>i�]>���O`b���ξ�+?mK�?�{�?%�G?�\�>Gӿ��!������	��=%�=��>>��޽�ɭ=��K=�ɘ�4Z=�n�>���>o>D;x>w�T>ϛ<>��.>r�����#��ʤ�4ْ��[B�� ���wg��{	��y�����ȴ���L�������<Г�z�G�^���T>����}�?�7(?S��>�?��">z|?�P�;o^>=�u�����b�-�"�h�7�W���%L�w��P��;�ξ�о�����)?�%j<U�l>�,�>=aA<cn�=
�o>{�>��E>��|>�E�=�J=e
<�	�=���}P<p$��Z>�
>pӄ�����e�4��]'�����+�?p̽�=���lK��򾕫��v��>O*?�&�>�� �������P��>н}�����ɽ� ���>P��>�ߢ<�������bg�^⋽��>���>��K>�]�2���W�ȽB҄>���>	8־M��=���>�?�vh?
�(?@������>qR>`ɂ>B�=+�t>��t>���>5�?�m:?��/?�� ?�J�=�*q��o=�#=�K��b
�������l�M�;���@\Z=t̽=�j�<S{�=qq�<"M�f�<�򅺎��>R�?}�>BF�>e뎾%C��OR���(�~%�=�����>!p�>��>d��>�d�>��%>��=q{�Q�þ�d�>�>�*m���r����=$&�>~nd>r�D?��?G�d�4�����=;��=�e�>&k?|$?ታ>S>��'���Ōڿ%�ʹ� �P�m=��=�A3��냻�O=�����ӽ�e+=3C>�C�>m��>݁>i>�g3>��>|�>bz�=n�=/�>��M;�Y����}<�ћ���<�1�?W;�R3�.꽘���ؿ��3��՞v�!��io?�n?���l��X����K̞�fd�>Q�>��>�^�> ��=�x���T�]�?��>?�&��>�d?QN�>�F���=���j����>O^�>"Q>AA��)�����=�<�>qh?w��>����Z��p�a�
��o�>����+�p-�?�\??��	�^����=#�W3+�W�-����>+q>t�޾7�0���j��M�I*�Bz����]<�?j��?�(����<��ɾ�������7��n�>�ͱ=��>p�>�7���ؽ����hu��ES2=�v`>�U�>�;,�c�^>�$1?�+?�z?��,?�z(?���E�?=�^>p�%?���>l��>�@�>���>�F�>z6�>Qo����	D��Ï��Y���7���Mf=%�>7��=X��7:v<���=�V�=>�"=�p<�Z;=q:i=�H= �s=�->�s>�K?�>?��Ⱦ<�x=,����W=Jν�^�S|���M��ؘ�~����ט>k�?9�H?��>?��>���`��=q����=�|"?�Z?�J�=�HR�Fҕ>�D��ײ��=�,�>��s������y�;���[�Z���m>���>Z0�'G>�O�?0�C?�T?6���F)�I�T�g���c=�D�;�F�>�`�>���;B��:���j�N�a��0�c�}��Qp�5<�&2>�>��Y>�t�=�2>��;=u
��������=��<�!�>�s�>\��>V(4>s�<wSƾ�����-?��qa���쾝�ž��-��.���=��<���>Ղ��s�lc���h)�T�>���?d��?,/?��<�L�<�5!>�A����j�3‼�>+��ㅮ�K�>�����о�!���(�=��?EG
?BHl=�sӾw���=��˿|�M�l�K>똾 !��L��T���u4��Y�^B>��4�����zBb�.Տ�ꈾ�#�5����
�x���c �?��c?�>p����8��D �i�	���=v��5~=F���[�� ��}���M�վw2�5z,����H���m�>Tp�������D��&;�0A=WC�<I&�>_�����ž���F�=U��>&k>�Z��&~���g<�&L?ی;?���3���<C�����>�9�>�L�>��>�k���q�E�>��\?A�7?�qD�C�� ��� A����?��?��g?{�����]����Yu�;Ӟ�>|`�>�}$?�����P��\��eG?�LT?k)?=�ݽsχ�z2���B?k?��W�^�b>���=k��^��<�[�ky=>獻��~>���>�����qgվw�g���5>x��>|�K>��Ͼ���S��>t��:A�_�E�%���X/���׻m�>�m�X>F}O>��=B.��u��?x����#�F?�8�?�2Q?h<?mR�����S��@Q�<о�>l�>�oY=@����>Q�>%��X�g�����?�B�?"��?M�\?��d�(rӿ馚�{��n��0FA>�ˌ>�nr>��:��X>��=vc��<>��l�=>s�>�5�>�7�>�nh>]\�>nU�>9W���P)�3ω������"�ۊ㾰
��c�{ ���P��K ������O����'�z;F
=�s���ͼ���=̿�x ?e-?�g?��?^�>�"�>�^=��
�<�����&G�a(����\�����mĸ��H������?ڽ����x޷>�.����>���>W��=��>xE�>��=�H>QC[>;S�<_�.>|�=��Y=weH<���g\=���>�潇ӏ��U���O=�{I���|c�e��>����M�ͽ3I�=�~<�C�Biv>��'>��?�a������o�k��>^$�=< _������y>g�?�'�>�[>>�EP��e�"ܽ����|<T
>��<�]	>E�+�m	��IdO=%�>[������=~��=i�*?.�x? ]0?Xk4>=�>�v{>���>��=/�&>>��>kr ?&�0?�%?��>���=N
V�>��<�=9!3��dI�|�ۼ�C�=������/�'�p�sT����=�G�=н=�4v�)�
=�G5=%K�l�?6�>�5=���>:9
�9(g�m�\�^!˾�ʒ�B'�<iF�>jr?�@?b�?$c>u�R>���<G+��Q�a�>)`= br��v�5�<4ŭ>��<4� ?}��>:�ҽ�b<7U�<W��<ܸ>���>�F?�E>����e�B���6̿��ʾ�"$����=p�O>��>7EJ=4t�=�ց=��A�����i�J>ac�>m�>���>L��>>{�>�W�>o�>iN>�=
>�)6=�g�����D2<s��u�a=�	F�e��=޸׽k�g�����ӽb��Ot�����i]��0?L�!?I;,��\"=��S�����ŉ��`}�>Y8�>&��>��>�_[=�w��в\���;��D����>�3[?]��>b�H���=]r=��D=��>M�n>*">Z伡$}�㌾\B���>@�	?6*w>A�A���^���l�#��U�>:�W=I��$^�?&}<?k.��wѾ+'�Cb�c	���c>�=�NX|����[:2��?.�l���$���v���k>k?�s?��U�<�4-��!���w���
�L��>��>t�p>ŉ�=���d��,EU�j��̽��->ƻ�>v�� c?3W,?V��>�0�?�;?w�F?�w>gf?Q�=�@>O�2=ZK>���>v?���x�>[:F>�7�=�_ҽb料wMn�F�Ӝ��9>?>9��=�I5>ˌ&>�&=ₗ=�O�<"i�=?>j0�=`�>k1�>�J>�"?b�?�Ծ5�=��3��3=�r����0<S���`\ǽ0��=�x�=�0�>�>F�>��?�C�>��þ������侦 �>#�?�n:?&C�>X��x��=�a��úŽ�6>X��=�ԉ����~(�lj�ʖ(��%�>uu�>p.�=g�_>ֆ�?�B?\;%?�ܽ>.�lq�V�$�&����X鼌�>�@�>e�=,	��6��jt�W_�3,��EH�EK��4�<a��=7�>��S>��=�#>"�;=ii��d�ὮG<d�g��ū>��>�j?C�O>¨I=΄��'"��D?����K�E���d޾W�]��8�=5>MP�=�?�$���{����S9�A��>���?Q[�?��a?�p-�樻�g�Q>�'>wd>�M���?���Cj��8&>T<�=�V���o���k=\ُ>�ڑ>W͝�SBǾ9�Ӿ�|��Af����S�eƄ>{ؾ����]�r������(q�Z���)���fO�q��?߽��
n���X������/m���?�~?�2�>�(Z���A����\�ž�If�;�d�
�h���h[?��������d�%��9�5�V������>��@��o��O{_�x0G������Y�<���>�۾z;z�7�kԷ<�|~>.�>��u�m�x�٨���>>��?�E?~�پ�!Q��y�<�>0	�>��>8f�>�'��Ⱦq�?R�v?�vp?=�<>0����Ҕ��$=�4�?���?�3S?�ka�,�F��YD��@��fk�>�7?.�>d9����#\�=�o�>�^?�j?yo	��+t�MB��2>���>�Lw�a��>�ު>���>��H�V܆�A0P�R�����pN�=�+��ޖ��7�L.<�}�A>4�e=\�u>d��=�ℾ\��>Xr꾛�N���H�ڷ��#���<8F?�+��9>"�g>E>`�(�ጿ���)N��wL?�x�?�nS?7�8?�J��;�-ܥ���=�M�>�>q�=����[�>���><��*�q�����?0�?��?�TZ?�:m�dZٿbԛ��k���p���K>{>�Q>Q�o��[>��	=�_-����[�=,3�>�,�>[t�>may>RCi>*u]>o���^�D���@����4�x��Y+��a���ޒ���+
�IS��t.ľi�t�������A�j�n�!�rd����X�>�P?���>0�7?J,:>��?���.>dh{� �ٚ7��uG�����-�zo�ܸ]��->�����?�<;n.�N�>3�?��F>���>Q�=��>�5�>D��=-�~=�3>��=�?>����.ܺ<`��|��=��=(��>��*����O�u���>��j�Ha�7�?��d����������W�Q.D��.7>:�>{��>L�'�v���^�=�j��>w�'������$�7>*��>�?���D���5��=P���|h��zB�=l*>��=�������R>�?j�Ͼ�<��(��=� ?)�?�/?"".��u>���>��>�*>��;>I��=��_>74?�m?YX?��?S��<ﰇ�$У<�/�<���'���2V��S�D<C���������V�*=�7*>U�*>��#���;=�ҵ=j����w�=m�?��a>�Eü��>}/#��U]� n�����#��}�����-?� .?nF?@��>Ou�<��>��o�ز���Ǿ��>JoҽHV���[��!�=��?���=�?��?�'<=���>��3>��۽�|��d6>ҪQ?m�4>�:���y�f��ȣͿ;u�)*#��Og;��D<�6=���$��<��P��	N��%�����	Ph>N��>��l>P�H>hO>�G>���>^�_>|�=T�c=@���pK��?)�5��< �-��K��e����W�;�Lh�"���3ǽ��ؽM�%͕� �b?_�?j��$A�÷y���򾚋¾]@�>���>���>�]�>b�>� ���T��;��З�ו�>{ML?�Q
?��0� ��=��<��=?�>�u�>�C>R/�NF��EĽ.�;���>E�>{�5>2଼Z^c�"�n�9!�/=�>��=��8����?u�!?z`��ľ/|	��A+�7���ߎ<vS�sڟ����X&ؾ�$��}ʾuR�u�����)>rk?-գ?���5n>�A�Zo���U���Ԉ�m=��鞽{v�>��>�Z>���>s��g̏�WG�� >�ov>��Q<���>>21?`�?�p?,�#?��?P@O=��'?g��<m�~>��T>f��>���>a��>&K�<��N>{='�����
��2Ƭ<F^�b�=0 >6]�=}�;A�m=�:y=>�D=�Fļ�i<<�e�=�*�<��j=��^=� >�:�=K�?�E?O�;9��>��	��Oc�ް�z�?>�B�	��6����T<+��>$�>v�,?�]q>��?����x�<�*��>w�?2?�#�>�Z��}�	>��xW	>!h�<s�
�y�ܾ�派#Q�JY�={V���\>��>Ɇ>�]z>�o?�7?j�,?�>�I;���z�"�8���f���y=�2�>~L�>V��=IM��+��>d�y ^���8�C��J�,��;�$>=��=�]E>=O<�=r�=�d����׽m@=f\˼�p�>�I�>@) ?�B>�H�=����k���J_I?Sc��%E��ϟ��оF�"��>�s:>#���?��
���|�q��z�<��s�>��?@3�?1lc?��@�j����]>)Z>�f>�I.<�?�����ꆽ_4>~|�=w!y�7��]±8�U>��y>��ν%˾�b⾛�B�D:���V��>v�.��K<g�����v='���'G>����nT�hN��d��!F��i��/����}�j�aϙ�e�?pMp?>�i���N���&��l��Ϲ*�XԾ�N����&"U������<��ު�,}��N�����a~Ҿ+��>x@]�4�p�p��z,�\p��
>�*?���a��������5=�Ip>SN�=������x�9W��A�@��N?�kA?��˾Ha�H�����3>��
?�R�>x��=!�¾�k����>�BW?"�7?ɬ�=�K���O���D=���?r�?�P?����$�R�����I%�u6&?E	�>GH�>] ��	w���>-�?p�??	A�>G��6(���Ҿ�j�=��7?x����;F>���>=��>]�Cо��Ƚ�&�=�P���>��l���#��̽<��=뢼� �=#U�>8�X����X6�>�T�.�<���B����{�����;��>������=�~A>R)�=�W&�S-���2�����KCG?�E�?9P?a@?،�t���H���n�>��>��*=v��2�>��>eL꾑<d��8�?W?�]�?^��?sTM?*�d�2Gӿ��������1��=b%�=��>>��޽�ɭ=ĘK=�Ș�%Y=�I�>x��>�o>4;x>K�T><>��.>k�����#��ʤ�/ْ��[B�� ����vg��{	��y�����ȴ���5���Ң��'Г�_�G�5���T>�	��c2�>��F?��?K�?p�>�?�>��r>�A?>��ž�Z�(pB��H7�oM���C���$���b�Vp��h��fԾ��9����>��ǽGc�=�g�>~�z=�{>N(�>�9=��s=��=ִ�<I�=�:/<L�x=�ī�:��<g>�Ż>+��Wyz��B���rG����t���f$�>'����0�T������}��DN>��>}��>>@/��b��a/�+�>8H� /K�o���	��=�q?���>�+0>����=6��s��'��t(>��0>��k<�Z����a�+d�=��?��h�S�u��;�?�_?�=?{C�[ph>Ѿ>8/�>(�>��Ǟ$>"��=$�?oW�>�$�>��>�Ze=�0��DI=z=���=�4�<�f>1Y��i���޽�:�="܏>OO�=j'���/<�->��?>�q����>=��>��i>:}=�/ݾN�c��M��ξy��=N��=4V�>R�>�?+��>}ՙ>��>__���U��/�e���?�D���s�pw���W��Z�>�Cb=&�%?�?�Wo=�KX='�k=�䖽p�>l�?��.?��J>^1�"��9�}	�&Ͽ�T�U3#���ż���<i�<�p�O��<Y���<�J��h�=<�[>��>~!_>�9>��3>�GO>'��>��P>�|�=@�>J�<q]"<�׽l#s=zX������;�?>�w>��Sҽjw������8������}r�2"?��?�K�Ĵ�!�N���W���v�><��>J��>���>�G�=�a	�J�V���=��1X�x�>hg?ٸ�>��D��=�������,��>�$�>E�(>���A	�tU�����<���>%�?��>o��Y�i�p��u��-�>'FL�\�Y�r<�?�0;?9�
�P��]���{K�u4��of>��e���a���h�b5�I�$���s�#�
��^L����>�?��l?�=��V�}�S���ޙ�n]i�g���J>~p4>�\�>���=$S2����'ӄ�*Gڼ��'��rH>���>�I�<�0�>��&?H�?�Pp?�P?�/?������?��=�I�>t��>1��>e��>�� ?�V3>;�> ��<�^q�
a�pH���`<���<�\=1.
>�]@>L1�=�*=�=^e=�h�,��4XT=@��<�I=o[�=���=q�>�M�>��?B����Eo>��i�o����=D��=:e������i[�g�=��>�ܚ>CU�>�b>���>K�.����X�փ�>�3�>��?��>H��x�>S���#��Д>�۷����q����	�
��;5�����>i�>b��>��f>��~?jB?�J"?4
����.�I�v�c+�J/��%=�#��>��>�r�=H�۾�6�\�r�w�`�^�1�Q;�.FG�S6�<���=��>!�A>���=�>[=�$��;�ؽ2�;<����.�>�f�>D?8z\>��=�����``C?Rn��DF�m-��}�ᾥB"�R�>}�&>v���J?L �l4��q&���5�l�>�j�?���?��c?//���ǽ�k>��>8<�=we!;aK������\�/�>���=H�t�⯒���=䭈>�t�><ʙ�j�ʾ�[߾����ʿO7P���7>�c��ѓ����?�������=��l<5��:��>ƴ�����U(�e��; ���Lv���P��1�R�h��?�1b?�0�>�A>��#�b1���|�'���!�����<���:f7�0���C��L<ľ~�㾉�.�/Q&�����g�>�� �`䋿���A�a�{�M���?����-��_�$����5y>$S�>�$��R�k��BZ�=ܓl?o�A?,����s,�;�J�u��>+�>q�>2�>�w�*E���8�>�U�?�:b?��
>L۔��Ǝ�]�g��0�?��?D�T?9�^���D�*�����<���>�V�>�5�>�>�����M>H�0?2�)?���>��3��*�A�s� ��>���>����mM�=j�>�@�>�ý����-�<�����;����QOI�_B=[A�=��t���弬=��?��:�����>_<꾌�N�T�H��������-�<�?��6>\i>L=>��(�y��3Ή�����L?'��?��S?Xk8?�\�������<��=>��>�Ь>�ʯ=�����>���>�j��xr�����?�K�?���?8^Z?��m�I�ѿӚ�����
ĩ�K��=R�#>��Q>���k�=�3��奯��@'��z���>r�J>�G>%6�=%U0>�� ><҆�|�(�!W������T��S��e��eu��7ܾ6)���$��)ԾȕϾ�4#�s�{���l=��7�6�y�ŲK�:�Ҿx�+�^?��;?]k�i�>��==2G�q������!��C�J��1��R`>���U��쫾��$�N�ݾ�>;a��<�X��
�=�O�<�G�>k�?��{>u��>�/�>UL��L�(>���=�&�Y�t>1;�=+�>c����o=W�E>�)|>o�=�'��C쀿�9�'P�:Q�;�C?>]�I��ƫ3���޾-
�����>�?_�S>҉'�`���u�x����>6<F���b�oQͽ`�!��g�>z}�>ug�=گ������4w�]f��o�=�@�>�
>��_��R����gN�=´?Vʾ�o��)�>��`?J�R?7�Y?���>�P>>�`u��p�i>qݻ���==��?�^�>��>g�?C�?��=(��#��<J�`�m{��-��m��2��켼 �����R�\E�=�B�<tk0=��0=�B�����Bɧ��0���?<�d?�:�>�_�<L䥾�q�^w��O���>�&�>k� ?3��>�E?Mb? Ǻ>/���x������!��ò>?j
>��E��R��7t���I>T��>�U?�q?�6�.4��3���87�
�@=V�>�j?bV<?3�?��>Ͱ
�oտ�A�u�C�[�[�o�=k(�=�W���n ��8,�󖆾SvJ���ݽ=_=�h>i�s>3��>�{A>R=��>���>��>;�_��?n����#u��y�j��f�����.7d>9�4>���V$������9,��F>�U�=�f���)?{�:?��f��%{�c�3�@���Ę�Z�?zOD?�?$��>Lj > ��c�������>���>E |?�Do?��E��Π��W=T��=��?Ԙ�>j�?�6�� ����Q���=�#?���>��>ͥ)��We��}j��:پ���>��s��* �?�7Q?H[:�h޾��!����'iG�� �ɠ>��Ǿ�ݾE���Ka�ۭ2�g�,��o���v?=�??&>�ȽG��8��+ɧ�����&���7�>�O%?�c�>v��>�Ç�V�����;�ȾT�������1k>�0>��>��-?�N~?�M'?�04?��=�Z�=�'��q(>Ui�>H��>U@!?Q�%?ғ>��>
�>N�=�'����ӽ��=Y(�>�]>�]z>/��=�QG���������pf�L1��Kg&<U澼X ��8��=��X=9a�<?<?��#?�Iý�P����;�`���l=�(>y�R>�?k� ^���N=�`6>8��>9�1?���>�;�="H��dZ������@G=�y?H9?D>�>I��<�=|=�D����3��Q�6>h}���[K�g@��"Ӻ������>~�u>���=���>�L�?y/#?ɗ���E���R�Zї�X���9μp�0?�G?`��>�q?x��" ����0���`@��V�������F=g���L(m>���>"��>IO>R�B�7B>����R��x�}�~>�?�(?�->i�Q>O{�po;!�N?��S���V˾/��'��<*��>~9>�D?�"�?W��c���L��A�>��?C��?U�g?{��Hƽ8R>��;>���=��<��E��Ƚ�O>ָ1>�4>�B[��aȾ����*�<�4>��>1�����R�ilq>F���<BS�l� �%�ؾl>���z����� $!�� ��.]i��b��T��l��lD��ר���~���>ݽ�ɀ�#�����?Fӕ?>??jq�>JC=��M$�ҋ���۽ܧ��5�|�ܾ���Ks���gҾ�P�6�0�����d���ś>{<X�����}�S�(������=>k�.?jRƾ�������l=��&>3e�<>{ﾏ������M�W?�9?����;����#l>5�?�N�>��#>mՓ��R�fs�>.�3?[�-?�5�(��1��<Ꮌ�v�?|��?�??��N���A��������D?@\?�>L���دȾ����Վ?�2?�t�>�d �G���&�m��>��Z?�J�'Y_>���>y��>[{ �P����b5�S[��Cw����;>�W���o�k���3��v�=!��>�ot>N�U������>�D�(�N�ةH�0��A���3�<߈?���B>�i>39>��(� ��sω�)���L?m��?�S?�k8?|X��F�����‐=a�>�ͬ>׏�=s����>���>�d��rr����?�I�?"��?pWZ?�m���׿%4���Ծ���� =m��=�-�>:�7��Q=ī�jh���X=��>�ܥ=�Q}<��?>��]>m�(>@�>�����%��������8>�������7Ŭ���̇���Ծ�Z������ h����+�a�1r���T��M���T��X�Ψk?h><�}>Z�>��5��=>���۞=�ڽu1�y�����X_U��E��e��f��d��=s���
?x��=�a>���>�B߼�^�>�v>�,{>���=Ԕ>Sa�=��{>g>D��>zk>3��>�>X�>%]�=�[��)���8�6�i��
���#??9y.�)ۖ�=R-��ƾ������>ɝ?�2=>�x%������w��c�>(�!�`�V�XIϽ��V�>%��>5�=��I�:�P� υ�=`���=Ei>�>�^p� ����<��i�=��>ӎʾ�`3�R�=[�L?aiZ?��\?�)�=t��>>�
I�`��$�>�?䢇>Y ?�2?��?��&?x�</��]D��E�.���}��8��o ��>�X>��,>��s=lE=5��=�񄽁�7�/M�������.�t1�#?�:B?�{\=�?{��昂�6	r��1,�>�R8>��%?��U?R��>�L ?���>-�?��N�����񾦶�>�`">׌m����������k>�;���D?sG)?\q�;����>8>D�=��>?Z %?��>�d�>�]>E���0Կ��0���C������o���#=	.y��Bڽ~��<Wy޽�/��/Խc�;9�>�=���=�=zF>UA�>k;�>�oW=篒=u=;=��v��{�F�T<��� }=k{��ζ�T����ؽ\=��{���&�� ��x5;3�'?�H?gMt��Ie�'Ǿ�U�/����:?'4�>��?�U?v����O���i��(���7t�>|�?��%?�?Y�F^�=����S}+>��>���>���>����d��m�Y�M���>�?�$?�-�!j2�uO@��Ɛ�b�>ҫ<�!Y����?[�;?�f(�W9��L������^�)��>q��>����wA	�l!ݾ�-��,���-ݾ���O���2?�İ?��e��>�=<�f�ɿR�����^�{<�^�T�!?�a?b�ҼM˽ +�� .���<M�!�]>?��=
�>��>%q7?��?1p&?�2?��Ⱦ���>Ƞ�E�~���>�?�H%?�E0?�?m?#��>���>�fѽ=}��0��8_��
>U�%>��#>6�=�{ �G
�=63I��r�8�fV�=;Q�G�)��Q�ǝ����=�|X>W�?;?_���:=��ƽ�`���殽2�y���>~|��G���|->�;�>)�>�#?(�>�^,>\�F�F�u�[Q�f�=&0?
�E?A�?%AY>ն�>�����ža�J�1��꛾$�}�����Q��|�=�>��K>�����>��?��?��-?�&���G�Z�@1�y��=�F���?>�Ʋ>��H��8���	�Wa���p��z:�������;Ӄ=�ƞ>�w>�\�>1>��>���=8NL��rH�C:ۻ��q�\�=�g�>�?���>�!�=Ω@��
�,�Q?�!	��E���ɾ����N���0K=|��>�h$�y�?H��n�}��ɥ���G�<y�>�?��?�k?J��s�����z>_�J>�,=����x��#l��|�<��#>M�?>��+�e���"����������9�û�ǾD�t�/NU>�Wҿ�	h��{���b��"so��^��|k�R˾v���Q�e�dc	��� ����]8¾mF�3(Ӿ�J��Q>�?Y�?b��>�	?>�"������K!��O=4ͬ��a����3� f���r�f�`�E�Ͼ����Y`.��S�����>��Y�3A����|���(�俏�O?>D5/?�]ƾ$δ�e��.�g=Sa%>%��<�8ﾾ���S���J�bW?d�9?@P�)����޼>1�?�u�>.�%>�)��X,�\(�>574?��-?sl�����9��񯓼�l�?* �?��6?u�����E��k��}�_��>�?.��>��E�x����½� ?��=?��>l&����z� A���>n�E?��@��a>���>�5�>#.
��A��ʶo��!w���:=��>��������v2����=�>���>�����������>�A���N�^�H�j������O�<u�?����4>i>�>>��(�����ω��*�Q�L?���?��S?�k8?�^�����;���픐=@��>aӬ>ޱ�=}��+�>!��>�e��xr�����?vJ�?+��?�[Z?5�m�18Կ+���,(�a����P>*�\>�E>�i���M=14�="r�i�1=�m�>�xy>��'>0�Y>g�> >'��=衄�[3 �n`��� ���%��T�Ϭ�[�þ
a���ș��A6��"̾j(��y=PQ�.�4����;ԖW�e�<�����ʕ���?�� ?�>�~�>.C<���=q� �_�ľ� n��q����F�w������뒌�>s%�kX#��=�
���"?5S=|�8�f��>
�><��>�I->��=�]�>���=�E0��7f>�>cI�>�Rz�>v^>��>x�{>��=�������g:��RQ�,��;�}C?�*]�7���ʛ3��T߾u�"3�>�n?��R>T�'�T�����x�R��>�2G�:b�'�ʽ�[!�#�>��>��=Ӳϻ�!�:rw�_��o�=���>h�>�m�	����w��=��>��о�.Ž�5�>Q_?�,Z?�Gy?�㩽�>KA�=�K�����>�=0>� ?�?��Q?�1?ٮ'?��"?&�4=\�qD��) �z��"!μu���b<> u>��r=�" ���=�>ޓ-;&��MBV���ͽ3q���+�>�?�o=?�,�>��>]վrd��P�;�=>���<4삾�j*?��?Iք>-}�>���>�=�����¾��Ͼ��>]��>�p>���r�!٪<L�C>� >�N?��-?��3>~�ڽ��=���>J��>\B?0�M?�i.?D�>n��=\3�&\տjZn�7�B��uz=��I�b��;�<���:5=���zq�<P�~�>�j�>�<>/>��>�>d�\=#0�>��>>j�E>�: >�0V����@�'��<>X��=��!=�K����<��>=�d���3�����G��Tw">����%?Ŵ?�� ��w���h�����7[���8�>��>7��>�"�>x��=r����T��b@�o�F�\��>��g?�j�>�28�v��=��.�D�+:�Z�>�C�>�>�[l�$�iח���<���>]�?��>$�3rZ�$o���	���>X�=�1G�N�?��O?�I��n
���4��� �MwN�uШ=klU>�پx����=�Z��:��u�7�پ�0�(?l��?��оQ�����^��9���tɾ<�����<3�B?p��>����0�q�~�=��������oR��^�	?�@
>�!m>���>�P#?^��?�A-?�PH?-�{�(�>;F�=��> ��>���>��?(4?���>��>�:�>bQ\>g���	y��4﫽�AY;H�=l$�=\��=�{	=�z�=\��=g=��|��$ �C����.�'�QF<�UX=��=��"?�L?�M�=��"=�4�H[��7n
>Q�J>&�`����)���y��	>�2?dCd?}-?5F�>P>G~�R��E6=yz�>c�?�C?A�k>T.�>~X@�8׾k�S=��D��,����}��:��cn8��p�=��>�5�> ��>��>�o�?W��>A5��%Ӿ�� M���3�ᭃ�%��>-1?(�>V�ϾxF+�\@=�k�t��ߌ�������?>Ѩ��P伪��:�q>��>��>�
�>����J�=b⣾�/��B��z�}>�'= �,?t`�>�3>�4��5&�4�I?����T��W�����о9�&���>�>>����+?�	���}�����OG<���>�W�?���?��d?�&B�2��΄\>W�V>°>\q<P�<� Q
�V���e0>��=={������z;Mv]>�Qz>%�ǽѠʾY|�q�:�l>��Do�O�N��m��1���+��IȾ����N��7�w=��
���m���#=����`�x���ž��p�ݽ`T
��?J}�?k?��K>�?�m��g��|�m������ֽʅ �L�������("�U� �<�Q�� )���#�Fś>AjY�:��l�|���(�eː��Z?>*3/?�\ƾ�ݴ�n��+�g=�4%>H��<T;�䮋�ư���0��XW?
�9?>�*���@���>��?Cc�>a�%>~����)�>�@4?)�-?�i�*���3��	��Mi�?���?��??�`U��B�����+�?#?�?K�>QI���̾�����?�9?���>2P�z���������>�=Z?J�K�E�d>hu�>%�>�������+�����tt���9>Wu5�]��8p���9����=&M�>��x>�xP�[D��&��>�A꾞�N���H�������R�<�?��5>7i>�A>6�(�����ω��*���L?暱?Z�S?"l8?J^�������ח�=���>Ӭ>­�=�����>]��>�f辎xr����?�J�?���?�[Z?�m�� ܿ:n��BbԾ<S�N��<O�j�Y�>�E����w>��8>3��M��`yT>
(>�";>m��>:�%>��=૿=�&���y$��"��9��A�F�����$��=�ċ�%�%�ܓ쾧=���׾ـ�QP��z�g�fD���쑾20��'���A��.i?���>�����>���;��<nƷ���H�(�{=wJ�q��qL���.���u��R��	/������V�=t���>��x=l�=	j�>��v=[Y�>R��>k��<&}Y>�U+>�>lQ>I�=�с>���>!'j>/,>^�>��=Z���񧀿U�8�[aP��;
�B?�Z�]��-1�?ھ�ߥ����>�U?�KN>�Z(�������v����>�o<���b�l׽��#��]�>�ٿ>���=K�V�vG��t�xj�(8�=I�> �>1�!�y���6�����=�ե>5�ؾ����_�]>;yf?ĺ|?��y?����&>q'>�bZ��}��%G$��)�>&?[�?�?'E?��?	�=��>��j+�%���^�C㡼d�ؽ�f�=2�9=�c�= �>i�;S2Z�>�Ͻ��;�����n������J��w?!�N?
j>�Ւ=N���Z3P�[�c���]>���)w�����>D?��&?g*�>;:\>�v��b���w쾊����>��>��7�A����>��>3���7?�"T?���=�p�����<�?�Z�>s�>�J?�?�8>/�V>���Y�ؿ�&�c2�u�������;�ѽC��<��=�oA������8K���c>ɑ_>��>vU>�2�=���>��>�<>w,�=�˨=YQ�=��꼍h���l��d����� >�'�=x��=b(�~c���7��K�<f�3>h��!�?$?HH[��=����f��U��&2��%��>(P�>�@�>���>[��=+�eV�\>@�&�T�v��>^a?=��>`0�T�=��c����}�>:��>�t>9�(� �b���G�<��>�Q?�>�`/�4W��[q��E���>�o�<oSW�4��?��L?�:7�r���10����<�,�p+
�ၖ>My|�� ���о��[�-�+Ѿ�����O���?m��?2_&��k�s��K`��DX��.v�����ܮ>�P�>���>�@�(G��9�5TC��̾q"�����>��p=�p�>�'?O�X?r�p?�k�>�b;?��h�f�>�hL����#��>Í?��?�!?�:�>fP�>���>�A�>���� ���S��.P�=?`>�En>��>�eM�z|���>3F=v�P��]ƽ��7>!3�<U���x,>��C>���$�?K�]?�ꂽY�#�nZ�=l�^���ݽ)~�>�*?�tҾJ1��_L>:?~ �>b�1?]�<?�>H�-<y9����U0�<��5?tL?�?�l�7�?Z@4�����M��¥����/��ޡ���ξ����d�=��$>�M�>���>�}�>P�y?�bA>ψJ<
/��5��d��96Q�K�>���>�a�>e؈��v��Bn�_������t�B���7��{����>M��>u3D>h�%<s��>H�c>�>��־�(6�'��<;�+>Խ�>��%?�>���Ѻ�<ܚ �gV@?𨧾���_/��t�����=l�N>��<=u��BQ�>+�!���z�#ģ�O�'�`2�>L�?���?�l?�Z��̙��>��=vS;=�.��%�#��ٶ���=�ht>J!>�	�'2��O=��=b�>��W�����'�G���ÿb<Y���<���������������M��)�����$2�����n�x�X���1]�ѷx��`��Z��������?�>�?`��>y�^>?nX��!������o��U̾�Z�5	�������h��ӥ�;$�Ly��G�x�q��K2�M�>��X��5���|�l�(��̒���>>��.?K>ƾ����C�d-i=�:%>��<oZﾽ������K��qZW?k�9?���TF������>��?� �>9�%>�ٓ�W��Y�>=�3?}-?��켃!�����p╼-�?���?D{:?�w�~_N����.�½�{?�W?ʁ�>�`�����[��߲?sY.?�̸>��վ�X{�C��z��>o�\?�C���>>>ǳ>�X�>ę⼽���w���� e���`�MiE>g�!����4���� ��=ɸ�>�an>�tC�Ǘ�e��>]@�g�N�!�H�������aH�<�?���4>Si>�A>��(�����ω�n)���L?���?ۊS?�k8?�]��y��Ӯ����=���>rӬ>��=���g�>F��>�f�^xr���8�?�J�?���?J\Z?��m�uݿ'���ƾ���{%<��W=�a>*���ϧ=>�8�=�'>�f>=2X>��3>�mg>:O>@��=:{�=7҆�yX%��2���E���F��+�V.9�넹�� 	��O�]��_������	�
�����k�u.��l�"�d�������������?﵋>n�ɽ�>-�!��j�>��� �V>���>�K�����B���X�(� ߙ���H��U���D�龭=:6���>��<�	%>"(�>�F.=��>�>P4�=2#j>���=�L>�Jf>��a>5�>]p=�2>/,Y>�"�>#G�=�턿����9���a�Ԗz�k.??z�V�I/��z�2���վN���6Hq>^~?4�I>�U)�6�����w�M��>Ւ3�ګ^�"ӽ�L�X+�>���>#W�=
&���'�k�p��tܽ�ȴ=���>��>��%������3J�=Y��>�1��Ǝ���>Ɗx?�d?���?74��q>�ݳ>6���<|��Ia�>=c-?�>�*?�'\?(?@y&=Zۏ�;C�x�!�0Yž�v-�o����l
>FE�<^�<;�S=�Y(>&�=$�`��TQW��A�Ç�$���"Z!?mc?9Jl<��̼�M��)�#�XZb�aw�����>#�����>�;C?�^O?#�=.�>H�3���S�ڳ���#��{�>�-�>�E���4��ė��p�>!=V>��&?�9?j��Rz��v,E�>��>rf?�"?� ?�i!?T?lu��cr�'�ҿb�$�
u)�����Ճh�	�����[���f�>}�<e�뽍꛽Y<=_�.>{*t>�]W>ؿ%>z>�A'>��>.pK>Ȍ>ј�=���<Up=$$��z=->�J������·�f�����*������a�s��	=g���1�?�?	%?�Mu����i�F���*D��Z�>q��>©�>e�>��=*���S��>��\7��t�>��b?�~�>�5�/�=�#�kO2<��>4��>2A'>�ނ�	b�>���v��;�1�>=o?EW�>B�TVT�Swp��^	�bc�>,�<���h�?p�1?��$��M��nX<����U}S�$��OR>��j�M"���*�r�W���]�?d���Ͼ�3�a��>ܚ�?�����޼�����ה��[��D��O���W�=���>�{�>�땾��*�ǯ��5���
ܾ�$!�S��>���=��>���>�Y4?<o�?)�?��,?Kk�n�>+>�w>���>?�>'?�?2�t>?��>!c�>�_}>����d����F:��ǽB6�=�V^>��b>������;%̗��|!=��漏W	�m�W<�>W=���=d,>
#>֫%=BI?R�N?h!9�*} >*�]=�E���>Nu=��?�9�s��HԽ�0�>.?�;3?DR?�\?G��=�t�=��ԾrU��Z?C�Y?&�R?k��Pй>���,�l�1&>N^���׽ۿ��] ����C�P�e��=89�>>M�>�(�>�ރ?<A>� A�:���C�H���p��cM��P�.��=��j>�N�>WȆ�Jq�1jP��	m��N����|�jĖ� ������=��O���S<F�v>g�6>f�k>��j��,���Q(�ѭ����
>���>ÆY>���>MQ�>�?=�;s�����Y�H?,���r��z���Jƾ^�ͼZ">�4>�R��?�]�U|��P����9�|��>>h�?�3�?��d?�(=����=�S>EM>��>I�<��9�<��/�j�Q=>�K�=�c�Aœ�@去N>M�d>~��.MξY��i�H�`¿�	k����>q����{�
�I�T�־�I�>=���4��[�������.
���ѹξ����0���5Ͼp����?�?���?+��>�
>x�/��Bھ� ��@>ˈ�_�>�y��e̻�J����(���.�R,о�㉾��2�C���>TyQ��đ���}�)�0	����6>�,??�ľj����N��xm=�>�FN<A2�2�����UY�s;W?�O9?=�����s�н�>�
?h�>��->�C����m��>Z 4?��0?*��.s��G������[�?e�?�F<?�e��ZF�	5�X� ����>� ??�>��e�.ܻ����U�?��5?�$�>m?�C퀿���&��>��V?.%A�u:Z>:O�>.ψ>�~�+@��>e��g0��בV��5,>m��!�ɽvH�'A�-�=�ٚ>(z>8�]�4�����>AQ��N���H�������,M�<�x?[g��>>��h>�>,�(����ǉ�����L?+��?�~S?�m8?q?�����TZ���܏=O�>��>WA�=���\�>���>~h�Brr�}���?�F�?���?*IZ?i�m�}���搿�v�'�Ѿ�v>>/:�>L@8��2E��W=>���2\.��Ѿ=��>��>���>�M/>�Y}>���>���!�QW̿~���S�M��"���U������8��!��v��C��4��z��=o�#>��q;"���|=ѽ��=�݁��}�<r?���>�1>�s>��f>`A���]�nѽ�/b���8�>��G�On���ۻ+���p�4D
�6{==��L ?��w=��k>���>rS;���>P�=K����>}�E>�?>��>O�>|��=�-M<F!�=��'>*'>���<�ׁ��z��@���?��k�=�73?V��VJ�:(E�4"���Ǿ�R;>�?8��>�������n�u����>Kޓ��
�J��ʌS�#��>�.�>��=�!2��\���SV�l<Խ?
>>�M>�z�=BY�;����Y�'�3=���>W�ξEE�=���>��e?��G?�E?�?> !)<�����T>'�=�?�??v�j>��?��K?��i?���>j�/>��ڽ��=	�J��V����>���=�~�$"�s�9=4;�q�=L�H>�5>�aA>u�q>�����=X9=;�Y#?�_Z?�O�>��>>W,�����W��u<j�]��>��>@?O=�>�$�>@��>3�>E�=�.߽�g��B��ڨ>cTV>�Q��q�a��=�ܵ=Q��>�KS?N�?R#�<�����|�=��<&��>S?]]W?i��>9�>r��=fM�q฿kck���S���ɾ�����a�=�np�qt�=�U�ݠ��!-�?s����7>+E�>�=�>D�>�*9>�B_>b��>�&>6}>D�>pfh�z�C��-���zռ£U�fF�A��=�G�n�������O��T|_��9�<K�9���>[?/j-?s�Q=�M��Z�4?�&%?g�?�:�>���>�>a���k��
x�x6���-Z>cV?��3?	�����=sƲ�C�=�]>"��>���=���=�K=���r���!�,û>��?�e7>��s�]�S��� �K�����>�m>��^�?>�J?�r�`�Ǿ�\)�<2'���$���L�g=mM��h�����ǧG��Ǿ��O�Ī,��<���>�Ƶ?uث�w�Y��4��䙣�)ڦ���M�4�g>�wN�\=�>�	?'�^�;7�Q�U�mJ���K_�>�&+?�n'>@�Y>�.?�a?�{?9)P?�u.?Jꭾ	R"?ݩ��O�>HC???�$?��>�Ϲz?��=�d���'��[�tH�����=^�>��R>l3>�Q>f�>*/���j޼����X/>�`>JԼY�=ߋ�<0Cl�<&�<�$?ߌO?����p�2_=l'x�Q7=�6=k>�=�^~=aYԽĉ�>��S> ��>�$E?�O�>4H,>�⣻�I��L6�d<��?�<=?WU>d><e7�>������5�1>�W�<�>Wo�����n{��a(���Q�>�>N�Y>m_�>"G�?-�)?���>0�����A��v����/d���C>I��>Qʶ>P1p>�>�[e������ct��z�>J&>����6�<xD�z�,>r�>��}>��>t���.��Ɓ�)1=�ľ���>���>��;?�?�>4��>%Ժ��:N�ɚG?<���>��[����ԾZ-���>�(=>����@#?���.~�A��~�=����>�;�?�.�?�b?m=H�/��LOc>�3\>��>L�U<Ō:����@����.>:�=�y�+ȗ�S�l;��U>�v>'��CϾU��{h�K�����]�iTԾb��B`���d���r����:`�=�I>�6�U���
�f���	>	>�C.��R������p�?v�y?b�>�p�=g�:�Oz�A�+��)g>����~o�=�~Ѿ�n�����w.������!#��/ ���J����<P�> ��f��eu�)<'��}�����=��3?g���N���&�[��=��=�+�ܟ�5[��栿������c?�v9?��ľ����h%�  >��?�E�>��>}O6�����h�>]N?��?�K,�v1���w��@��<��?ZS�?@?w�I�l@�'e� ���U?#
?n\�><����_ξڪ��??K9?�>�>�w��섿�n����>��[?�K�v�a>o�>�h�>�"�������Lݒ�g4��p09>,�@��4�=�e���=�6��=�y�>X{>ŖZ����m��>�+�}�N���H����
����<!�?R��MK>�%i>�8>��(���7Ή��9�>�L?���?�zS?-i8?LU��Z���駽Hǐ=��>�٬>&�=����ܞ>�>�[�Mpr�+���?qI�?L��?�_Z?Y�m�a�ο_[���l�}.ľ9>b7�=�A>�޽����jq�G�<��d=�*���a�>8�>*L>��>l� >��>����j�"�Ѧ�K���:�i��/���W�����������w'�����գ8��2l�R�ٽG�ӽ�F��z���5L>C�?��>B|�>��G>��)>���E��%�r�������9�����̾��u��,�3�g��x��|��b���^�?��a<��=���>��
����=6��>�N8=�+&>�VH>��>�w>>�0>I(R>'>�6N>m;�=��~>��=̈́�U2��-�9�1*T�� �;�AE?A)`��B����3�gZ޾�f��,t�><�?�2T>Y�&��͓�� y�b��>M�A���c�?Eս���0�>[��>�)�=�"����b{�����)�=&/�>�5>(T-� ���q���a�=V@�>�ʾw����%?��b?�?�n?�;F�.=�>��R�7�v�4����=S�>���>\�T?�D?�;?�Ĵ>l	>N��+ֽ�g=�������p�~*���
=6�m�{>�/>V�!=؀W>Y"�=Q� ���=�e'=Bo?�XX?�n>V#�<1ﹾ�_��dA����=�J��W>���>��s>~I�>�7�=�]>�Q�<���[���XC�t�>��z>g1f�n������>FJ�>Ɏ;>~?�I?L���\�>C��>�j>4"?Y�S?��
?S?�=w%�*��x�@�ۼ��s��k�߽ Ȯ=��8����]5ҽ�3X=�8���r>O�?1��>� нp,>���>�ȑ>si�>J�={!e>u>�Bٽ�b�=��j�=�':>٧�=�!#=)���v�=�X�=8.�Y�/�Ε��d=ȴ�=��?9�)?<�k��KO�������� �(!�>�.?�?�d�>�Ň>�Ʋ��+o�mz\����>S1X?s�?�'��Ug=)(7����=� �>T��> p�>/�=�{�)��5�s��>V?��>�kͽ��B��J`�̙޾o'�>�;<�y���?�%?�8�֛=��F��g��H1�lu��t>������:�ȗL��R��@bO��*N�+�;��?��?j{Ӿ7z��i������*��kz��5�`��]�>��>X�T>Y5n��y+��P�my��#��S��;#�1>ex�=JV�>�J?(�+?�jw?) ?�m ?r=��>�?,�<��>��>�>yF�>�6?�@�>���>�i�"5<D��+�DҺ;@0>��o>�*�>d��>π�<%M�m�AF��ݛ�Fo����Q>�=�j�����/a<!���Ȋ?��P?,�@�����>��ƽv⫼U�>N9f>�s@>:����>\v�=��>�U??J�>9�>#����g ��:�;�! ?��6?�l�>��=��7>��8��L��=�R�>����J��a娾I�̾�ؽj��>�}|=��>���>���?��?m�>0���._�}<��L>������H�>��>drC><�>�6G��r��S���|���-�n0%=r��ꮝ����=�V�>���=�{���w?=n�@�ྌ�+���*��:վ5�A�V6?�e?��1>�̺>���6�'��`I?o����e����oʾ��$�l�>:7>�����?�t�-}��!��1~;��.�>	�?dK�?��d?�F�� �ʛ\>E+R>0�>�|<�n?�v��0��d1>�~�=6�x��̏�~/<�_>�
}>�:��%�˾>�/�@�Fد���o�ϯ�=�!]��	����=*5��u>M�:`u�̀'�tž��KYC>;;޽`g:��������}�,�t�?��=?�8?�E<�e���ͽ�a˾��3=����$������L]��(��}Wھ����捾��R��l>���Bܢ>CY�q���~����-�	Q�'*�=�?]����4��=��b��=]N/>�c�
��u��*���5�̦N?�`6?^{Ӿ���.��4�">��
?�J�>�->1s/�t|��2�>��A?� @?�=��������	�L<��?���?M@?%�4��L>�����C*��| ?�?���>�s��a��=�罗_?5�<?Zק>Gs
����O ���>��]?�<K��fT>^S�>z_�>b�������W:������,�w6>t�&��(���i�V�6�s��="P�>W�x>%/^�����E��>@�7�N�[�H�������i@�<�?;��6>,i>aC>��(�����ω��*���L?���?M�S?�k8?�]���������̙�=y��>�Ѭ>c��=���d�>���>�e辻wr����?�J�?h��?L[Z?��m�A�ӿ̱����Ǿ�R���_�=(�>z�;>����u��=���<�E5�Bݯ<��>]��>�_>]�f>ZgO>�w>�ʂ>�u���$$�)���|0�� N�^�=��:ox�Y���Z:�D!�}Jž刾��޻!r^�I>̽zg������9M�:r���,=��?�>��>p�>�:>}Б��TҾ1X�����4�#�~���������]Y�W�I�rƊ�����ԣ=���c'?O�=!�=$�?��[��]r>l�>:] >WOl>@�#>#ѱ���>N�L<��=�v~>>=�Og=�v>9��=����t8���d:���Q����;��C?�_�c���up4�0�ݾ�����>�r?�wS>%'�⓿A�w�b��>:�?�!�_�AĽ� �4�>�
�>^Q�=f�ûv���kv�������=U)�>��	>��H�M�����Ob�=�"�>�s׾F:���W
?f h?l�E?k�[?�z��&�J>��w> O�>`�w���G��>��>��?��B?�m%?���>���\L�4x�<��<����,��4��=+�(�k!m��"��{n2>V�>A���p���J�=�6�=�O>�*�=�?7vb?�/�>��>{�o���>��L>�D�/?���>�/�>���>�N>`�>פ7>�>��̾�W6��/�>�Wu>�Vs��T��R?=Ú>X��>^'7?��x?&2�<3����z>�����>�?�:�?|M?�?�1�>����ſ$�4�xPE��9y�1�[�d�?=RL�f�3�e\���V�����p>tL?ۏ>$ʗ��BŽ�~�>���>e�>(�>%t*>�,���4�6�y����=P>Jc�E's���k��m�=5>��<pК�Ӭ����z�}}\��,?X,+?�����Q�������먴���>`^�>�:�>K��>h'>qFݾ�uL�u:��e��+��>²X?~� ?��3�vP�=�#<��r��#�>~R�>��b>C�нf�齟C>�O�G=�>kR?�>�K��a�T���Z�lo�M�>�g�=9-��p�?d�?����Ǡ�-�X�����3�_��=�0��<�Z���[I���b���)�x{G��*Ӿ�X��`y ?O��?g��c�Y�~�'�.s��J䂿��:��YL>!�>��?.?S>ъ:��N���[S���ܾMW��C��=%D�>��C>�Q>l�[>�?�V?q?	�.?>:t�{?���>y�?�$�>B+;=Zt�>��?�y�>�t�>(� >��=ME�vM���ɽ�.¼�+>�f<>a�7>�2�vY�(ͻ=��=.C��Cm�T��:E�=E떻��R��9�=��>dS?��.?][��9@����Hp��HZ>��=	��>��[>��=���=��<���>�?O�?ゑ>�����������7���?
�0?�m?_��>�C�>�|�l��cG_>3<�>{H��������T!�qo��[;F&��:�=0C�>\G�?� "?Ì�=�!�.�J�KD�����9Eν�>�H>�2<=]+�>^$r�2{��]ˋ�Ùx���W��E�Y�&��H��I�=���>pO�=��.��>Ôc>n<���,R���B��6M��w�>݆�>��=?�S=��>���5\9���G?$������w��'/��ďz��3(>�/>�wҽM�?��ý�:z����/�Z�>Y�?�B�?�_Y?+�O�����s9>�n5>��>wI=��*d�珞�ܭ1>J��=����uߑ�V�a<!F�>�_>���헶���޾�{6�����\ri�
�>+ா���=.	��~��>���r�A�ǲj�/�=/E�h�0�}�d�tƬ��R����@��|�?�zD?��?[+>t,��,pľ�[,�V� >hR����/�OH ��0@��S���0=�tɾ6"��Hk"��1.�%=�@��>mdP�㏿V$~��)*���ۼG�/>2T+?�T¾
���*��N�=/�$>1_<������>���c��W?#i8?�w�m1������~>��?M��>�!>�퐾݌Ƚ�̗>#1?�/?W�F��`���,x��b»?�i�?S�??e�N�~A�A��i�W�?WU?�	�>jr���_˾�
 ?t9?���>�5�],��F��P�>�b[?O(N��`a>D��>�b�>	��&���mX*�jj��xtj���9>$�
��O��f��r?��/�=fˠ>0�x>}�\������>"�龛�N�|�H�s������<Q�?�K�G�>�Di>�>d�(�������� ��P�L?͒�?"�S?f8?�2����������N�=��>QǬ>\L�=�����>���>˖��ur��<���?A�?���?7uZ?�am�U�ȿ+��?���K��<�t���=�N��*%o<���=�-<>UC>Р>N�s>��8>��+>���> �a>
�z=[���)�$��L��n>���qb�Z-��3�-�Ҿy�:��C�hl־�}���������藼RN�"�p�~D�dU��t��Ȩ=S?���>e^�>#h�>곷=�K����U��k�������������5ɾB�|�T�t�ь��#\��zB��~��te?h�=�B�<_��>�9��F@>%��>+"=�>�j>ٮ5>��%>�>�QC>#>��M>��/<܊z>o%�=_-���	��P\:��Q��+�;�wC?�]��;��Q�3�l+߾<N��e�>D�?�\T>�`'�������x����>*F��\b��Y˽=��_V�>а�>�#�=��û����w��H�b�=��>�B>K�j��"���X����=2��>Qtp�mI����>̪|?8e?hu?�.�>}�;?�)ؼ/a��1���R.����>�a�>+	?�]W?g~[?N8?��<������[Wh=sнJ�!���z=��c=��=��.�����Eכ��V><��\�'b�?��=�=�=��'��hF�`?�^R?s��>V��>��$=�3�)�*�')�=N�=���>+H�>�;�>S��>���>e��=�o��P����˾F��>��3>�~N�}@��dW���/�>B+3>�[?�J?E9���ޙ<#�[�E��I��>�a?ϩ+?�q�>���>�濫`���T�F�6�)~��A�3�$>ꈾ�*���C>;��>���=NŐ>� ?��>[��>�\=>�����I_�>���=�_">��8>��=U�>v2=�>>i=U�����#�$����<Za�=�v��7`��h�q��Js�����s.?��<?�y-�݊߾nF�v����D?"߻>���>.��>��5>��&�%ʏ���о\I�]
?Hw?KR*?�S��K�8��S��=��1?���>;{>/������蹖���"=��?�<�>��}>�7f��EW�IeV��.ԾD��>��8>��ȽS��?f�r?��:�mb<�uL���������y���ڼ)�������uc����N7r���漍�!4?���?�¾�.����j��F��� N��־AȎ��f?�b?���>�uo��,_��0W�B�k�e���{�ݽ6{�=#��=_�>��?'^1?>�?�??��$?�x��:�@?�M�; gu>�4>.h�>� ?��>�D�=��>�k>�3>�\ܽ�F���K;�ָ�G, >�6>��>��=q⻞%r����;|�����e�Y?}=�|^=5��=�=]h=��S=��?�@%?z������x�;N��@�T=�X>C>��w6N���=�&>f�>B1?u_�>?��=C��:2¾�� ��b�=j�?�a:?���>��z;�j�=�_���h��I=��5>�ʖ�%�y��̾_�R��%�>�h�>�D�=�r�>�i�?�*&?�;*? �	�\�r������7��c�����>�-�>~P>5j?�Q�Ϯw�X`���G���C���ɾ�l8���{<u��<?\>�K">3�>���>��v=>�&>�88�������"�>0�>p�i?AB���>��y<T��!PO?ݾ\�����ľ��x���t�='��>����?v;�������򥿶�F���>O��?�-�?��d?�s�}dֽ�Sw>%�>	��<cv=�����O<Lq�=��>�{�=t�{�֥���Glj=�]>K�ͽ_���Z��h�N�O����[a�LH��m���W����Nð��@нԎ[�����)�J��������Խg�˽�V����ؾ���|B����?�}V?*a?�ak>s�1�W�a�9�+�%q9>8�5��oپl���Y����M�N�����׾9Ƽ��:B�ic��^�����>��Y��@���|���(�����+�?>K5/?`ƾ�̴����Ƹg=HZ%>�q�<�6ﾬ���ܮ��j�cW?��9?$R��&��sί�>��?Es�>ſ%>�(���9�%�>�74?5�-?�/���:������l�?� �?\i??O�׺9��]	�� T���	?�$?���>�x���ܯ��ϩ�j�?�E?�+k>��̾�}�����w
?@t?D�k� s>��>k��>h���΃��oϢ<���G��<�,�=����d7�φ&�Gw����^<o�>!ȇ>V��������>L�F�N���H��������n�<�{?t��n>Qi>�a>_�(�����ǉ�3���L?Ώ�?ѐS?+j8?X��T��Q������=��>�Ŭ>gӯ=����˞>��>^�tsr�*���?�C�?b��?+PZ?e�m�{˿�]��qt��V�����=�{�=��d>�8��K�<!���G�����v��>�t�>�u>�Zj>n�p>��;>�{W>+ň�c�&�o���'���/i����F�cV��]Y�>n��+�(��c������!���@��I��j�U��i轒���D�%s罂c�>�0�>-�>Ϳ^>ڱ>�XW���Ͼ�­����8���*�#��Sn���@�pY����u�Y�(�=�?�=0?!v�>�=�� ?7Z���>Au�>��Ӽ�A�=��.�!}�=\� ?�(�>/�;>3�>3�j>Q��<|�j>"_=Qy��e/��+\7�Y�I� �;�A?g�[�|՜��.��Aܾ�3���z>
?��U>N'�P\��/�r��8�>��e�%U�[1���!�4�>�w�>_��=����d"�eox�-����=�n�>ʿ>a:����������=\��>�,�������D�U�r?9�Q?��$?~{=ҷ�>���=�?��>� �>��X{>�J3?�?^�>ݶ?b0	=#_��"�pHE�
�j=�Ӫ�_b� ��Q��d����>�oK>RUo���l��hr=�i7>��꽶MI��>5�	?4�T?�(�>\s>������5�O T�,@�;�%q>��=j��>��Q<���>��>��>��G=Cǽ�Z���]����>5�E>QwS��2c�!Z6��{>\M�=�-S?U3b?ۖ?>�Ž����	��>�?�o?Ρ%?���>qĽ�a�2̿��J�aT���0�2�s�ds1>ͫ����ƾW�2��_���PR��tY��9�>
=�>���>���>��t>iqI>�+�>�^>��<�~�=�,r>��߼�Lʽ��!=$����m3>��>�A�=������n�Պ4�_y�=ş�<�n�9I���?�O?�9�����ӌJ�3���S2�23y>�) ?�<?��i>�b>�Ξ�YI���)���b��!?کx?b��>zc����<K���O=�V�>��>HA>������4�����I�;�?�>��?^�>�r��+�h���[�D�ݾ�ʗ>�#�=�=�-�?%�g?[�&�����4JF�s�;�~Z ����-h*�T�N�4e� K��,_�������/���%�+���?Rc�?�B����Z��(��+���k�����[=Mn�>.��>/�>&���8ž���4+l�ؕ�
�>���>6��=�^8>l��>59?R�i?�0<?�hI?�eu�K��>�R>vd==�i>�4K?f|?�_�>�tx���>�@�>��>R����־K�νQ���f:>��`>�k(>ђ�=�F`������=���i<1��=�D�<���=2��:ļ5�[�<�F?&,?_� ��L�giܽF;A��*�=��j>L6>'?>����ʽWɓ>:ȿ>3uM?��>�Ř>V������۾ä��6�?	�>?s��>#7=��²>bS��͐��>;I� ��#>�����`���傾%4>��>H)L>�9�>+��?�3?��>끸�Lol��/������=��>��>���>)�f�)5���l)���y��Yd�nn/���G��c�����+��(>*��=�D�>��>��=}G�y%���E���ƾW?��>>j"?ٰL��͒>�o�	v	��	L?ݜK�7h�8�ɾ. ھ5j��>!�=�)�>�Lȼ#�?��憿�A��� (��?�6�?��?w�b?�0x��߽G�!>�K>*�>�?�<�/�4/�=񚖽&�='�>� ���u1�U��=�V->�m>�����o�������Р=譲�b�w�4"�ug(�=�z�bۚ��7���J>����ʾe�I����l�Ҿg��h����;��i�������[�NW�?`[?b�?Zn^>�������k��.��N�#�)�M콾���� o_�.Ս��O���������*d9����\�>��Y��=��`�|���(�|7��|y?>+/?�cƾoִ�C{�2�g=��$>˘�<rGﾩ�������1�!eW?�9? M�O����S�>\�?M�>n�%>���//���>*#4?�-?��꼆����,��ד��S\�?���?��=?"�,�u�6�ͮ�����7�>�)?֣�>2kK�;ԯ��A5�]?y�D?V�>`��o������3?~�U?��n�8�=>ա�>�O�>�v������䉽���B�4�7b)>� ���B���L��p��2�="ؐ>ɕI>�Q)�c���k��>�/꾻�N� �H�������pv�<p�?���QK>yi>�M>��(�,��6ˉ����L?T��?�S?�i8?SP�����|��=��>IϬ>���=���-ܞ>i�>La�u}r���[�?�J�?���?`Z?�m�9Gӿ��������F��=8%�=�>>��޽ ʭ=s�K=%Ƙ��Z=�d�>���>o>W;x>��T>қ<>��.>o�����#��ʤ�2ْ��[B�� ���wg��{	��y�����ȴ���J���{���,Г�w�G�i��U>���վ��"�tH?mb>�k�>L��>��A<l���I�����l���\�ƾ�V���I���V��Ž��a�5��ܓ��0�����=@4�\d?��F�^��=ۧ?���2>�#�> ��n;x>�ƅ>v$d>.�>��->a_>�D�B&�>}��=��{>7u�=�%�����X~:���Q��]�;��C?��]��)��i�3�lS߾6���$ӄ>}?_�S>��'�������x����>�F���b��̽�Z�,S�>1��>4+�=_���{s�ߤw���h�= ��>�B>g�������%�=�7�>$]̾S񶽨��>��k?���?��Y?R�C��?2W����>܁1����;饣>K��>X=4?�,*?�y)?#�+? �<�c����r�T`�=�����޼��]��؍�  �h2�O3�i����;ͽ�C��w�=�>�	<�p\=&@�=�n?��<?崉>�k>�����:�
_*�z�a=8�<�P;>��>Ȉ>%��>E&??�>�3�=2H�=_`Ծ����k[�>�I�>�Zo��N�����
P��hT�>�v_?��Z?jj�=�=(=v> n���K�>r�>?�g?я?�?�d޻P���ѿ�����r��<g3��}�=�����[X=�ov��8Z���Y�7�j{g>i�8>�D3>+�>jψ>h��>��>��=>���=8!	>�=��˽%4C���}=������<;΄���X�IϾ:��4�`���������:I��J�s�*�?Y�?�j��#	�d�Y�e���x��5�>��>�4�>��?��=���@�C� ����.��<�>�n?l�?�l��[8=M��<�_�=�Ğ>u�>]>+��qF���5<���>��?��>{@p��hc���l�u)
�K��>�V�=~ @�S)�?=�J?��T����`�8��e���&��G>>�詾/X��mA�+f��'L��"���A���侤�9��x!?I�?�����3= f�����i��q�Ҿ��I���>�$?�֑=�]����پj7��!þ�(;������>�\=Iq�>�?�i:?p?�/'?~	A?���$d9?�ڞ�Yx�>K�>6�?zQ!?�>��>5��>:�4>�s>�Em��,�:S���b*�R�=�	�=݁�>�5/>w�=ԔӼ%�=��g=DU�.�h���7���=j��<��<�	?��2?~�6�I����?�<�պE~�>�P�=Ǹ>���� <Ւ?�p�=;b?Qt2?�~�>�t>�l:��׽��(��d���;?ޭS?��>3v�=��n=��-��=����<VC��*�H�-ʝ<jl�w^�06��?�=�!@>/i%>7;�>�oX?e��>γ?N%���c��V��s��_¾Aז>P��=TR�>���>�R+��SZ�
�T�ITr�^�L�bK0�F����t���?>�{G>��>p�;>�qU>&*�>�������G�[�C���>�?�"�>�h=}��>��]�q��ƲM?k�=f�H���4�n����J��B1>��?V�=�0�>_�>�1g�2��
���J?���?�b�?dHw?�~�7+��ગ=8F�<{)>�k�==/8=��d>m`N��Ƀ>R�ܽ������]���<H�>�c��_��,=]����>Q�����w�X.	>@���*v6�>�u�ޥ��m�D�kz�� �z�&���r�{'s�9�<~�9�k���p��#^�� ⾻J�?��T?Qو>~��i9;�<���� �(�E���}>����@�����@/	�䵾=��ɹ;���Q�ArI��͛>QiY�>��!�|��(��d��'B?>J"/?�lƾ4��� ����g=Z%>Ἧ<M�¬��	����>��XW?�9?z6�I*���D�5�>��?5b�>��%>���Y��� �>�A4?��-?� �
���/��԰���h�?���?��??�8M���A�+��Y���?�c?�"�>������˾��RX?"p9?C��>j��d��n����>�o[?c�P���`>�w�>�>���OO��.a �D����و��:8>)���#�mkf��;���=��>,�x>�]��R��Z��>8꾔�N���H�E������g�<��?L���A>Ii>i4>ַ(�'���̉�4&���L?җ�?օS?m8?�U����秽�m�=���>��>���=�����>��>�f��qr���B�?�J�?��?bZ?�m�=Dӿ������~�����=�a�=i�>>�$߽
�=�LK=Ȝ��Y�=���>p��>��n>O<x>��T>c�<>/>v���#�#�Pɤ�{ג�`YB���n���ug�~	��y�����Ǵ�g�9f��������G����p>����D�u=��?;m�>���>d@n>х�=^w��D�ﺾV�۹�������m��Y2���8T��qܾ����� ���s����>�9����<od�>_�\��?>y��>`g�=�$�=O�9>[P>���>k��=&�3>���>Q��=��*><��>�>�_s�֭t�[19�?t�������F?�ڝ�?��_��=<��h7����p<c?h��=�_4������p��>�>e�`$�܈��(�<a��>p��>�+?>v�L=�^�9��j�D�'�=��?>�.>��K�E������X>�Y>
������d�>��q?�}l?0)E?�]��|&?�f4>���>�.��t&��
�>K��<�>}=.?��0?͛-?�=ihľ�"V���K�d%:��:��a[�Z�ؽ�e�G�>����B�";@p%>���<x˽���۽�,==D�]��!?�K.? ?:>�A>Y����x���?��F>�#G�(�5<R+�>5�>��>�|.>�&�=��=T8$��L��z�f �>��>�,w�Ė�Ƴ��0kr=�d?o)8?�du?�仉R���=GHB>	�A>�l<?��_?b ?���>�,�<~7���տ3��*�7�K�$,9�̓=h�M�#�,��&3�}N��8½c�<U�>���=WF>�?A>w�N>/�G>��>��>��5>	��=��h=D��=�	��1�=g<��S
$=��=<�^=(Qe��t��W�����V�����u��V<��*?dN?��~;��_m�`���A��j�>���>�M�>�?D;�߾:�9�T�;��q�o�>"�_?+��>������=�V=�z=l�>X�>�6>�����,�7#��	�<�*�>.�?�ߤ><���_�!n��x�Ig�>\�o=Mp��Iޒ?�?�*�4���{Q��Y�o� �X?�>���+�z��ؽk�(���&�32�e���z�^��"2?�8�?	��L&>Ij ��״�����Cb���&l��W���_?WGL>��<�	����_���]��Β��iн���=}�P�$'�>|�>��3?,Vu?V??�,9?��ɾ�\:?u1¾���>�>t��>�K-?�@�>AF�>�l�>�Pn>�e�>��]��ġ��x;m��\0�>z�>��	>���<�`)>��W=�i	�D��=Ե����W��i=�#,=y�ϼ2��=(o)>J�)?��6?�R�5]��x���ZK���>[��>D�>
>o�>������>��>�r4?�>?2�>ы�<t���)C�z�b���?C�:?��?�c>�=H>n��HS����E#0>in�z�ɽۛ/�\�����X�*>;!�=BU�>��>Ǜp?�=?�d�>n�C���>��3��#4���@�j�9=g��>n��>X�==Q0����|�4~�:8��Ci�����D��_�<>^|�><�=�\>/8�>��~>uˍ�M�"��R������*Q=�V�>���>�����Ta>�㿾�_Ҿ˼M?�*�����ڻ��qݾ(�Q�)>��o>�AŽ��?��ʽ��|�����KF-����>B��?���?Ʊf?�Z���/�k&J>(O>ɭ/>�<o�����`��m:>�B�=8I[�������;.�g>SU>�x���߷��ؾ�hm�a���5��|�>��辪XȽ�_ݽvX���>n�
���t�ͽ��T��m?>�F��}����H��nހ�P����>T��ݾ8�?��5?�l�>,\d=~G#���Ǿh���"J=�f��I�N={r��M?���I�̈́��G��㸾��3��6���3���>�Y�4��?�|���(�vd��X�>>�'/?�pƾ�ȴ���>�i=r�%>K�<��Y���k���ƫ�82W?�9?Y:쾢���i���>P�?�M�>��%>���E콚��>�4?�-?t����5��`Y���c�?H��?�@?aL��\A�bD�|��B�?��	?���>���M�˾41�l?��9?ٸ>-����|�����>�5Z?~�O�(`>e��>��>�mA��%�$�C:���r�:>�b��
��5h��<���=I�>`�x>B�Z��X�����>E�d�N�èH�d��8���B�<.�?���2>�i>�=>�(�	���Ή��)��L?���?މS?uk8?Y�������Ё�=(�>Xˬ>���=f����>I��>�`�Vtr���?�?�I�?W��?�[Z?��m�X�ϿҖ����ȾZ涾Uk>��+>;��>D���2�>$^=I����b�;~zg=s�>��V>��g>��8>$� >��E>K����?+��s��K����R�!������{(�'v �����������]�����<�>��_�oCr��D7�{�B��˳�+�N�5|5?-��>�4�>��>��=�X���g����F������\��������������|��^�j�(:J�#�6<Ƶ�	?���R��<�I�>uM���4=�>�>��=a)>+�j>���=��%>W�>�j�>_�>;1W>�}����>�M�>�m�d̎�	7D��eܾ�d��G8??MǾ.y]��%����/����W�L���?pY>��G�l���Y��*��>�,����`���Լ�I�'D�>;>�>�*\>�[�=�	Ľ���Q߭��<�1X>Ԫ�=���0�/�6�3�`��>��>���T�ɽ��>d�i?�b?s�S?b�}��
?������V>Np.�R�0>�A?k��>�*;?c�P?Md?�8?U�5=���a�z�넂�㞼��<�` ��Z��Q�;�5=��S��g/=�b�=��=2�=)z�=�fU��fٻs��=��&?} ;?2>}�	=����x�"YW�e�<Mǒ��6>�" ?�2?u2>�0�>��>���<�����'�|)9�#��>��>s�y����\;>��=xm�>�RH?�LO?�@��x�F��v>:�W>0K�>RO?��Q?lZ�>�ʹ>��A�R����˿1���T�Ңu=q��<�b_=)�$�D�=�	>B��@��sK�>Tc>ZӼ��L=�s>6U�>Tw�>�v�>�<�==xh>���="@=~_0>�g���=�ї�sH�>G�W=�R�=Ѱ�=1������Ί���$s�9{��bh����?h�?���mF�SL;���������>��>���>ۛ?܈h=J~
�q�F�#�8���2��>�>Ìd?�f ?;#B��J�=*�ͼ�8<D8�>/˭>u�>�_�����{�����s��h�>7�?�"�>D[!�H�^�c�o�\��t��>r=��S�ؼ�?RK?�,����M�?���\��~�AҴ>S�z����=,u�:j�D�{:��bžN�&����/��:?[�?A'�ۆ9>|*�ּ���q�N������>ډ-?���>6���k�c�e�=�2Qо㟇����"�I<l�g=&P�>���>l*Z?�\?��>~(%?'nξ,�9?��H�?Ϧ=���>G?��?�#�>3�>�4Q>�<>���ʣ���=�	�<\x�>Ubj>!7J>�	�=c�ü�D��	:]�"=$k��(��t8��['<k����>�<�E>�"?O�L?*оY�����t��j�n>�	$>�F�>0V_�S��<a'�^�=0�?)�)?b�>-�w>�r��霾��%)���?rba?�n�>�4�<2�=�L�Sy�;��ݽ��E>�՘��)�J�%������J�#��>p��>���>�J�>?um?�?�>!?7ˍ���4���w��D�������Z���>�͑<.-������]�����ڡY�edd�}Q<��y���n<0�=B��<:�=̮;��>���=�y���潎��=⒄�#�7;K�]>��>��=�y>���r��PJ?g���1��]�����Ѿ@�&��p>1�D>�� ���?��t}�?����@;����>���?5&�?��c?�D�����%_>�jQ>G&>ϯ<�M1���ؼ�q��^�:>j��=��v�5G���<�Z>��t>�˽�{ž�$�)�2��s��T���#�>��վ�� ��,�=��ƾ=H<>���g�`>6����v����K>�oŽy�k�����I���u2�^��?+�Y?F�>>M��H>�>�ؾ��	����=�ĉ��>�Sŧ��v�����s������o��;�*�i,�nh$�A�>��W�Q����|�W�(�~�����<>�U/?�ǾVŴ�q��h=�$>Í�<!�G����������ҵV?!F9?&$�]���G�ڽc�>��?��>N�&>�<���-�>}o2?�-?��἞��Tn������;�?t�?[@?D�B�n/B�Ş�Y��z�?�.?��>FX����̾"ｆ+?߾6?C�>������6��`x�>%fY?��Q�ͩ]>��>ǫ�>J�å��|�� ��<.��0>����B�g�n�:���=Eg�>�z>��Z�ȑ����>0	����D��0=�H#��D���.�Q�?}����g��F�=�i�=�5�0S��������q]'?��?�M?g�??@���e��`xY�� �V�E>�zo>ܯ�=��*��;�>�T$?�����H����Յ!? *�?q�?*R??ዿf�̿ޘ�)��㝿��=�+>W�l>��M��L�=Pd̼��m��<?>���>� L>�i>w_>m�f>�D>b����*������ԓ�6rX�tc����﬐�NA
��Q����� I���G��{$�<3/�����
T�/H�\o���	�������D?�%�>;�>��>6�<V9��B0��0�<�̾;������7��D���i����o�䈾ђ��~��=�?׾8�?���Wp���%?m#�аg>�}�>�ߩ=���=,cK�_0��ֆ�>Oٳ>�W�>�2><�>3����> LJ>G܆�o��	�3��q����2�6�W?��]�|.�����3�����ξ��z>5-?��F>������ӽ��w�>�~<�.��͕�:W��D��>���>2�=w�->ڼ3<ֺY��� ���=�x�>
�6>t��=1 �h�޻td >n=�>���n�>ֆ ?�'l?�B�?�h?�_.��8+?I��=��|>u��==@�=���>A�U>UL2?�QB?��??b35?��=#m��F+w���<ـ<u�>�W!;�C:<8����k����2�>\W>`=���<�3e��R
�\�=B ?�I?���=�U~=s�m�.W_��G��#>����h2T�%��>�G?�v>൦>���>߉=r�=��ž
|<����>x�>ˉ_�T���˘����>o�I>Z�>?�*N?0 =�K@��A�=����O�>q�(?��[?'��>-E�>u�B�#=
�k'ҿ�)�e�,ݩ��9����'=գ����<��d<~n���̼=��>Ф�>	�>v"�>ި\>Ň_=�!�=�z�>f�p>bI>��>���$i�����v�?-:��#>!{���=vcM>v齸S�����h�� ���󢶽��?u�?ǥӼ-!P�n�b�����hC���2�>e��>���>b�>f6=|
�4�]���E��
c�;��>�U?*?�cH���Z=J4�(�=��>L�>��a><�.�nv"�����f0�3�>���>v��>�G��g^���g��
��$�>l�=�P&��y�?�Ho?*�;�K[�E�>���4�M!"�t�>��
�Z�������C��l!�9���94�s&�W����?�?�K���F>+�꽾���ߟ���ʾ&��N����	?$��>:f���tھ��9�۾���8哾��)>�W�=B�Z>T3?�H?�$�?��;?�;?ъ=��I'?�r�)�l>>=��>h?��>��>�؜>��(>�0>�Y���Bþą�����"p>ud>p��>(E=Ī��6�=o�<�˛<ּ�=�ӛ=d�==���=)��=|��=�|!?��B?��澌� �l���A�y8>Ql�>��?3羾�Ⱦ>|����Q�)�$?��m?�=?`�?�<>^O����Dԫ��=?PBI?~��>ǯ�<��!>�G2�2d��=�<��>�q��/�������y��_Ǽ�.�>�&�>ď|>��>�
~?- ?��t>�hd�r�@����&S���`��c?>�k=���>f4b��C��{��v�R��3P���5��_Y��Z[��B�=?>�>�jW>wh�><�=7<�|1���}���о˛�=���=ص�>2���;�쿽[^\��]K?)"��	_�"����IϾf�<��u!>��d>���GF�>�?ɽ�mw��ؤ�mF/�*0�>�	�?�h�?�f?��:��$��L>o�[>�R&>�q�<�P!�~��������H>Q¨=�Fe��j��te<�UV>��g>� ��U�����۾�缊��&�b��=�=�,��V��������N���6��q���6�=��־������>M���/�0,'��[��Ƴ�3���|�?��i?q�>���=����E�����,n>{���b/�ž:�*��l������{��7F��l,��T��ԃ�>���ښ���e�g��0�P�r>�b1?�^ݾVU� ~9�['�����;�� ��
�Z���U蟿&Y���b?p]'?��󾺞�XŽ�&o>��	?�9�>�s�>.A��|v�y�P>�,??�=�/m��Ԍ��Ep==�?�H�?�!??}H��~@������k,?
�	?���>Ů���MԾl�
�}�?A�4?	$�>���\��������>�>\?W�H��/_>�?�>�x�>��罍������Q���pk��8>o�*��s�Tcb���1��V�=o֟>�8�>�R�>Ȱ�M��>�@꾆�N��H�'������N�<�?c��3>�i>k@>>�(����yω�1+�j�L?���?�S?l8?�]�������Z��=���>�Ѭ>a��=����>I��>�d�xr����?�J�?t��?�[Z?��m���ѿ����>�ݾP��of>��=�v�>Wc�O�>�Z7=ng��*�5<8�>�W�>s�7>^&�>���>o�/>���>����Ry#�wI��������L�C��R���j�x�^u���� :��~k���$^�l(׽m���E��B�; ��u��'��<d�?L�?���=���>���=�m���s���Ⱦ֪��s��ؽ�o��J"���߷�����þ��6`G<��k?i ��zn>ַ?�+"���T>7K�>@5l�Eb�>ѓ�>b��=R�>�I>�۬>MO�=E�>�k>c�>Uk�=�=���P~��5�v1Y��_?<�C?�:[��+��g�4�Bm��3��`1l>��
?�B2>B$��G����v����>$�)�Y]�+
꽾#���2�>19�>X��=��P;��?��]m�|��W��=~^�>��*> s�x���'�k0�=P�>��mb<RI>ȫW?:��?A�c?־,>�� ?��I>%��>,�Z>HO>��>%N�>Ge?ʦ<?R?V�*?��=�r��Ϟ='H=�N����DI)�]O�8���7�]=��u=;�=�>��>w2���r�;�>r���8�eT=I�?5M?�b�=�b�=�u">4k2�q*1����=I0H>�ۓ� V�>���>��Y>���>�)?�}^=jʼ�z���W6�>D�w>�]�i8��:Cz>{	8>�m�=�%I?��$?5���p̼�i�>W�p=�(
?~q?��N?�H�>=��>�𷽹��d,ֿf5�5�'�Y0����ݼjZ>1�B��,����!>�3������<��=�[>��U>`�>d�G>�7�>�>{��=���=�)>���=Up= c�<�s�=pᅼ�h=�����*1�8��7�ֽ���Y�=��ڽj�)��-�@�?u�?����s��.ig�*��`�� �>�>�w-?���>?U=3)��Y}X��5[�y�d��J�>��P?��>�c7�:פ=lE��<��>���>Eph>��6�<È��4��ϒ�$Ȳ>{�?�G>�S��r;��fm�2����??��=Y�Z���?oy?4a$�(	ּlr!���j��.��\><}=�\�)߉��~ƾ(�T��s�����n5���%=O6�>5�?OC���0�3���_����g�u�����$>�?�-��|���/ ��!�l#�Zg�gͿ=,aM>�X=��O>�;?�+?��=?S7-?��>/�$��>�p=�_�>_q�>� ?7�?UD�>���>�rF>��C�󌳽�T���9��0��<oS1����=X�=��]>�6�<X
=z��=CK=9�4������<l�/�Ue�=�s6=uͼ;�9I>�7?�Y@?�����*��e�(>�j���=���>$x�>����J½[��=j~����?�W?_�!?ls�>�s-�a��Ҏ�Lܼ�?�b-?0��><�f=p>�뾌�x���=qv�=o,"�ga���섾�>ξ�|h���?�b�>�Ry>	N�>D
c?��?��?������P���a�����e.@�м>�]>�W1��p���@�tHH�GW}���a�&��7ؓ���P�!��<Cҡ��3<=�->a/>>��>�wL>ٹu<�z���5��hd���Mn>0!<>٧ ?|"=�{=��:��
H?�7��J���ľ0됾4Z��Fl^><��>TI�=���>�0��:Ki�j���H�����>��?��?R�?�ӽ%q9��ޙ=�`>�)�>z��;�ٽ��;=yt���x>�{�:8���5�6<�w�>5c(>�Խ�l�������Z�&췿^#M��0t��������4q���d��E�+�8�o�Z�,E!�7�K���)����=Qg캁�)�����@n����?��x? ��>�f>G"]�t����%���
����A*/�%����<��#>����E���վ�_��Zu��<���>kY�X;���|��(������{?>2/?[ƾ ۴���s�f=&M%>��<J(�����������WW?��9?�A쾚-��K�[>!�?�U�>��%>����>��B�>4B4?	�-?������/��pU��`j�?���?��??�?N���A�<*������?�?as�>����A�̾����
?QY9?�K�>���/�����
2�>o^[?�N���a>�a�>iŖ>���lJ��z6"������9���8>΢���#h��<����=��>��x>�\��{�����>X.��N��H����V
��H�<d�?n�� >�Vi>f7>��(�d���щ�}`���L?J��?��S?�g8?cV��`����R`�=m�>���>l��=s��9ݞ>���>i辽jr���+�?G�?+��?�PZ?R�m��̿�ۖ�S"������O��=��|=�(>�;����� =!(�=>�<�)�=�e[>к�>���>��>(g>�l">C߇�nU$�ڨ�^���H��<�����bӞ�5C"�!�k�����-��KSپ�{Z��
J��Hd�0����mE)<������=�|$?���>:��>8�>��>�`��	��d��x
ľ��O��
b��\���8�������-��k��2�Y<�/�E{?a%��6�L=�� ?��1�Ӑ>o��>w�b>k[�=�.a>���=Wcs=!#7>X6>�6>���>�=r�>�3�=�����x{�e�L���~������eB?q]��>������������n>`=?��!>}�,��x��g�j��P�>'��'�"��F<i��>��>��<�ڻ:���㠾y+���=ER7>H'D>�9�<�m�����{\�g�>V�l��H]>�o�>3�:?��q?_�P?v��s�>�S?A������w��>|�?�)�>#��>�P`?J�R?��>���=֤b����~+�b�\��q��+�N(2=U1�q�S�׮=���<t�V=2�=%	�m��6�V=T?�x@�6?S$[?�uj>�W�>�ձ�{J�H4{���T�U�>޴����>`?�[�>��>�=+>ș;>al�0X	�N)F�]�>�X)>�I%�'s�L*�;�f�>�W�>R_?�n4?/`/<��8����>��>M�?ȩ*?.�K?)B�>d	>��<�n�տ~�V��T[�f�v=5`�=&�>�>��~<�J`�=�
�=�9��]�J�̬�����>�2�>6��;<ǽx��>���>J�->0ۿ=�>�=��Y��L����{>��>�-��|Ļ�)�uoq=�=1=��ɽ,ym<��D>���h|>;,� ?M�-?�&4��bn�n举�-��Jʾb�>��>;}�>�,?���=�c��]��oj���4�h=<�Y?�Y??�z	��l=	:��5�L�[Ԣ>�?�`>��A�Ց���k�����M��=� ?�m�>��|��� ��|�҄�,<�>4K�=a2%��{�?{�??��� ���,�Y�;/��I�=�"�;��8�%��$0��nL��N(��&��JS���K>�5?���?G3�D�=�y�����]�r��⤾�Od>���<�'9?�4�>�(��žĜ.��?����뿺<�E!?y�+>��s>�?B�>X�??��?1�?M\����?As�>�9����>RK6?�c?�� ?Bp�>��?[E�>���;�	��!k��P	>�^�=Qij>9vp>	�@>���*�o�ֲ�=�<�Ww���,!����f儽@9x����=�rZ>
�>�?�@?�창�B�=��������o�&�+c=�>��O��S�����=��p>�t�>��$?>W�>�ޔ:���q��	�0��=Y�-?��T?��#?�D=��>�������ۢ>Zi��f��s;k�����q�� ��<*<�>C9�>���=,U�>#��?8�?�rT?�qn��iU�����vmR��^Ƚ����^>-�>qZ��	Y:��@���g�F�V���=�'H���g����=Dw�=�g7=#'->���=�c/=�+Y�c�c>^��a��=�p�>[a�>>˳>��>x��>v=>e}Q�4��=�I?���Ag�蠾�nо\@���>��<>����?���'�}��	���D=����> ��?���?@d?��C�@)���\>�HV>��>�/<3�>�A�o�����3>��=�yy����o֞;p]>Ky>��ɽ��ʾ�.��H�i��	y]�MG	>b���v&����Bҫ��%>�p���8/�����YX��N"��ۚ��=h���������[�Ƨʾ�=�?�t?��>,��=/�?�~���Y�n�o����|�����j#�\���<g����¾�{�j�l��7�����>#�L��͐���z�KA*��%���1>��/?	YƾJ0������=�=G>�R-<���k��=��N��M-Z?�j:?Bi�v� �\�����>�}?_V�>4d%>*č����+��>G�3?��'?�Uּ!⍿�����tؼ��?{�?�U?��U��i���2�Z�羳}>�d>/��>���[���ۇ>f8�>ty�>Uه>�-E��ܑ��cR�.��<�m�?�4�|t�=���>b�>�9���ľ�u����ǿս'��=aj�=�hY�zr�=>��x��>���>1�>קԾ�Y����>&,�>�N�ןH������m��<��?L��'>�i>L>��(�����҉��S���L?Ė�?��S?#n8?PN����_�=���>xĬ>���=���d˞>���>�Q�rr���V�?�D�?���?�QZ?b�m��Eӿ/
������������=E�=��>>|߽���=��K=������<���>���>so>�3x>��T>��<>��.>����v�#�CƤ�	ؒ��`B�'�����Rfg�9|	���x�P��	���N꽾��������Γ� �G����8M>��Â�V�@>&4�>]��>���>���>�;�+���<�8¾��O�I��� ��>�tЇ��}��c4�Ȩ��
���	$�N��|@�>����%<�U�>dN=磔>��>-N�>_¾=0��>\�>��V>*�>�ڐ>AW�>���>��=�T�>��=v���H�n�2i9�Z��d=���<?��R�ߍ��%E0���꾢إ���L>0[?��9>��"����3|�xd�>���+U�?p�s�,:��>m?�>�~>�ފ�����c����S"�=I�>�->"�V<��R��l�{@&=�u�>�s��wI>��E��y�>�(&?a�X?~�>ȶ?�>'����)t>j��>��>:�5?ڦD?� _?$W�>��<��r��t��~r���ݾn���2�s��I�=��=)^�=����r� ����)�=��I=�9�p{�=#vk=�>�7?�B�>���>�Q7��3�vf7��O��Y5D>ɏh�L��>��>���>���>.��>��>�"��)���yھ��>hH0>m�[�E%~���k�~M�>��j>�e^?�D;?�ҽ�����ڼ��^=��>� ?�?^��> �V>�u��ź��ܿ�9&���`����>�9�>���<�rҾ�z׽��$>��ֽw�X�3�T�.��>*��>��>0�>�I>��=��>�>>�?>���=��=��0>�5�=�ߦ<��ҽr���D9E=�[���ֽ˶f�B���fx�= ӽf���>(�=�C*?FL!?h��6mɽ׶��?�:� [����>0��>�o>h	>�&�>;W��_��̀�4Ҿ�5a>�??soM?��h��x�<�ZO����~O�>e�>p-�=
��KEw�q����.�{O�>u�?�,z>_`��uP�k�G�x,
����>:~=o}d���?"�k?6о����º3���>�"]O�i"�=�;(>E9:<����(*�!R�9�U�@��P��HT=��7?�)�?p�-��֢=�����3y��C:��´�>S�޽��>�Y=�U%�(��b�\�lc&���x���b>�?�=Y�>@�(??X?~�`?��>9*?"Ґ<]��>�Ӎ>�?�>�>,r#?�'?Z�?��>���>ߓo>��޽m܇�����S�=��P��]�=��>��{>��#>��C>�_�>������)׽��>���=�;�=��|=��=]��;���>�Q?��ֽf��F����{���>y�>Q�|>3��rv=j����A�>���>�j3?||?TԒ>��0���ݾ}2�wW�t?~{?[?������={-�?M����q>̭�>g�[>{ ���: >����7�b=���>`X�>�M�>=��>��f?uf�>$-3?dwо.R���m�J�2�eS�A���H�>�I�>;��=,��3�G�y�S�v�P�g��=����D��<��=Pn>��W>FD6>�!�>�ʻ�������4���Ҽ�yj���>b�c>)?�I�>xsd>w���1G�)]7?X���d1��PM׾���ū.����>���>8��=��?XՆ�;��ܕ��f���>~�?���?7�p?b�S�����p�=/��=��w=�!�� 8� ýu۽���=��>H;���}�2�j�$�">�w>���Ш��󾋰1�b����3p��[�=w����垻��j�J������1쾣
��I嚾x�#�,����ݼ� ��C� ��+~��Wվ[���l��?�q?nn�>np�>��wt����89��c美.����~��=&���Ծ3
��8��x��Y�{���.�>�X�0Ǔ�1Bs��*�7"��Hv�=�(?�A��w�ɾ�++�ߞ>j�w<��/�چ��鎿옿B
���n?!�2?+C��u�����)>Ǘ?���>��>���m�F���r>�t/?�3?����������g|0�ʳ�?���?�jL?�"��}X�;�ܾ}�J�п�>{��>hO�>��W������5�F�?�~?�P.>J����^�8�c�>kC|?�A���8=>��>q)�>��3��Ⓗ�G�;7 ھ�N�T�_>�K>6tg��t�<��`��	�>�D�>��$>�,��Ve����>@�N�N�ϩH�S��E���*�<І?u�� 1>�i>�C>��(����(Љ��.���L?[��?Q�S?Kk8?S]�����v������=H��>�Ӭ>L��=r����>���>�f��vr�e�H�?J�?(��?.[Z?�m�L�ѿ�쟿d�㾄���Xּi"�����>*��������=R�{���^�(>�>�>��t>�s>�H>�Q�>~>g;��_X�����h̤��|q��+��qӾhC����iY��)�۟��s��G>Y�T=O[����c���<���ž���=��?f��>h��>n
�>Ę3>�i`�l��������־[�/�P���֭���=���5�.#/�a*��鮞�1��<��5��>��%���5��>���$�>���>1D>��=+v�=�˔=�|>n>���>�q>�Ά>\m=�\�>Q�=�.����R���5�S�uI���WU?�����־n��tFʾ^r���#>�3?.83>خ�We��}Ā�7��>p�Q��8���
��e�=Jb�>x��>�->Rݜ�68�]M���ar�K�E=N>�>J\�=�W��_�/�[vq�Q��>f9���r&>s�3>̳E?�v?�P?���� ?��>�=����m�>�\<>qǐ>�]1?|X?f1?Xb�>�՚=[P����ʽ�o����S�aaƼ`P���;��w7���*=�A6�_U�=ݭ�=@[j�㝽�==9һϑ�<S�=tE?��/?�p>�`?ƞ�6�&���M�>DC�ƪ=(��&	?L��>���>��>=��>d��=h�ɽ������z�>�MB>��M�Ԃd� ��(t�>:.�=$d?"��>��!�ᅔ�'���u�=4�>VH?�k.?*�>�{���Њ�ͱ	���ݿfUC�[�S����n�Z�=�0>����М�<�6)>O�����ѾozD>6��>�l�>�>F��=	L�>|��>7��>qq>>z�>��->��>L�<0�o�(����[�+V�<+�(;���	�(���F��T����'�Q6R=:W<:�?S`*?j����%��\s�o�#�\�~��=��>_>�>��>�œ>��O��j��`�:����>ʍG?f�?�[���=�j��}�����>:��>���=;���i�?�S&�da����>�T$?y��>�`Ӿ�T2�vY������>Fw= ��1��?��%?�!��>Ѿ� :�<�����Q>)���2�,�����X;�� �"��������r����<ͯ�>{�?F�澿�c>�
��"K���w�#
��Q�=��?�3?=��>*��U���lUC��=V��c�d~�=?b�>Ę�>��R?�?;�e?Mu?yS=?��l��j?Ӌ�>8[�>�Y>�@+?��?��?�&?��(?�Ɉ>�o��&1�����d��=I���u|>B�>��c>���y�>*��>3�+�W��%���!�:�1�=�w)>�c�=��>l�%?�*?��n�V�I>��<��>��=��>R��o̾O�ɻ<�>��>	�k>!?ޱ�>x�{>���R�-�I�޾3��=��?]?0��>��罌t�>!�j���u>3�{>#��=�L%:q����Q� �<F�>\?�O>��>W_?⑹>�`"?�?Ⱦ��4�>�n����#��y�����>��	?~�轿�[�`��}���c����!�>}�
�!�G��[�<�>++>�==g]^>�˯=��n��f�!>y�Q��/�>�P�>��2?|��>�T#>'2־ܪ%���I?tZ����f��&�Ͼ>j��>�eA>���?�
�{}�ť�/?=���>�0�?��?7c?�LF������\>QW>��>:5<�X@���&���F5>��=k�v��y��jO�;�bb>��y>zHʽ2lʾ��ྩ�?�F���ʘu����=,���n��t�[����F����0��{�=�^�;>־��>��="|�=3�ͽ$��\�b�����?�i?+.�>��>�U������"���=������b��a��1}#>xrᾚ ��`׾����1��5-�6���Ġ>_�E��𑿎�{�c$��@���P!>f�&?"¾�����g����=��>l�J:.� �6��Ja��F��ˑ[?>8?�h�>������2>��
?�7�>�6>F����Y�l��>#k/?/1?J���ݳ��w.���&����?��?b�D?��ܽMmE��7����Q���>ӹ�>���>���w��5^��V?-	?�T>h�=��A��d�3�8L�>�d}?Kc,�Y�0>�"�>�o�>}^��}n_�!���k��'/���<A��=���|	,�}�޽�>e�>��>#e#����	��>��ھ�sO��^C���e,(�<�8�)?T� �q>��>5>%*��2������u,�i#<?F��?��W?�D3?gJ�c��5b���a=���>��>~�=&R	��$�>I��>���_�^������V?%��?��?��N?�Pm���Ͽҧ���⾪IҾp>)"���I�=�C������"=�w���d�+M�=�M�>�3�>��>�o�>���>f�x>����Ћ$�����Y���:*�3�)��*�^刾��e��)�m	�7���%�=\F�=�-_�/�N�="�����@�$ m> �?:�?���>���>�R�<���Q���5���Z������X���i��nr����,�+^�ɝ	�[��'�d�Wh���I�>��p�Γ>��>��<_X�>���>�*>cq>V�>E:F>��>��P>�I�>K��>d��>���>2�>�	�=���nl��q9�@B��vn�d�5?��V���Ǿ�7�c� �㨾��D>sb ?��.>�����������>Y<��b������=^�>T�>J(0>��<*��p<f��ə��<�=���>'7>��=�_�{����=k�>��߾4_B=	�X����>�vv?j�|?�=�>a{?Iz�>CC�=(�>�a�>sB�>:ũ>��?�L?�?�ε>j�=��7���,<�S���+��p==1�=P7ν����=�?V>�s�=$�<6�=#��*G����|=��>�`?�@?��>�$ ?gƪ�.2(���G�}���=ΫJ���>�l.>�@�>,V�>5z�>���=�9}��x�4��=�>��>a�����W=ߋ�>��>P9[?�'?\�#�EЇ���ü�ߐ=9�>�B?	�&?�Q�>y��<0.������0}˿G?��.�jn�>�Ӌ�d$�፾q �<��=�R6�� g�t=	> +�>���>�ۻ>��>��	?o͏>���>C,2>ң=#	4>�v�<�<������B<���>X#�<gά=��)=x�i�h=���aɼ������H����&�)?��7?�H���W`��2��'��Y#�&�7=�Y?pD�>l�%=J_�>1�w��Z��L6��~���u�EH?��B? �s��H�=��R�B�H�(X>(
?Ƀj>�𷽥ͫ��ܓ�I�;�0�>��	?j�>/�l�� 9��탿	t��|p�>�{�=`���0�?�lQ?6`�S����!����Zz6�(Y�=
z��pA���	�4���S�,���%�&���>ǳ?,߷?R��9Õ=j��˰�E+�����C��>�]�<Y��>t�B>��2���-�e�k���%�a���?>%�>L�*>�9�>�_B?޲�>U�2?]�!?��6?�XE>/�>��2>1U?�?l�?��#? �!?�?��>e��=E�q�W�$�zƦ��>>{�P�t�=�4>��m>t����_=?�>�3���o���л��4>�@�=I>%�=en>&|U>��?�B9?H���$��̣=&��:�h�=���>u{>84��F89�%ǰ�y>>^1�>`{"?_��>�">�� ���t���b�=�!?ޘ?�s�>;pa��U*>?ḾvSj�V^{>�>�>�L,>co���~?�c�J�t��<	v�>��>�2;>���>f�~?9Q?�iy?��ݾL�J���x��T���}l>����>�>�=���=(+%���T��ne�ʂD��E=�0o��fE�jug=87�=@>>U�.>�>Z�!>lC��)8+=tp��2Y���k��<>�X=�W�>C->���>*h���n���I?���� Y�`���aоgC�f'>]=>�e���?tx���}������*=�C��>�|�?��?C"d?�D����\>Y'V>\�>i0'<��>�<����/�3>>^�=��x����~ �;]>�my>�qɽO�ʾp=�# H�N:���G�H�2=8@7�>��nƊ��3���c���{¾:ʅ���뾁n���ֽ~���ɽ5� �Ĳ���^Ҿ�g��П�? ʋ?`y�>�_}>n��s�Ӿ��̾�+^=J���=�_�9D����Q��W��fϾb[ݾ�&�M�a���Z���*�8[�>��2�Gʑ��~��*��!��C�>��?�þݲ����n��=�z�=n������2���S��`�罫�]?�4?z�,]쾐]ʽG��=�?���>�k,>�γ�����rѰ>��$?U-?�qc��N��Ej���0c�C��?tZ�?�>P?�y��+�E���־���H�>�%�><g�>@@��I֙�ˏ>��?i��>"J>���^*����W�s�?��w?�H��)>F3�>-�?��G�Նž�Sý����F���V>��>2(C�D�?>�A̼�c�=	?8�?H��������>�&꾻�N�5�H�3���F��<Z�?Qr��>i>�P>��(�L���Ӊ��A��L?ܘ�?ҔS?�b8?$`�����h?����=���>ެ>� �=�$���>��>rz辎dr�^��?u?�?��?�MZ?��m��ҿ喿C@Ҿǩ����a>���<��p=~]����=G�'>�2y�	+��RЏ>%q�>�Dt>	޴=��T>�5>�>�P��0�#�@����Ƨ��#3��F!�yB.�;�������R��N���u��W�}�'Ԛ�a�ٽ�1�e&���-��u3�n/����>@-?'�>��-?�*>ѐ�<囓���$�d����Ͼ���Oi߾�������oǧ����3���������>}E=y���U%�>�[ ���^>��E>���=�>`@�>P�'>�x>)��>�>�z�>�u�>U�>��>w�
>�����r�<�;���^�dH$��^??�9L�)�����!��>œ��m>f?�:�=A&� [�� |o��b�>�����-%�vD>Q�>u��>��=.���O$�ޮϾxiY�[ݽ��)>��F=3�0�=�Q���|��1��˜�>�Ӿ�آ=��r<c[t>	�?o?������#��m?5�?ӡ��V�>h�
?W��>,3_?A�V?>?�0y>���<�dB�}�����>�#����~x=�'�=#��>����Rl2�#O�=2�]����� #>Ձ��a��"��=��?=Ms	?P�E?=w >���>��¾VB�<I�.	�ǒ>>�It�=��>���>�j�>�١> +�>�ܛ��X�Cξ󈾠c�>��'>P-M�IP��8�a+�>?�=D�c?R�?���=�G��)]�͠F>U??{Q?	l?�	?��>�Sʽ�� �Y�ÿ���g���s'���H�`l�����.*>
>�>5LļLBT>�K>*�y>�DN>zu�=4v�>�=kC�F��>�Q>�i>82�=N=��^�=�9&>�G>H~�����<}���hK��ߞ��&��<U����L�,�=���z�0���&?51?4b^��=�{Խ�Q.����\�:?�)Q?��=
ټ
�>��<��t��L��V�C���l\?H�a?:|��zp|=�l˽�Pӽzô>��m>}�$>���=6�.��K�����=D?�� ?���>��t�,���i�ʾ�ʐ>��=����3�?��}?�����X���>�Ӫ	����Q��L�Ͼ��&�'�@�%x]���L�>�)��'��>'x ?���?����\>W��񠿁%���)4���>�ӏ���>*�J=���=��?�J�����䭾�;�=eF?�$>�v�>{?>p
?��K?h�+??U�c���>�q>A�?{��>"X,?�m'?��>��>���>��>!�����ϙ��j�=�χ�@�=ۗN>p�(>��5��!<W�>J=u�t�=���=�y2�mj>8>TK>Ca�>n�?_�3?�c	�i��<R_�=\��@T�=lL>Nh�=|�H���A�G=���= ah>��A?H�><C�;�W��L��mӾ���=��?^�?l�?f�v=rb�=yU���,Ⱦ�dv��}�=:=�='�O��ˬ�T���Lq��6�m>i�1>߷�<EF�>�0}?��>�M?�о}`C�"�h�i�&���7=8
���iP>�?>�������6�o�o��Њ�}�,��=��z���><V�<P;�=�"�<ܙ�=��>��m�aT��
f�=���=����1B�>�8~>A�Z?��[>��8>օ��_#���G?�՟��[��Ý�R�޾J��}D>��b>�°�JI?;� ��q��{��xb;��>F!�?�y�?��c?��4�F:�_(W>J<Q>G'<>��S:�W:�4��8`a���w>4�=2�����[�45�<�x5>�ۙ>A^���:ؾl�˾�"�?����;C����=�˼��`��%������`�ҍt�p���5���������h%��:���2R�W�f�z泾u��i�?h�?}��>!I�>�!�f|ƾ����VP�M�⾈ ���{��٫���X��xؾ�o�D�쾹�\�~D8��Nͪ>�'��8����l��������͸=�*9?�ے��#˾^4#��f= n=VJ��z�@������7C轣�m?�l6?s�ݾF���T� �+>/?�s�>��M>vw�75
�R	�>y�;?{�,?b��<Y��'&���ly����?!�?�%I?���"tC��þ=�Z����>0Λ>��?v�^�|s�x0���?^��>��>N�.�º}�#�D�[8?kI�?�J���=0��>��>N��H��=����5J�_ ,>\��=���������/�e(B>�M<>P�>{v�G=��
�>5�ݾ�6M�c�J����:�4����;#?���k>8�W>:��=�h%�_���5��\��RC?�~�?��V?��9?����&�W{����=�q�>n_�>��=k���>���>��վ4�a�����w?���?���?�QJ?��q�f�Ͽ0���'���N���[#�=2�>z�w>[�s�=�5=��Y=�<�>�4�>���>�V�>tÉ>�JA>��Y>a��ғ'�ύ���n���N��4��������W�3og�� �"��S*��#��� �8s�#��vH�j�����?�8��n??}�>
��>���>��=�p�����ľ�7ʾd�� ��E�hL���:��H������K���<��ݾ;Q�>�J�=rK>i�?v>�b�>�}�>!���)�<�u꽔?H�	�<n��>"L>�Fܽ]؇>Շ=2Y�>U�=����Ƀ��
3�F%�$�~�!]4?ӟ�;�Õ��'�X�v��<=	�>r:$?��>'��.����r�߲�>-6+�J!<����#�� �$>���>3~�=�$��؝������_;q~>�#>MW=������սj�u=���>��R=>�H�><^I?�9k?2X?>� >먎>V���)T>ψd=�e�<8�= c�>���>'�6?&�A?Q�>-<�< �[���=���;�Vf�{�<��ѻX�=]�r����<�\��ɽX�D�$>;F�<o9�=�e.=���6� �=ү�>�}=?w�;J>$'���$�C�B�5�=�k�>4�/>�w�>q'�>o?&��>R$�>�&>��2��J��E2��?�1o=W�/��و�3���,?t��ᨻ>�}&?���>����wv>��?�*W?�[??!d?8cI?��㾻o��	�2ԿH�#�2p!����<\@�1�`�2{���,�Uk�ah�<vhW>�P�>�6u>��J>3h>��8>�%�>~�N>0�=�@�=+N<��.;�S��<=��^`q<~I8�$���7켋J��茓��p��]S�rf)���Ҽ�&�>rI?�I��97����Ǿ4�;	��P��>v|�>�[�>��>���3��V���k�K�ƾ*�J>z�?��,?B��#z4>��e�6�H�Vu�>�X�>.�%>jc���f�=�`����(�>^<?zvR>���n[!��xL��<�غu>�������ϙ?��3?����{f�����0������<!E���
���0�7�r�]�+�.���.�+��k@[>��?���?L�������7��洿W*W���<㐚>ik�>�)�>��='f��2l��'K�bH�Nʷ����>|�?b̃=q_�>}\�>�K.?؈?\@!?G1[?%�X<�Ni>9`�{y>c��>�m�=�X]>��>B�)>x&�>ȱ>!}#=��)�_�k�̺�=��0��y�=�s;>�?�=!�=hԽ��,=��=���!
�<8���߸=*�+=�I�=��=|O�=�6?U��>�˾�?E����������G���Z>H8�>B��>��K�>=��>q�V?�F"?p'?_��=o����
������o����>e*.? �i>��l��ء>�y���̒� 񒾯=��'�'�վ�0ž���s�=�$�=m�>$�{>UJf>�n~?�A?��"?y2��~/���u�YJ*�����]l����>���>y�=ܾJQ6��Ms��va���/���#��kD�CF	=1��=e>e�C>ci�=�{>��=���טн�"`<�@k�"m�>��>m?S]>0đ=�0�������I?�����h�4砾�nо�n��>�<>����?<����}�Y
��nE=���>��?���?�<d?��C��3���\>IV>��>1�.<̕>���ㆅ���3>Q��=L�y����D��;��\>q:y>��ɽ��ʾ�0�eH��~ؿ�o�����=	L¾S�,��)���������*��3z;��� I��v�����Y}r��Na���'��u��G���?�I�?��?�*x��M�^��"n2�t� ��X����=g�پ�=k���WоK�澿G�OA��*����Q	�>THO� ���T�x�G+���&�=�9>��/?JD¾I۲�8���O=��>�@<Q]���J��ׯ��-�ڽ$�Y?�9?T�ᾴ����)����>�Y?��>�0>���x��xh�>f3?�.?�� ��
��I����?���Z�?�c�?�>?^�N�]�A�b;���5� ?l�	?#C�>;ꊾ~?˾-�n�	?��7?ŋ�>@=�߃���r��>SI[?N��Wd>.��>���>�+�
���[x��r��&]��w8>@惻����k�GF@����=���>/�w>VrW������'�>��nI�}�R�2��Jb�e;���p?��s9>��7>�
><��)��s���z�L��X$?z>�?�!Q?N�C?�����]T�e�=Z��>ȅ>w��N5�����>���>Z\��1><�I̾��)?��?4��?<�?W��>Gӿ��!��������=%�=��>>��޽�ɭ=��K=�ɘ�3Z=�m�>���>o>D;x>x�T>ћ<>��.>r�����#��ʤ�4ْ��[B�� ���wg��{	��y�����ȴ���N�������;Г�x�G�^���T>�����\+�/�?:�?�'�>:�;>Hl>�T��r12�.��������n'��6"�����}�Ǿ{~��I���Ӛ���3�6�q\�>"��=xAv>���>� ��Y�>>F�V>�'ʻ�?o���i>���=l�>#�>���>��>fz꽱��>���=�ہ�����6:��C��u�h�	](?�}W=�G�=���Tf@�?��<�?3�?6�>�<�������|�4/�>Iƽq�Y�
���HĽΣ>z�>N�=��%��%���f�?K��� >	�>�\q>D�d=�� �IPA��ϲ�>]�>Goо0��=�mw>(?��t?��6?.	�=�!�>(N]>���>���=�=>�R>���>�??�h5?/*+?]��>E�=�Z]��+=��d=�;�5�k�s+������x+���<�.�ۃb=?C=)qg<��k=,�4=0#�����;��<���>�SC?�!�=�=[ ���*���[�~�b���>��[>���>�b ?�?�	�>��>CЋ=�7Խ����*����i/?:ё���#��ʃ�}�ľX�?L����>3_5?ޱ�>�Gf�o�
>�?�_?z�S?�i?݊?#�H���Ѿ���H��#4�4� �TNu��
�=�q�=��Ҿr���R���2�w���J��"N=��>�J�>���>} ?!�>]=�>���>!(�=r">	(^=�S��@�������� >C�įX�nh�;pa=�u)��}˽����y���	���U	�ώ?��?nν�q����F��+�����l�>c��>���>N��>�,�=��"lP�s�[�?�þ�t�>�{?��?bW/�	/>�d�?ս���>�?�>�>\�Y�ۏ�#���NHf=*��>�K?�P>s��7A�27Z����l�>"���Z���?��R?�����ž��4�e�������H4=p���'v�=V�����D�M�����N��?�o؇=j�$?��?YCҾ�0���nھ�C����b�`�� ��;<>T#?I�>}Hh��Z�K�?��
�~ࣾ�:�>��?D	��J��>ܑx?t.l?�?xt�>�;<?���{:N>Z��v�>�^e�?Cb>���>]6?\j ?��_>:�9�2����#پF�L�|��Ø�>C�$>?g=~� <ӦG>q��<Y@>�G��<6P���=��=��<G町�_g>�e>R`(?�?u���ޟ��G:Ͼ���戽��=Q�>�Jj>�bD>D��>�˻>�';?�:?���>�!�����������*��+����>��?
88>�L�:��>�V��ݙ��ݾ�18>�9�R.��3���Ⱦ�׆�
;,�(HK>�	�>,�W>��~?	�%?)�!?-�p;h,9��g������?��v��@�>�ʉ>�F%;@<��]1�R��Zc��e%���<��=�;�Z=�E�=Y,>��@>�(�=v>�=6�=��(��#��=R� =� �>@e�>rC?&�f>���=�g�����K�I?m���hj���sо�F���>�<>����?�����}�:��G=�ʌ�>���?*��?=d?��C�i+���\>WMV>��>�&/<^�>�[
�c�����3>��=�|y�Z���;�]>Cy>s�ɽ�ʾZ2�i�H�Ŀzu���쵻Ǳ����P��n�dŹ��h���D��Xg��D+��}��%5����ʾ����՟�.1%�N��o��� �?+o�?��>E�n��lK��!��#�m�=|�̾�*�������=�舾gx����Ǿ�3��Eq���/��$��a�>iB)�����j��g-�3D����=�E?a����&��������<l��=Y���g�&�1s��M������=�_?/2C?D-g�s)�˫���>�?Q4�>Ek>LE4�a?c�$ө>�"?�? B`�����MɅ�S�`�	��?��?)�M?4w�;�-�݄��(�;�4?Jt(?��3=�S�W��]�:�^ ?M��>�>6��P:���K��a�>T��?!�����= n�>��>b��<>�̾�w��v�:,��>����=Ǐ��i>-�h��ҽ��p��u�=��>�D�����Q�>S߰��:�$H��_�S�T��~Q?'��[^>]�>LFf=�-��S��ꕿ|㙾��/?E�?�8e?]??oUǾxL���v�"p:>���>ˇr>3\�=��Z�x��>Z��>����L�����7?r]�?��?C�:?h}o��z������m���`�Гz>Tr�>�[>�tg��|0�+ʣ����=�<L!�= _�>��>r��>-G:>�1g>Mi>�y����'��x��S펿�PF��Q־�Z8� ��'�9�`�����
��&�Ծ#U_����<���=�גľ{r߽�~��P֬�?b,?G;"?v��>�m�=W?�>5#=v�¾)[��5վ&�1�R?���
���������xr��p��j������o�P,�>�V?<���=���>K��<}�I>q�>�p	=h!<>7�O=ȳ/=�㛼���=��F>J�Y>�	m>�3�<�*�>q�>.[��֒~����5��x�B�3?,��p�^�sD9��A����K�EÒ>Z�?�b>�� �����*�z�N��>/,�?Y��"	�󘽩J�>(�>D0.=��$���мʒ[�)%ʽ��=��>d>B�k=�(����H�J�e=S��>4�����J>���>�?X?݁?�I?u�F>|�>�>�=o�>^3��I9>��	>�@�>!M?�Aa?
�a?!�?�f�=Mw��q�<)ܮ=�B`��7�=Ū��}�=5�1�5��<͍�d�-=���=-$�	��=g�����;��A=)�=��?�E?Ut{��!�=�~<x�%cY�f�j<�>�j�>^ܻ>� ?��9?��>=��>�]i>�>㋡�,> �9v?�MM>�r�6�j��{>��}>�|7����>��5?#��>��W�w�>1D ?��G?�S"?�ai?�Q?;㓾�3)�� ��.ֿȱо��վ��h=~X�>
�������	��vҽ���
�D�K:0��#߻Q��>~�=��P�*W���g�=�!�>�y>Fol>�R�<�y��P8A���={�(>��n;q��<>`������K�q\P�$�������=�ԁ<j'�> #?�e������������Z��E2�>��>�t�>~�>��|��!�;H��
c��u^�>U#|?��?%k�k��=��Ӝ(�� �>�P�>�z:>(�U��<n_���K���Z>l��>��>i�Z�V!5�c"F����R�g>��_��b>�?��B?�?�0=��;]�/	�\K�^���v_c��ڽ�M־j+F��U��6�6)�Ne��p��>t?iE�?hӾ4�#<|Ѿߛ���"j�om�IͽVQ>��?��4>�#���k�.�D�V�$���[�>���>/P�=�i�>�,#?��?��a?#w??b�VM?ה�=Z%�>���>��
?+�?��>Čr>=�>�	;=��0���
�Pd���^<�̼���=��*>&�$>�e�<?�=0AB=���<��?�{��'҅;kDe<b=���=L��=�k>	PB?�/?%���M����Tt��y���<� �8��>���>)��=4�?0��>�W?�Z�>��1?b��>&]�����ľ�=�_�?�6^?L��>�+��v>����Z�^3��Ur>��콘Ӿ��#,R��9���Z�I��>W��>cz_>�7u?4�<?u�"?��߽"i/�g0e�3���ʳ:ꁽ���>t�>}�=9�ܾ�3��/p�@W���$��S�yR���=�Y�=��>X%F>�y�=�?S>��:������{��<�g��	�>�ʥ>x	?�W>c =���8����I?�x���c����0NоU~ ��)>ƀ<>k��n�?Q��\�}�����@ =��k�>;{�?���?�d?��C�qH�8�\>��V>�T>�33<��>�vP����o�3>'	�=z�6����;Ŝ\>�x>4,ʽ��ʾ��㾊�G��1����o�Y�D�,`��&p�������k���\h��n���X��V�H����l���펾&���c��۾�-��+(���i?)In?�"I>1�ͽ��G�ɂ6�v�ξ'�=�o��ٸ��7���Mi,�e�1�Q����������hO/�k�}������>�tE�m덿�Tw�ݑ0�O�I�~�5>r�1?g;ϾH;�����r�<��>���[�-����a��Do����\?��;?z�־y|����]�>)�?���>�4>7����~�|�>ۏ.?�E(?V#�9m��'d�����:�^�?ꈾ?�<?�	>�f<7�=�Ə��;�>{�?ؓ�>(ҁ���۾pjN�l� ?L7?w�>��Ct���l���>�V?8fJ�(�f>�1�>�Ì>7�����KQ�c���IX����:>��<����}X���*��y�=��>�2l>(�T�������>�����K��A���@X�~=��?m���5�=6�L>By�=;�%��Պ�����K��?"L?��?�HS?Qy2?���N��e	���ml=%?�>f��>s��=_��b;�>��>����Jq��t���?]��?W<�?~s]?�e���п���������C�<FY�=��h>�����a>�:8�>����ʶ�4�=���>mN>��Q>�-�>S0%>7���}*�m ��a>���+{��1��#��Nh��[�ʾ�� �����k:��K���b�
,F=>�ݽ�|H��>`�)�t6��w�n>�!-?�1 ?!9?���=v�>�׾��>"��m���-�%F羇��f`I�~�[�h;f>�0M�Ku�=��R����vs>4[8�;i�>��9?E��>>��=4����7=�H�>]�<�<"=aV>iȊ>'�=���>�+�>��>��>��k�ZY��Q�5������k���<?�*{�- �=�K������=�n�>	?��Q>Ў�Ҩ��ڄ��Q:�>��x�B��S3���H�	ץ>��>U�=��vP<TX`���%�n �=%�8>��>�`=I�h�ET-���<o6�>j*�5�t�W_�>X��?Yɋ?�E�?���>���>�U��L��>�2\=fCw=;��3I�>�gi?s�M?;�?�@>?�y=a��S��=ڙ+>�'���i����n��=���=��M>+��>qI>j�>�5X���>W(�=�?`��É=�W�=.��>ʶ>?7mb>����@���LS�>_\���=�T;E>z(>&�>/�?��>�lL>�o'��f����ž�]?��>f��Ҏ�'h=>(#�>�{H�Y�>KoJ?���>�о<���N�>�|R?v2 ?��l?�BT?���� ,�@#��Կt:i�������y�>8B>?��ч=�[g=LV=��u�H��1�=C�?�ǎ>�>.�?�U�=��>=�X>�$>U4��I�>I*>>XHĽ� �;����c=�� ���a��z[�J�!>b�	����'��Ak���*�=�0?�?�;,=~����ƽ��;$u��3�>�w�>o�>'h�>��o=h9�1�X��X�Z�9�}g?BZY?���>m�D�^~�<���[+��c��>��>ۻ�>"�!<*bu�js���y����>F\"?n*�>L�I�KT�H^�����F�>uf�G<��q��?$;?��
���þ�JH���n�8��-=��؏Ӿb����8�X�M���T��A�7�����w>�N?V#�?eY������c��β���v��nK=��c����=��>��>#l�b���}/�
����=��B>h��=�e�>c�6?_�#?W�;?(��>�o?�����%?ܦ!<�e�>��>N?��	?h5�>�H>��O>�Y=�y�=���ӌ��2<��.<��>v>�~�=��A<׿=O}H=CE��V��
���j�����9�:)��=�Z=��=q�7?3XC?�μ�ۺ�����H苾�5｜�+=e�6=#_�>L%ܽ=��>�Ǳ>A�B?M��>>m�>������5�����R����Iֽ�?D�`?š�=$�W���>ր��:���{�wz>)j���ᾔ]�bB���U���������>7h�>�{�>e{c?�Y?Jo+?O,U�'d5��2��X��X���`����>I�>���=�c����7���w��85�i�~��=�+���-=��% >3�>ד�=q(h=���׿�=��<<Y:�?���Z>� �>y7�>��>g<�>l͡�.���	6I? ���O�Av��C�˾f���>��>>8��-`?(F���}�z�����<����>=�?���?�d?Q5@���<X>M�Q>-�>pf <�B@�����q��6>�^�=�q��r�����:^>�΀>�뽽��ɾ��߾�t@�zʸ�d'c���ٽ��d^����������da�)UȽn����뾅��1_!��H[=�Ή�q�̾�a��`e���?�͑?,��>�$�:`A�eX-�����=߆��ߐ.�I!��qܔ�줲����g�o�$��|D��N���ᾉ�>��V�N���|�a5)���ļ8�8>� 0?�}ʾI��ӂ��h=|">!<���w��L]��&&
���W?C:?���O����U�l�>��
?�`�>��,>����*�>)�4?�,?���eW��q���Y��D��?
*�?��??�nN�~FA�G�����h�?�t?��>oK���u̾\��?n�9?p�>���5�����80�>�-[?N-N���a>���>�O�>���#����(%��6��ZY���U9>���i-�+h��8>��b�=�Ҡ>��x>�a\�ᮾ���>Q���+N��QG�QE�F��!��<�P?�W���a>6�g>�f>�&�R-���鈿C���BM?!q�?\Q?b�8?���y
�y��a�=�R�>tͫ>�ѫ="<��W�>l��>��律�o���r]?���?�?��V?mn��п^��Y�hI��$>s�>'vd>Nlp����=*s=�ټj�W��70>	Й>&&�>yt�>y�}>�sg>��*>���V�&�}����-��B�G�����X�K��$���B����3o���D��"��h�G��uF1����4mY�>�1�R��=_C?�"?ߨ"�y6�)R>"dY�g>N����(q�����ؾ8cоk�6�����Ф"�`����Z���Ҿl�?��=�h�>0l>����h>-��>+���[f:>95�=�#R>�:>�_=��>V$�>�_�>�P����>+$>2��IR��Y$>���P��N����7?bz���=�h3��t����>�>;�>lD�>8�n��N���!��>��#���#�4ӽ�Z�v$b>7+�>X��=�:�<��
��彭�L��P�=�1�>�5e>M#�=i$��*R��=�,w>�#��	->�Q�>v?�s?;�K?��v>�?l��>]��>.כ<H&�>J�>5+�>~�A?��d?�j[?���>/�=>����Ӹ��&=KB��h=^MνT=>I!���<���N��K>IJ_=:�=��3=���:�3�;;�T=�?��4?��W>7/>��k�!9��c�;q�;��<��i>XlG>�z�>(�?V&�>3CQ>L׃=ro���վ��ћ�>��>��Q�5��b�<��|�>U3*���?�?"8>hVW���_��1�>`�?ޚ(?ڄg?�=�>"������o��տ�|�a������������=��&���3�z2�������D>��>s�?���>��>���>Z�=���>�>�=���=�Aw������ m��h
��J��7�e��w��L�/>/c=>���IX�HAI<���=��=����f?3�$?<���y���O9��4��L�ɾ�Q�>��>[̗>k�>�����뾤�x�y�[�u"�(�f>�U?��3?�Z����/>a�[�Ն�5�>�4?��>�����)����"���D=���>�Ĭ>(�>��&�UE�u$�x^�ޘ~>���<	����\�?oU?�S˾�;����է!�.���ܡ=[���x�b��,>��73�Z4�����bI�«�=�|?~_�?�}1��)�;��ξ�����]~������6F>80�=��>�G=>Z�n�^V����,�N��ڵ��$>���>��A=�>D??�s5?�M�>a��>����?��<<Q?���>���>�?CC?@��>ٷ�>@��<D���� ˖�ex	>�F=7�Z>/��>^6�=~˺�f�#f�<��H=Ws.�H=�<���V��=߱3=<�=�-,>��=��"?nE)?�b���H��A�s�u�;��{���ɜ�>s>�S�=H=�?��>I^ ���>F�?��>â��8Q�v:��^���:��w�>��i?���>a�P�Xs>�萾��:ξ�;ʻ`�a��Ew�S����վ�ȩ�{s>�>�>���>?&P>�?^?��D?~ 0?��K�:1��D�����D]=(/p�vP>���<Jﺒ�|H�*�m�3�D���
�c܋=��C��{= �A<�F�<f�>�"�=�>>l��<�}ǽ��҆>���8&�>��>��?�?d>�e>�Ͼ�w���I?
����j�i�Ctо�T���>h�<>w���?`��/�}�x��KH=����>~��?q��?�=d?�C�i+��\>�RV>�>�/<�>��vz��K�3>�=!�y�c���}�;G]>�By>ˢɽ�ʾ�1��H�s�n��!]��<��OG=����qŁ�7�R&0��u��c���l����<q	�/��W6�=ň�=�$R��z���?��?x4�����Ҿ��=P���<>
�s��=-c���Ȱ�o��a�����y|�j�Y�p�9�M���o�>JHU�|���{�p+'�������:>�&/?9ƾK��;����t=�%">+a9<��>����G��?��W?�9?�*��E��k�佋�>'>?�I�>D�,>ᐾ�0꽇�>�2?$,?���VV��̚��W1����?�r�?s4G?��=-�M�re1�:��Mxa?�4&?���=wc9�;b��wO�<z�?��(>	��>�%�,Es�m�7�[�V>h�c?ރ�^\�=Py>�bK=4�Y�"��	�	>v������,�>�l��C��ٽ��lý_�M>��>��]�.��b2ھ~��>�P꾝�N��H���������<�?w�48>�i>fJ>�(����r͉�=���L?���?݁S?hr8?oN����h���w.�=�ئ>湬>�0�=��U՞>��>[n��}r�V�P�?sC�?���?SZ?ԓm���ѿ������t���,�=H�>�oV>[���j��,�=�8=���P���&{�>#�l>!�n>��s>�0C=���=�U�����S�������K/�%����t����'���O���޾%�Ծ�о���>���e=j!E�����j
m�����=�>}�>GZ�>�L9>S�
>t�X��X����1�j��'	�rs��p3��ɾ�]<����f�B��������=t�(��G3?0g8����=�;?D2���=�[�>�H�;Acd>�_�>�"�=kr>��>b��=�>)"v>�c�=�p�>�S��T���l�y� ��&��<kg�>����L �#:>��x�3���Q?;:<?�T�>al$��i�� ����>ǎ�(s���y彌���!m�>�9�>'�g>�=/њ<�;���v���qM>u��>(9�=�=m��m��C�����s>��>0P׾a��=�Zu>(?�Uu?	6?���=P��>w�[>b��>���=h�K>��W>o�>�?C|8?��0?4��>lX�=�<a��*=V!:=��@��fI��P���7����#����<�A���G=9�=��5<x�[=�p)=�ɼ?��;��=_[?�~?H��>���>����Z�nM�w���9<�눾�f>4$R>�&�>��?��?��>����
ߵ��ҵ�-�>�sc>z��偿�|�<֥�>�g�>0�'?�KD?�z=����l���
>Iu?Y*?�?��>>l��=��>��b@�����&�@�'����;^0(>X���%
��>�5`�V¾G>>GU;��F<n<>�]�zc��Bv:��:�>5�(>�r�=�#�=L*��m^�@	���	>S�f>y}�<���;TK>�
�������Z��;�Z�=0�<ڬ%?�-?��.���>e����,��־�$?v��>�1E?�%?~��=M�nt�S�{���q�?��?R	�>�� =!>g�=����$6��_�>	���T���s�>������>�7?h��>���>�Ӿ�kq�m���t�s�>H=�咾�@�?g�C?���୅�����[a�~��?����S��5p�n߾d.�0<�Q��)����3>�~��<N�?y��?Q
���0$>D��Z1���I������/\���r�Sq>�7���˾0m��k��
�&�
r)�Mn[:O�>�_��W�>���?c�(?�X?��M?2-�?���/z�>Q�>/P?W0?e]�>��>3�t>��=�z*>�p7�D���ې
���Ҿjِ=?N�:�� =]�> �C>o�=j��<�<$y�=E	��$��3z=-��=�j�=)9�=��V>qa(>I�?��S?I�d�1B>.yM>�3v�-౾�>�:ݼ�j�������mG>U�>�R>�?n]�>J'K<L��3�ξ>��Sc>Y�;?�>U?\6.?�RO�}�>��)��E�C��>'�u=����נ��nZ��Y���I&<&1?CXG>H�ƽa[j>�C�?>:?55?R�R�J���7k�3�$�D>�<`D <��> �>Q7>��޾s�6��s�Q�_��:����]��a<-�<>>9>��>>�+>��j><��<�4ƽv���v =v˽��>�>��?MI>�^�=�㟾���q;?�ԧ�nfľl��w8��z�ξi��������ľ���=�x¾-փ�P���)�'�̎�>�$�?��?��E?z���F�<�?&>Z���N>YLT����9������=��P<�=�:�x�A��=��>�@?J�#�������K��<VѮ�:�u�lt�;i�;����������}�ѽ����ɶ��
R��7OG������� �^��{���R���x�?��Y?{�>�����=�=o���־"���Ц��
K�Hg����z����������1����5���h��3����>�d��j��z�i���%�uK�?�]>��>�Ȥ���9��K����g>���>3V4��p�@X������_?;%?ҿ��H��F0����ʼ!!?��>J��>OZr������r>�}#?�@?�'F; ^��Uj��D|���?x�?�_\?_��=l�C�j�-���Ӿ��'?�1N>g?�c
>Ǉ��^�.�IA�>9[?��?<Տ�D����?�=�s>e�n?R~R�|��>�x>ao�>V�y�������p�=>�ub��=^5�i,ֽ�� ��c/���R>��?���>y���l.����>�A꾓�N���H�s��[���R�<��?��5>�i>B>'�(�����ω��*���L?Қ�?9�S? l8?Z^�����˱��ŗ�=���>�Ҭ>A��=�����>P��>�f�lxr�����?�J�?q��?�[Z?��m�����y'~�'� ��"о�K5>�Y>�}k>ZF^�Hc3<m�=�'>@t.>�W\>PrE>�;�=\P>�J�>.>����P�|�6��.}��qß�v#�޾Le�������T��a�ξ~s��FG�dć���)�c���2U2��&4��n(��r̾�l�=G�>���>�~�>�m>���>"�����iν:4�������������=���=���p�[���z�a��<��	�*	?�l����}=���>A	��_�=���>z��<��	>�[�=���;�u'>8>2��=���=��$>e�=���>��A=յ��'9w��5�h���xJ]���+?;_[��3���m6����YF��J��>�?G�s>�'������`��>�>��4��w�h�)���>H�>���=Yg�<�����s�b1�yI�=��>��=g����9�����
�='�>x�վ�:�=F�u>X�(?Ɏv?�J6?�ޜ=$�>}a>�W�>)��=ߺJ>��O>Wl�>Y�?��8?��0?}��>��="�a��=�{9=3?��R^�ى��Dἇ�,���<�0��<=%�_=T�;��`=<�L=9�����;�:=M�?G��>؈�>&�>ST���c�#vm�U/�@��<wc��8��=���>E�>A)�>J?��>��Ls��
qh���>x<>��X��u�lP,<y�f>���>�c1?�s?E�3�&�f�3�� D�>�M-?O}?�C�>��=�N�=���=�+�
��e���Y�� .>~�z>��i>��=�m�����=�#B=�O�=�=���=�s�=��>��B>�#�; ��>���=��(>��=^
��Q��T��C��=է������ǽ?�9��{��Vd�0,=(6o���B�)�<K*�=�X?ٗ-?��V=0�q>��O��U0��ľ�?Y��>��??7��>KF>��&�tz��;u���	����>���?t�>ND�=��3=oJT�Lz6��<��t>�[�+=hE�>3?x�O?��"? �k>+݌�Iz\��}���y澊j3>=}Z=�˪���?�&>? � �L����Q܁�^jҾѥg��$�"nľ��0����t�Px������l���&���?	��?y��띐>��G� ��P#��=H�]�Z�V�r��L�=�	�� �,h�-�쾣E���j�j9�=V�>`R<�Ơ�>�z?�	�>�>q?�J?���> �=x�?�m>Մ	?��?��?P0>���=5���<����)����RξF=/&>�
�=
�=�*y>���YW�`��=LJ�=T$,=H��$�=�B>��=�W�)�G>�G�>+&?�?�g�i��>-�r��߂��S����>W�p=jO������=*q�Ҍ�=�>�-?�=?��5>�}$�3��� ��*E>�H?�<?&�
?�4��:;:�̯��ݾ��>�8&>���ﾀ�b�~��0��@?sO>=�ѽw��>�K�?�?���>���������1��]�ž�:�>��}>���>��>���>m-�1P��4|��:X��H�"���ц�؀%>��>��7��>"X�>x�>N��*R��#�&�ݽ��u��
�>Y��>�?���>ð[=����^"���;?E���s�;䋽g����/���=���=�Ƨ����>ك��?��Ѱ���6����>��?`+�?;6?�E�\�򽾘k>}��=�=��>�um�]�h�����nQ.=�A>agɾ����>��>2\3>J��(P��譝�.L�:�3����}��ⅼ��>�9�(i}�Ľ���~tB�Xѽ�e1��V��3��1�	�f�#�}*۽��Z�����S(����?ׇ8?"|�>D7>ۼ*����)Pa�d�[�����j۾e����9����p���[پ��_��/	�ˠ�>Ps���⍿4pV�m-1���5�mx)>	�>u2������-5�Ms�o-m>%|�>8�b��Ta��B��P�=�a|?�J-?�v���۾K�ڽġ=-g+?�a�>^V�>�)���<�u7>$?��4?�Z> ��ɋ��j���Ѽ?`��?�<[?�Ҡ��z1�4����a���a�>t�(?�ܩ>a�ͽbm�L)�\��=ۜ\?\�W?� ��K��7I��5?G1�?��	�H]v>)͢>���>Brؽ=�:���O= x>�鲽�R;=��K=/�ͼ~f��*���H>���>T�>T�ľ,������>UA�W�N���H�<����1W�<�?���5>�i>�@>I�(�����ω��*���L?Κ�?ʊS?�k8?�]�����ݲ��E��=���>AҬ>\��=�����>���>^f辰xr���t�?mJ�?X��?�[Z?��m�CIտ�3��Ј��Oؒ���F<�_�=���><J��j=�H=���=f=iI�=|>�x>�=>��>eA�<R��=+����<����6���>I������d���a=վDa�6���h������vu����4�Ŏ�q��4C��=j�X��a>&V?o�?��>;�=9�>� ��
t.�d2*��� �]8��t�@��/�JVk��2>�����4þ*��׹��b?�=���>�6�>!�1=�Ol>z��>��;=��->��=5!�_3
>,�'=F��;w�B>���>6==>��>�y�<����&�����p�@��6?{�M�4��(�<��v���V����>ˤ<?���>b���/���S�z��>�ʼUZk�
�����Z��>	?Ή>T?�=O��= �r��m}��>u�>4=��T������]M=�d>c��>G�Ծ�?�=S�u>b�(?��v?��5?�d�=�j�>maa>�h�>ؒ�=X�M>LYP>Wć>>?�t9?�=1?���>V�=N�`��>=w?=��>���S�i���f�ؼ��%���<�.�_-H=S�s=K<��a=�\>=�ʼ�B�;�=Ep?W?ऄ>o��>�׽P~g���c��Ӿ�<���ʖ%>��>$��>g�>g&?��?������j����>h�2>��k�����"�
>3��>I<�>�Q?m.?[�?���H�t�L>�>�?��2?��?	�8>r-�<��=Cn ��⶿/c#��d��$N>%t�=#��<�����{<&�>���>�@���@��x�=�~0>���="G>�ި=!�p��>�<����82�8Pd���ͼ����w^�u/�D�t���:t�P�xo��ؾ��I��:�=@Q$=q���q]�:ߺ?��9?�6"��=:�l��!�h�žr�>X�>dZ�>^��>�>R�4��r�޷^�_��c�>�?���>2;���=�/��n� ��:��Q�=���0O>���>�E9��?��e?�'?!�>L�q��g[��������>	�*=(���k��?*�[?b�	��]_�z���o��^��<�3%��l��$ ��T��(�_����Ȭ�����A�=�T?d�?���p�>��2����K���B��'���?�UO>�}��6�9���g��U���W����I��=%��>�0Ƚ.?��w?�7�>�c?&4[?�?(�<>7�?�+�>%?B�"?~�?�"=A`H���>�xL�>	�;<����<A�yx���e5>��>#�=�j�=�T�>c��=o���{�<�X>�ü���g i=a�;>��H<�0�=8�=�;�=��?|�)?c,���g�=���I�R��TӽF[-=�Ͻ5���}������ȅ=Df�>/��>�m�>#�=j���%�y	���}>E
;?Ɂ#?�96?�v�=�>�.���Ͼv��>�<"��z�`<���RP�*��7����?i�>��^��r�>�sy?�?��
?�3���;�'c���0���c>��>U��>�?�tC>�����M��4��A�e��(��9!�:U�DϜ=:�=`}t��Z�>+��>�g'>vZ�"���p���X�9�����>\� ?�8?��>��;~��n	4���B?�Ě�Bf��
�m�+�ľ8q��Ϙ=����PJO�c��>`�I�kX��~����\2���>p��?F�?jQE?�<�C��缪>�g=B7�=_��=Y8��+��Tņ��U�=��@��r��
9��fY�=�,�>�y�>�G=�.־�ݾyϗ��T���ꅿ!E��Y$ɾГ,�}�Ľ�þxp[�<e��u;��d�2���0�־��?��$��7Q�[���n��#^��Ǻ�?f�#?I��>�J�=�(I���оvxy�z������U�?�E#��8ν�a������zT���妾w���: ������>�~��ŋ�����C?'�-�]�c�}>��?�L��\�龑�1�����Ֆ�>�ҏ>!g���j�k���ܖ���x?�(?��پ��վ	���[�8<0�?6��>�ˇ>���d�S�*�o>b?׶A?���<��������+��?6�?�9c?�!����M��x��56�[�>7��>ߠ?v���]i3���y�~=,�y?�d?����4O��GJ���S?ۖ?|�`�G8�>�N>���>T�ֽ�������	���䊾�༡eI=����Jþ ���\#=��> �c>�����ɾ"��>�A꾐�N�تH�z��>��1U�<�?��05>�i>�@>@�(�����ω�*���L?ٚ�?B�S?	l8?^�����j�����=_��>lҬ>���=�����>���>Hf辤xr�O�w�?�J�?���?�[Z?�m���ӿJʜ�8���8��I���=]b>!��_�"=��=;�<Ճ-����=��d>RL>+�E>�ރ>�5K>��&>CI��n
"�삔��F��mW��)�q=��*\�]����_�+7���Ͼ�ž>5�)�Ͻ�g=bu�c�-���<Yľ�AU=ر?�<�>�[?��A>���>�%�3�#�ۢ����Ծȥ0� 	��sl�|b˾93L�^��=燑��q��I4=�����?w�9=�`=.�>��/��B�=��>g=�=�M�=��=W}<�LM>@�;sA@����>�>�>d�>�э>�#�=B��5z���5�fN�\Mڼ��-?vU����0��S!���Y�>��?�Y\>�(��-����i�r5�>��W��Lt��{��7��8��>��>���=�=G ~�z�/k�pJ�=E8�>�>�'7�c����νה�=���>�־F�=�Ez>�'?�Yu?416?��=�O�>��W>�.�>�m�=jR>N�c>�l�>��?	�5?.a1?�+�>�7�=~^��# =-V=��=�'�E�Dۨ����������<��E�CB="�K=��0<%N={a-=d�¼�<�Y=L�?�-�>��+>���>�W"��d���r�N
+�����N� �2��=�1�=�e�>3�9?��A?�p?�+`�bmξ%�M����>�
>C�u�Q�a�/U�= Sy>�>�9?D"?�w*����V�����>3U7?��>��>A,�=F�>��=���-�̿�jξV���A ��倽���=;!��ֽ8�=Mh��&��mj��kya=M�L>��X>�ݠ>��>&�#>���>�PS> w=�cc=�Kx=:!>�5�=�,=+EU�����f	=9=�^���� =����Ͻ��3�6�9C��?
lC?����� ȽR�>�+�"�K�k?�/?�?6)?`��>p��n�k�
�d�C[�n�>���?�,?�Y8<�h>0�@�����=�b�>ޡҽ,�<m{�>�H�����>�L?�^?9�O>gQB��\�Je���eǾr+?�>:='���l�?�_Y?z�-���I�a�)���t����F�ڽ}���l��t徒�����
��ӣ��pJ�^�=� &?K��?�u��>����ିѓ�AJ+���޽'\�-�>n��=�;2�e�R�e(V�_d�<X>=�F���(ڇ>�T~�}r>�8�?��H?�<?��N?p�M?�Oa=��>���>��'?)?=�>�>���>��6���U>�՝�"I���������7�{=[�=Y{�l(=>י>uF�=��>i�M>!qt=�n�������,����=Y�=�>���>�$�=D~?Ad'?W����є=�8�=��n�I����K>� �>�v.�+ΐ�؜;	�j=��[>���>8Y	?�Y>����2�6��2��=�)?�-\?8W?K��2��>�A�U� �3��<�ɀ�2a�*B��K�� ����fT�>W �>T0>��z>�?^�4?�+?������sr���Xi<p=W�>~
�>��4>'�;��6���n���^�&^@����S�W���a<j�>]�F>��H>��=ay�=3�<���z�#ƻ|�����> ��>�
?K�j>w�=ز��V�
�EuF?2x���+�Ќw�c7���_��a����=�#v���`>W��;�v��a��/���?�*�?J6�?�%?��C�z���s�> v�=ph�>��>B���_���=�|	>F�d;0�ޝ#��:㽫Žw�0>K,�=KGi��lܾ�#�̦��=Iz��7�=�.��m}��I#ҽ�����Լ�`�,�N��鿾��}�?1�������4��2�D�gk��|o��o���Ɩ?6�W?M��>�0>i��Ǿ�;߾�<=��nJ�(@�����/����O�����뷾�%ʾ����V�I����*�>�`�i��3�q�%�f���$9*>Y?�þ�о���j�v�R>S��=]�ž���d�����Z?q�6?�0辅{��t��(
>�H?	��>qF>�v����� >~�+?�(?���;a����<���d��>�?�̼?�mL?��=��3���a����cz?�Ͳ>�}e>�
!==���y=��>�f?A��>&a��4$u�(]� Y�=��_?$����>�&.>�Ok=C���LaY��?���	;�/=��z�>M�S���!�����ܔ��`M>b��>���>c-����?�+��>�@�a�N�p�H�5��q��V�<�?^���5>i>�@>!�(�����ω�[)���L?���?��S?l8?�]��7��󳧽y��=���>�Ѭ>���=����>���>�d�|xr���F�?BJ�?L��?�[Z?�m�
��X-���(���{¾���<
@&<��>UB3�*�v=��3=I{=�̑<��:>�e�>�%>Ag2>�G�>n�>���=�W��L�"�c?�����#�0���cY��ކ�f����r�/���V��:���������f���	�"e9��
ȽV�Z��G�>N�>��?vռ>q2漎T�>�Qd���@�F���*��G�<�����������������=X�\�h苾��W�Ԣ���m�>�L�<��>���>�M���=t�>j��=�B�>=�\>v >>"P>ɟ<�u�,>ŉ>%�>�=3_�>���=�b��Rb��_�9�Cp^��ә��>?)�Z�����3�D��M������>��?��s>>#�4���"�l���>� >��	c�t�R�Ky�c�T>�>h��="i�ūi�ys���ɽ��j=r�M>0&>`�=��W�X�-���L=��>ZM־Q��=��y>`�(?�w?W�6?:�=��>j�a>�4�>+��=|�K>��N>h:�>�j?s�9?�]1?��>�f�=�+a���
=	�<=T�>��oU�����!����I'�!A�<��1��tH=��v=�<�k^=s=E=��м���;;� =L�?d�?�Ps>�>]�}�n�g��Fm������c�]k���RD>�QW>It�>�A?��?��>��Խɱ�:|����>��K>H�{���p��^v�/Q����>�Z?��6?��J�pw��=�=C�>c?�<�>Λ?��R>\E\>��$>&a��Dп�]�/����[�S�9���</oH��r����F����n,�@�<��>>�g�>d�w>��%>3�	>��>,��>�D=�>��=8n � �D=���߶�=z����͞=ݪ!�>b�<jS�!���ǽ]?��a�f���x��o��%�"?��<?h3g�`�)��+���Ǭ�x��l�?�V)?�B?&�?�օ>ZW(�y�^���m�)j۾��>鹐?4�>��"�\->��R�NU�.�`>���>_]��fn�=�DC>V�ýX�>V\/?�z�>t(�>o�*�������R��h� ?\j=	ӟ�	��?kC?qP"��?g���B��/����(��K���r��������B��$�ݛ�<�ھ����Q�;!�?���?p��r�>�􌾂˫�.%����W�ϽJ�}��>�	���Z�)l2������΀���˽�U�>쥾q�>��}?��A?؀a?8qD?�GS?럥=�T�>�n�>G�K?��?���>��N=(f�=r~��ƾB>q[q=� Ӿ����hƷ�e�A= �=u򽍷'>�g�>��.�h�:����:�к=_ߏ�%� ���h=�i >7g=S��<��/>P>u�	?�;?����-Ž�|�����<p�Ҿ}>cm��4��渾Pn��S���O�>��*?Ay?�V>�+��l��I���V>>�?u�m?m?��彪���K����þ~F>r}�=��;ڼ��C�@��ƺ��㾼�W�>��=�7=ddb>"�?b?T֘>~�>���ßo����XO�=���=6�>~��>�~�>�@ѾC;�'a�S�N���R��6���h����y9�>e��>W^x>r�=G3�=�=Gp��=�=��1j}����>y��>�N?�>��Q>
倾�����8?CeK�(���g۽�g���)��D�=��#>���� �>c����?��96��p�@����>�>�?�?r|?�0�k����>M$�>�->���= F(��O�=�3�͋=aA>������þ���=�H=GA���ǽ<���B?���ĽWֻ��^��!�=�AҾ�1��J� C���*�I���y��sM�.G��{��\��M	����8��.l���L	����?�>?L�>�;v�N�^Z�k����?�A��Qw���
���p�Kx��=��K��hKо������O�F3�>����$���dp���Q�"��9^=��J>�Ǿv�&�	�C��Fu��۴>WE�>���/�A�Z��~�=PZ�?&,?�ž�
��B�����W7?-h?)��>�@m=bJ�=�f>n��>	3?�du>$?��s~~�W��?��?�`R?�H�o�`���<��z��ƥ�>�n�>	\�>rA�;��Ҿ�ჾw�l>F�E?�*?����ۋz��pq�^	�>z?j�F��m�>L0�>��=(g=�a�<�=����9�����e=�%��
h����c��T����]>�`?�(�>'�n�9���>�A꾙�N���H�������TR�<�?��5>7i>�A>=�(�����ω�r*���L?�?]�S?+l8?T^�����0������=���>�Ҭ>���=�����>���>�f辑xr����?�J�?���?�[Z?�m�B�Ͽ,������(� T~=�].=ƙ+>g�as���<-MH�Ws��/�=��t>�K>�J�>��>��>�Aj>k�����*�U���������*��e ��L� m����0��v���b�����*������q ��p=e��=��<�
�&>�׾�i4=&��>���>�r?7�>��r>v�=3)��Z�rB ��<���6�y�!���оQ����C<��=HоR�;=׾���>��>#@>p:�>�mO>��>犉>�>�c ?�;�>X�=@�h>��X=.s�=z�=���
�=�/�>٪�=�0���ނ�T$8�M�9�p��<��G?\mk� 좾�.�����6�����>}�?eG>�� �Q���<|t�e�>�e���j���ֽ<M<I��>�l�>j�={�꼵�1��,F���=}��>�C>TWf�����[���y�=R$'?8½Up�<��0=P0?��b?"�8?o{>R^I?�~6?��>�H�Kڭ>���>G�>�mD?/�-?��4?���>���=�<l��<>������=G��m�?�����W*����=�=��</=�MA�z����=�1 =ς >��];���>r�K?�H�>�Ӿ>�о��l�]�D��|
��,=���XT?��A?P,?�^�>��>��v>c�"����x?�q�>��;>��C�	L��V�f���?n��>�hQ?�@?Ȳ �[����=,=k>U��>n�>�o ?gA?�I�>�f��T;��mڿ�em�E�F���>�а�{ѝ�z~��_�jg�J�U���A��G�=��>o�=6H�>�?K?��5?��>'�t>�\k>{�	>�5N=9V�/��#^���=[i�=�&ֽ|)˼;/<��<M���@��;�&��}.��Q���?�q?�2�LX��;i�us���ǥ�X��>o��>���>�u�>�:�=���FYP�a�=�_TB�y��>�4f?���>}L3�;�=*�1������i�>Ӱ�>�;>�l��m%�\��x=�<^��>�V?�R�>����^�b�l�Z��Ô�>�r��W��=(�?���?��� ��iS��#Y�s�c�1���ϛ=��s\?��4�̉]�+\}�'�o��1+�{��t��>҄�?�R>}��6�	���w��!��+w-�o�E��nW=�ȫ>[�t>ʌ>7�����O��k�܁�b�;5��>l�L>�.�> M�>0c?SM?R4<?;�/?��\�?� �>�>�>�7�>R"�>��
?d ?'У>��>�t=m�+=��+��ͣ�TY>��O=�A�=�T;>�{>�Ba<8V>���=#Ѽ�"m�˥��}1B�K�s���=�
�=��=4X6>[�?�y)?��z��������`��=�!�>��>2���
v
�\�k��f�>Rh>י?�6D?�?�>���=�4˾?���T�̾�^� T�>�:?���>k�.>M�e>t]̾��g�>��>��	������]̾�Q�hZD�IJ>�?�>�$�=��>Pjz?�1`?�6?�2.�����à��5K��9-��*1���?�t�>l��=@�K���y�����D����J�&��ب�)�R�4_r�� �=���>8��:Ť>6m>D><
��3�=`�}>'d�>�9?:�N?���>�G�>�w��m�&�I?���(�+���$о���/>��<>�z�4?p
�Ф}��ҥ�9�<�\��>O}�?إ�??Dd?�C�����~\>�V>�^>��"<�p>�=���酽=b3>���=@�y�9:��)Ή;�I[>��x>>�Ƚ�Vʾ	s�<G�Ae���"M�6�	��0��t���<���o-Z��w<;Ws��u��5ҾFh󾯢Z��l���jA�����������E�?mrl?��>��>I���C�����3�s>dp����������V(�'$վjo���6��O��)���2� ��>�!�z��� Հ�+�3������^:>A#7?�c���]ľ_��_u�==iV>ӹ9=%^�鄿�{�����
�H?��4?V\侩<��0/��%\>+�?�9�>��>>�}��OJ��l>xe%?��&?(�= ����A��M�:�ķ?���?uD@?G�?���;��7"�/b��<?{�	?��>@-��_0̾uu1��(?��B?O�?3�ž{{����-��>�+?��A���=3�>��>�p�=
�7�
��=� ��nv�Y�M>q�"=����]۽&�M>�s�>��g>�C���r��5��>����9D��qB�_5���m=)?�fϾ�>�/I>r[�=�|(��+��g������I?��?��P?t�5?�E��e ��t����	=o�>��>�(=,@���q>���>D�Ӿ�e�^�ﾝj?���?��?@6a?@]��Rɿ+���|��E]���>T�= �<>Ʋ��E��=�|�=6�ͼH.��!>��w>�(F>�}�>Y�b>ɓ0>x�>�ψ�dS#�g������-�+�������2�T���ll���n鵾b�󾵎#�{�K�H���C���~��B̽�r�HM-��?_(�>/t�>�7~>�~a>��;���-��5��*���;�l� �< �n���2����a ��^�q�������>��>χ<�8�;���>� "���=���>7��N��=�>Ay>פr> �9>��|=�R>X��>M> �j>/�>:Ř��i��z���D���)L>�
M? ���ž�k[���T�U�M��F�>��E?��>��վ��S�+�j���>=ꋽ_�
�g�:=���=��>G��>X>��O=$�m�U־ 
����^���>0�o>u=V¤��콥�,=��?3���*=Xf�><?|-N?*8?L��=}��>7�?�<�>�ñ�u��=�݃>{R,>�6?u&>?b?�3(?���=]z���,�"��NhN����<B�m�G7����{�`ɽ�(I���=��H>]P~=J��<a��=���_�����o�>K�+?;*x>c@�=xI�u!E� �J�d5k�}��<t�����>@�?�#,?35?c�m>�w�K ����4�ճ>&.>|��V��- ��'>H�>��c?E
 ?�a�=����c+8>��1>�ʬ>oW?���>���>�f�>'H;> ��$�ӿ��#��E!�|7�ߦ���;��9�^{<� �1���د<v:Y>BY�>�2t>��G>o8#>�\4>H��>��@>d�=[�=H �E{�	
P��@*=R���	+;�oa������<��s��������/��:�vl��B�üMt?Z?�6+�C� �v�L�K��ux���> ��>F��>�<�>�A=P���uO���1�3G$��6�>�Br?�}?k�-�ዚ=j�&� ��<x��>u�>_K&>cA������c�"|=���>��?��>$��� �J�"�_��t����>�7v�E����{�?�C|?7 ������$5�v�y�)�^�Ᲊ���ӽN։����[l��bS�S8ԾM\S�P��7�켼�>]�?�F�=��������k��sG��쐠��Y�;t���8?��?l�>��ٽ���s��\2���Ҿ5��Ӡ�>���>��?m|$?��t?��?<�?ܤ�;�$�>��>�M
?� �>sq?�}?l�?��>^��>�፼��`=�����f��!�=����A�=s�;��=.2>'p_>z]Z<�>�yb���o	�-c�+�ͽo�<�"����_>�4 >rN?�� ?(6d�A8(�~�=.4 ���A>Eh>1>��F�C���FSͽ��>>�#?nG<?���>Az�=w<)�)���#ʾ��� ?p�F?{�?�M>�G#=�A���=���>;0�> ͡��r�����f˾�oy�T��>��1>�~>�Ɍ=�^?�oH?�!�>թҾ�kW��Ӓ�4$E�kqz�/���?��?l8f>�)��Y>���a�(����kg����]}����=��=��伹 *=J�D>R�=H�=8J��[>�+�-=޲�f��>��>FW�>���=���>������ھ�xJ?㎝�ܸ��H��/J;�(B��6>s ;>i��4�?5��\�}�"���<�Q��>���?���?GMf?��/���X>w�V>��>��<�,4�*��)m}�1>���=y�n��d���!�*�W>(�y>_Ǻ�<�Ǿ����+���ƿ0h����߽��*�π��L��k6�Ϫʽ��E�ja�"x�W��'�&ž/�T�?%;�����ƽt!K��9z?�p?\d�=���>��P���Ͼs̳�WF��v�脟�u���w'��[�N��s�ȾT���E��ᾬ���*��>I�H��#���J}���)��KǼǾ9>|�1?1F���'��5��9W�=Ƚ1>�=�澕���b_��r:���Q?��6?>�����[��9�%>^�?�W�>U<>�l��*��U>��/?��(?M��7��@v������(�?e��?��(?��\�Z�a�!��4�J&�>�1?m1?�M����׾�Q��?�_<?Xh�>Gɩ��,��ȭ���>0)<?&O7���>��>�
F>߇	=�������=���翽��`>��&��>�J����2=�#�a>���>�>yo?������>�A꾙�N���H�������TR�<�?��5>7i>�A>=�(�����ω�r*���L?�?]�S?+l8?T^�����0������=���>�Ҭ>���=�����>���>�f辑xr����?�J�?���?�[Z?�m�B�Ͽ,������(� T~=�].=ƙ+>g�as���<-MH�Ws��/�=��t>�K>�J�>��>��>�Aj>k�����*�U���������*��e ��L� m����0��v���b�����*������q ��p=e��=��<�
�&>�׾�i4=&��>���>�r?7�>��r>v�=3)��Z�rB ��<���6�y�!���оQ����C<��=HоR�;=׾���>��>#@>p:�>�mO>��>犉>�>�c ?�;�>X�=@�h>��X=.s�=z�=���
�=�/�>٪�=�0���ނ�T$8�M�9�p��<��G?\mk� 좾�.�����6�����>}�?eG>�� �Q���<|t�e�>�e���j���ֽ<M<I��>�l�>j�={�꼵�1��,F���=}��>�C>TWf�����[���y�=R$'?8½Up�<��0=P0?��b?"�8?o{>R^I?�~6?��>�H�Kڭ>���>G�>�mD?/�-?��4?���>���=�<l��<>������=G��m�?�����W*����=�=��</=�MA�z����=�1 =ς >��];���>r�K?�H�>�Ӿ>�о��l�]�D��|
��,=���XT?��A?P,?�^�>��>��v>c�"����x?�q�>��;>��C�	L��V�f���?n��>�hQ?�@?Ȳ �[����=,=k>U��>n�>�o ?gA?�I�>�f��T;��mڿ�em�E�F���>�а�{ѝ�z~��_�jg�J�U���A��G�=��>o�=6H�>�?K?��5?��>'�t>�\k>{�	>�5N=9V�/��#^���=[i�=�&ֽ|)˼;/<��<M���@��;�&��}.��Q���?�q?�2�LX��;i�us���ǥ�X��>o��>���>�u�>�:�=���FYP�a�=�_TB�y��>�4f?���>}L3�;�=*�1������i�>Ӱ�>�;>�l��m%�\��x=�<^��>�V?�R�>����^�b�l�Z��Ô�>�r��W��=(�?���?��� ��iS��#Y�s�c�1���ϛ=��s\?��4�̉]�+\}�'�o��1+�{��t��>҄�?�R>}��6�	���w��!��+w-�o�E��nW=�ȫ>[�t>ʌ>7�����O��k�܁�b�;5��>l�L>�.�> M�>0c?SM?R4<?;�/?��\�?� �>�>�>�7�>R"�>��
?d ?'У>��>�t=m�+=��+��ͣ�TY>��O=�A�=�T;>�{>�Ba<8V>���=#Ѽ�"m�˥��}1B�K�s���=�
�=��=4X6>[�?�y)?��z��������`��=�!�>��>2���
v
�\�k��f�>Rh>י?�6D?�?�>���=�4˾?���T�̾�^� T�>�:?���>k�.>M�e>t]̾��g�>��>��	������]̾�Q�hZD�IJ>�?�>�$�=��>Pjz?�1`?�6?�2.�����à��5K��9-��*1���?�t�>l��=@�K���y�����D����J�&��ب�)�R�4_r�� �=���>8��:Ť>6m>D><
��3�=`�}>'d�>�9?:�N?���>�G�>�w��m�&�I?���(�+���$о���/>��<>�z�4?p
�Ф}��ҥ�9�<�\��>O}�?إ�??Dd?�C�����~\>�V>�^>��"<�p>�=���酽=b3>���=@�y�9:��)Ή;�I[>��x>>�Ƚ�Vʾ	s�<G�Ae���"M�6�	��0��t���<���o-Z��w<;Ws��u��5ҾFh󾯢Z��l���jA�����������E�?mrl?��>��>I���C�����3�s>dp����������V(�'$վjo���6��O��)���2� ��>�!�z��� Հ�+�3������^:>A#7?�c���]ľ_��_u�==iV>ӹ9=%^�鄿�{�����
�H?��4?V\侩<��0/��%\>+�?�9�>��>>�}��OJ��l>xe%?��&?(�= ����A��M�:�ķ?���?uD@?G�?���;��7"�/b��<?{�	?��>@-��_0̾uu1��(?��B?O�?3�ž{{����-��>�+?��A���=3�>��>�p�=
�7�
��=� ��nv�Y�M>q�"=����]۽&�M>�s�>��g>�C���r���S�>{���5���@��nF�l���ْ��M?����? �5?JS�>�0�߽������KE����*?O��?��G?PV<?��F"�Rm	>��"��>h	?O��cbǾ��q>��?n�:�&�`�AK-�Ӈ^?���?.^�?,�Z?t��&3Ͽ�-���L��|���p>�K>{֯=�q=��<�˽��	��S��򫤼q��=;Oj>t�>Ȗ�=��>�E>������ �����\��]�3�yH�g� �Q�I�9d�nJپ�:5�rr��[��1�����݇=�p��~i�<2��D��qƦ=ӂ�>xL�>���>��^>�qF>v����S۾�
�����d��Rwﾗ�����V�����_h�:ڙ�9�1�E=����>�P=��6=�>�j���`m=���>�w�=�&>&W�=Ê�=�q>> �(>[I8>�
3>�SK>�>��[>�}R=�愿9W��s4��>��r�;��:?�}�\ڒ���4�cž�����p�>�{?*�M>��!��3����t�$n�>���R�_�ǽX��b��>���>���=�>}��ʼ�{�i��T�=4��>��>�����v�_)&�NE{=5g(?�"Ⱦk�]=d�>O�>��2?�?�>P�k>�Z?���=Tj5�a
Q>��>`cn>[,?��?X?��>�%0>RF8����[��=���0\=İ¼,f�	���5=�\Ž䙧�e�Ӽ5N����;��l�<9�	��BO�=� �>ԄC? ��>�=pOv��'�Qo�qֲ���K����F6�>~�?./?��>%a�>B�>���=�en�?��Hs�>��=�8:��~���<����>?�?��b?��#?"f�>$����h3>/��>|��>��?��?�J�>,*�>}�=��
��ѿiOK���J�'�:�<�'�ᱽh^��<�x���ݴ�����LC�=�q>OW�>x	%>ɟ�=/v�=��>�([>_@�=�|�=�ޓ<�G=��=�"n=L��=��=_Ə��g������E���#�VX��Y4�<�'�;Hɗ��;?�`?rnS��g�юN��0��9��5�>��>��>���>f]�=�[�wA�f+4�$���; ?��k?���>��<��ȴ=q������;3��>:�>d�L>�`�d���d]����=�B�>�?	-�>�2����V�8s���鬆>����Z����R�?X�F?���UϾ�ln���W����L����5Q����b�/Rx����uk��n�����
?���>��?�G�=�����E�����dx��Z�^<VX������n�>���=�oἊ��ZV�nj����#�1���>ʨ?><�x>*�0?5}&?�*j?�K?z�?%���7�>P�b>��>J�>���>�
?��> �:>F�K>��=����i7����F����=h62>�S>bQP=M˓�_���B��}0�Q��=�}2��$���=�̇<ŷ+����<�z>˧*>�A?��&?� 1�=�������Y�y>r�>hs�<�>�=d�Ǿc��=:3�>�9?GP<?5��>�}h>� ���u �ҡپ[��=�*?��(?��?��=�|�<��޾�`��!��;\˴>6>M�?�ݑƾ�Ů��C7�d�=��9>��=~�H�h�~?���>>�q>�G� ��f���M%�3�0�^ަ��� ? ��>-H+�L� ��F�V7t��*b�:�Z�'<�ص��m>�e=����l>"�>�=������<�I/=�U?����=���>���>O	?��>�rq>l��D�*�E[?{�����|��c�Ҿ
�q<�k>���=F����K
?[
�6*��㎿Rr�c��>[n�?��?kT>?��� {�K��>�]?>���=s�=����L$=K��60>�Yq=O�L�0h��Mk�=@�>|͏>P��=�����Y�;k���̿���,о	x��'_��;��C'�=K�Ց<=/@�IϾ'��:��S���ҽ�ѷ�B���$��*^��b?���>Ȫ>�Dr>�ej�B4��0��
���M��<��9���*������Ė�j�ᾐ}3�@9����E��B�>޻T��x��b�|��2)��<ּ�3>��.?n����U���n��Ox=%>�"<x+��z���)��_
��W?"l9?�1��f��n<��)>�?Ɉ�>�(>�Y�����2�>�4?-?���BC��0ي�K-/��>�?L��?�7?z)��N:� ����J��'
?�X?�5	?��n�h{Q��q���?GnF?���>������k����j?x�0?I����V>���>!s�>�Թ;	Q����F���L�B^��Ap>�O�<��b����c�c\>n�4>�A@>|H���̾��x>����AP�L�7���9��]���� ��:?A�3��៼ʜ>�Ӱ>�,�������|��,ʥ���2?�H�?Q�_?q�"?�p�����Tٞ=d>'+>��>�x��7��ø>��>,?ѾA�]��ܾH�+?ވ�?�b�?
}3?r����ȭ�q|��gY���������=��=<0S>�m����=�=��=�n��k >�Ԑ>"CK>��R>١'>�@>a�N>K����6%��	���c�� G��)�Ȝ"��z�9��� �����������{l�����.�U�Q����	K���N�+���si>���>���>���>i�7=���=Ƒ��Z|�=�u�a����!��Ѿ�8�A�ľ�]R��L�����ѾLM<��Ͼ�/?�=v��=�o
?�!������>�R,>�Ɉ=S |>�Z)>�;�>P�g>�=?>ܲ�>8�->|�=���=!>����y��K��r��#P����?�a���}���U�|9���
Q�P~>n/�>��*>��#����o��$�>d=�f�8�C�X�<=\��>+b�>D)�<V� ��?�;�>v����=�L�>wF>��=�>ݽ\'���߼��?}���9Q�>�w�>7?L�W?T�(?�9���>���>םN�')½a��>��>���>۴�>��$?)'S?��>��6>�o��l��<�ef=��^�9�������@�f >���L=��<��=/��=�%;=4t=)ٽ&����>Z�=b��>�]9?��j>x�>��5�2�(�h2?�0����`=��漜n�>���>�?�� ?�l�>�e>����������3�>o׷=]�v���i���|� �?��>WI?uT+?k�.P���=�>-��>4B#?��?�e�>���>���=���zjӿ$�2�!����;*���;��<���M��D<7f�-������<��\>��>�p>:
E>��>�:3>}Q�>�EG>�ׄ=$�=��;Ͷ;��E�!�M=��}|G<	Q������MƼ��������I���>�[��)ټ�?��?�)��錽��h�&R��ͫ�T$�>���>���>��>��=����U� �A�lI��N�>H-h?�0�>�j8��"�=��3�o�U;��>�9�>k�>��g��~��ɗ����<���>F�?ua�>�1�I�Z��o��
���>v��� ���1��?�Di?���7����;�wJ�����)��)>�%�8���JP�$�X���5�D��xz�q�j>MҲ>pX�?������Ȯ�����皿��o�ku>Ӝ�;=��>��>1�C����Z�4�澋����=��>���>$<�>G�*?E�?7+2?h(?�?<�V��k�>/S8>�Ĳ>u��>4\"?�v?|X?���>)&�>�mt>����������9v�=�
��F��Rp=iS�<�G��<!A=�в<����;;��X<��{<~T<�\�=�0�=�w>C>ˊ�>
cB?��M"����=�5>�r�>�>��=�1G>u���0��4+��g�?t�E?B�!?�}>	�߾�b����os>�{?V�"?���>�~=l8>�2��)�ս�� >x><"K���ʾD
�7�����)=��h>�?*=쪅=�DZ>�}?�7>?u?.���1�Av��+��Y��Ɋ��	�>{k�>�1�=�޾�86��dq��_��14�I�{��(=�U=S9�=`�>�:C>�$�=G�>!��<C��~��!�1;N�]��>�2�>G�	?��`>�̖=2᩾��<?sT���:6Ͼ<x�1�=�/�>b�/>�@׽�I'?���J�������`�>���?��?2a+?o��X��y>/��>/�K>��=a��GV<�V��p%6>fC^>�Ƚ��þ���fu'>�S>�Eн�����
�$z޼�洿��=���9�%I��
��c�M2ȾSW��ANv�A���.$V���㽦̉��諭�hx�����n��VϾ�%l���'?�>?��D>� ����"����ܾ�\ܽ��<������������׾6L�W��(����?�0C����k]�v羰k���P���E��n�}����_?�r>�z��i߾,F>s�>�?��F�v������=�ɽT��?.�5??ڎ��������	����1�>�e�>�F?���<XI����=2F?�\?!��=(l��^���n�>^��? �?N�:?��J��D�l�]*�0�?J?c�>kj���V;t2	���?�7?Ƅ�>�������������>$�U?��F��e>���>7y�>@�ŽA�����D�풾�xм5�<>V�7�7b%���o��B>����=�@�>�Wg>OY�X���+�>r���]�'�F�U����/��&�G=p�?z�Ծ[�#>��}>�,>r`�����Ā��u��@I?�f�?KP?�$:?���O�cĽ�#=<�>S��>g��=����,`�>��>��Ӿm�l��?����?˯�?$M�?�S]?w�m��vο������ؾ������=�= �0> ��%�R>��>h��8�:"��v%>O�>u��>REn>�ȉ>Rl2>�� >i����H%�څ���ܟ��L��(��-�E�A�>>���X�-�6��,m���ƽ��Ex���
L�� ��!�0�H��S�>��'?�'�>-#?�OI>���K.�̂������(���u��A�Db�J��)�ýn��~1>/*�����V?��G��>�B=)�1�>�8>���>6�=_+��=�C>V�W>��[>���=�=>ڱ�>�t�>`�7>�}�=,�>$�>�y����Ni��%>��Q�hT??$hA��2��J#��a����"�'Ŗ>�!=?�6>�k@�]����*�����>t���\�h�¬���/\>)[2>���>�X!>ZP:�%n� ���f��h=LP>W��>�=�Qp��[��)�p���?���>�ܾ�>ۛ�>Z�?��T?�s�>���>F�?'�"?(˭>�\�>��>�`s=}Q"?5�]?|�?!��>�$���vR>>�n>ǵ����ܽf�0��G<���E�^<a���c�V���/=���=�;H>a?>q���dR<&��=\U?�$Z?D�>t�>�\!���4�=aV���W;��
?��I>��?��?�~?���>��P>�_�����5���潙����>	Q>��i�$j���۽�>��=DL?�S?�j�=eܠ����=i�>J�?M4?��H?� �>ɾ��ھF�	�<�̿}���G5���齒��==`�F�>��s�4��ߢ��9�v��
>5�>t$�<���>��>_�R��>Ԃ�>��&>�8>1W�>��&>)6�<��<?�m�r,3�Z�����ʽ[.�=�>��~��=N/輀���!w��h���g�=(?�?�2�=<K>�i�m��{n�����>5 �>l��=7�>
�ݼ���Q8_������X�Q�>�*i?�� ?���w���y��謔=��G>�J�>�r�>��=W�˽4����=&�	?��H?��=�6����j������=�t>��<"��u�?>��?�!g��#���׈���#�x�8���m��@-�g��v�f\4�-om���G�,NZ>�/�>�!�>+�?k���$�V�qվ�n��cF��^E����>�?�>>�>3>�N��C�%��"F��zľ�SG��zx��>߯�>�� >�آ>�w�>M	9?�1?@<V?s>#��>1�>�Y�>>{�>`r$?�>?�C?x ?�� ?�ι���;(<>���A�=i}ս�=�=~1>���='��ɕ>���:��)��<h��<k��'³=�Q�= �!=?�=U��<3�?��=?ǖʽ�2�L?�AK������R�x>#�=�� >Դս�@M>�m�>3=�>I`e?��>L�%��2'��u�]3�u�u?ubD?� ?���<н�=� ��Px�l 	>�޷>*� � �4�������/� �Pq�>�=�>_ߐ>�9B>p�b?�iY?a�&?�<�=^�E��d��'i���u�@�2�ؠJ=�V<�o�ʎ	�a�1���a���[�L�Ⱦ��.=�.�a�>h�=\�.���>qӬ>�[5>U#��������_�,��3���G�>�;?���>.<�>�=G"O�����5�E?޷����	� @��lʾ^���*��=��!>�r���>��%�����*0��>=����>{��?Y4�?�#f?��1�.���p�=>�;I>��1>a����:6�<���7�9�1�A>w+�=n�_�-j��SW=�aC>w+�>��뽯ӾX�y�:��﻿�oj����X���k'��q����+��ؽ"ǘ�\����(��ꐾ�~v����������'��uY�P�������fW�?�KG?L�>��=���W9���M����E���;4�о���_..��9-��W������@�)�ܾ<�۾��>.�`�W��c�^�>��d�=	M>gy0?jm�����������>'\V>��q=���o�~�@���~n9��1T?��U?��1�Q��#9�U��=�{?���>-�w>�s/��iW�T��>�.? q?q��=/����v���^=��?�ݮ?q�@?uR��TD���1���?7�?q��>�F���Ǿ��὎?�9?%��>)��]��b�����>�gZ?[�K�nJ^>�Q�>s֖>������B���l᜼�>>:�����]�i�T�>����=c�>�l�>�&V��A���Ƌ>$�ƾ�b0���!���
�s�/�ݽ�9�>����x��?8�=F�U==�K��c������.T�0c?#ٳ?	@?L�)?�䔾�Ӿ2nf�0(#>*�>�n>�2�G1��
>x�F>_]��p�8 ��?�>��?�?cza?؉q���˿?�������y��.�=KM�=��C>�b@�`F�=:3�= �޽$�J��>5
X>P��>��>[J�=2��=|��=O,��w"����V�n��)b�M��n����/�꾧T���/�K<��	���h� ؗ��|��}��4�C��fb��n޾�a�>A+?}n�>Ds>O�:ք�x������[2���#��j�'9��5�����<�`>�'Z>����M�Q,��(]?�y��&��=}"�>;�=�e�>]<�=���>Lܗ>V�r=�i�>�>ׄ>�=MҜ���D=��X>���>��
>FV��Ƌ���O����=�`�sE?!K�gu��Ax/�~���(l�ޗ�>/�!?m%>Sh2�%������Ô�>~:��{�j%���7=8��>��?��L=�.�Ou���Ɛ��X�[/�=�>�>�
:>?�x=�i���ҽM��I�I?�3�!���;�>}�b?�/�?��}?��?��>%�?�@?P�>���>FG?�c�>J?��?{��>'?��>cǽm@l���Q��\�����=��ּ�νL�=���<,�=�C==4��=ؘG�9׭=��=�U=<~>��>F|5?��>�
Q>\�پ��T�=V��c޼�l�>	!��m&�>?H?1
 ?s��>�޳>���������㘫�3��>�I^>��p�e���?u���G>h>%�D?n�@?Sl'������>�m>f��>zNV?��;?��>��g��nᾁ����ӿ� ��h�;ؼ���C�"�<@�k��ͼ�2�:1�2�(!�T��;ߐJ>u��>��z>�u'>!�>��*>r��>_x>t��=�D�=�e�C)%<ӔL�[ �<a��;�u��6����;���,�{���ؽ6
z���S�B#��$����>K ?��>U���ќN��	��׾�/�>�W>}�>{Ә>�#�� �c]�P?��,�Z�?�q?~?����T�Hɽt�0>u�>��]>hu�=U��=AA �1���t_>�	?l2?���>u8G��o��φ��{��ʄj>%>4���E�9
�?�v?w���]��9D&�<�7�9�Ҿ�n�dC��3��G) ��5�>?M�t��Až��6�ߗ<>��>&��?��B����<+�_�������4���-��6��aZ>�w�=�ե�8�߾���Jkξ+5=�>�]9>�_�=��><��>Mɹ>�V?&3�>d��>��_� �>LS�>�?k��>J"?%J1?
�?���=Ōf=ĵƽ�8��I��@H���WM>KE>��P>�ؙ><�#>��>7�2>�#�=���>��4��ͽ~[T=Z�>�@�=p(S=�|�>��?I9B?�,�ī��n��M�l�U=&8�=�f=�{�;v�eqo>,��>���>H�7?چ\>����3�;Pc��7ؾ>H<�z
?V�@?��1?��>־=�u�
�;	�e>��>�)����f�����������>���>}=>c>��f?��??��?my)�)�7�Fh��X�$����!<K�>��y>���=�Y羦�S��󋿲�i�a�%�s�S=������=̯=���s<�S����=�	E<�I>�Hܽ�x��s�W>���>���>���>�K6>LvC�	6�mɾ�5'?j�[���S�����Ⱦ�zҽM�=�5=l�&��՞>2M���g��?��j�M�[�>��?�g�?q�u?�?����Y�>zi�>V��=�C=D��S�ٻ�ڽ�%>t�>�܅�=0���[�=J�W>iW>d���y8���о`�B�5�Ŀ�*p���ܽ�;I�n6ؾ� ����ۍ�C����ܽ'�ܾ�r9������/#��Dg��T�>���������?:�`?&|>گ�=]^F��8��r��<��=�B�^�~��Ŝ�#3#�Ӿ�%ž���������
�Υ��ƾ�8�>�Z�PA��e�|��k(�z���@>8x/?��žu3��IX���h=̤%>"��<Otj��������<W?n:?���:8�����>�?�>�%>e���P��
�>}O4?�z-?%����U������+]�?���?B�??�]Q�0�?����E2����	?��?�Q�>g���c��0����
?��9?���>K|�����Q��KM�>��Y?�G���l>9�>��>�w�ÿ���9���u���u��{'>�rh������X�V�2��l�=�{�>b-}>�_V��í��*�>�X����?�R�/�g6����������V>#�=a��<�#���oD���������K�z�9?>�?�_?p�-? LȾ3 ¾���:<��=,>�q�>��#>k�,�+5�=��t>�ɾ�]��r�W2 ?I��?#;�?��Q?���#�Ϳ���������N����A>y�=�^>���<�ڒ>��M>ŋ>�&I=�)5>7�>��%>6�>G�>�>08!>SĀ�i/%�Z���/��&G�����> �a� ��#�{Ⱦ#g ��/>��:��T�r/߽im��:����g�4Ѯ����=b��>���>ȧ�>�e�=X^R�K�����C~;�g�RX�������g�����l�0��_x=�O�=B�������)�>��|;,��;Z��>�{=��=//�>�3>E��=R#�<@~>��U>�`�>#+>��?>0-�=.�=���>'��>?���������B���V����<�(O?����d��
�Y〾�s*�H�>^�9?gf�>���ڝ��H���L�>g�1�}5���ؽb�<�)�>�?0��<�55���Ҽ�QϾ[8/�u�;<��>��=�^5<,���+��gQƽv� ?	���aF	� �>�%U?�y�? �s?�Q�>X%�>T�'>\2?Χ�>�o�>]ȗ>�Bk>�@?-b�?=5C?�]�>�>Q0�\�Q�ܫ=�o��ݭ�*��bɽ���=���=)�z�|��� !�#���J��^~
=T����A��-�<��>ֲ:?�ȕ>��X>�e����I�>#O���=���>`Z>Y�?��>�Z?�3�>z�?�f0>�D����䢾"��>��>��v��&����=�.�>�?>��c?�O+?�)/���O=���>�>?�?lWS?Xe�>�;}�Zg����޿��<�ב�>q�NRS=�6�=qVf��=S�?���q����<y�>�G�>�qq> Z�>�QO>C#>F��>-1e=�A�=&4�=y�]c$=l�;�󂻄���&��y�v\�����B��;v���|�����J�UO�H��>�G?�ܣ�Y��=Fi���쾠2�lĔ>��2=�e>X��>�`̽�����n�4
D�;�]����>PNg?���>�|$�;>3;������=<M0�>ܘ�>%�6>��=���Mf�ñP>:�>��E?�5�>V����h��	���37���A>�[�"z��#�?��N? ��/v�������*��S�r^)��/��du��O&�%J��2��,7�;5�D�#�^[>���>$��?����!X=���-��q���PR��1�=4m�>��>}�	>'F񽱴��i(�����7Q��B����M?�>�>�y@?��?a?q�?��/?;)˽<?r�>�e�>���>��?�V?�>��>�Q�>�ۢ=O4ļ���o���˽N��ek	>, />�H>�>���=��->%�6>^����Қ���=]$�=,8>��=dy>�)t>*�*?T�:?�	Q=��[��2���j��'�>�b=���=7��={n���0�>�v�>,�,?�,?�G?�y����"�#�R�S�������03?`?$��>3�S=+�=V���yL�ó+;��B>f���������Ҿ�OU�q��>�^�>Nb>X9_>q({?�8C?2#?�,�/�-�M�u�
Q+�9]Ѽ8�;���>n��>�`�=߾�3��t��a�L0�� !��k?��=uq�=)W>�+>6�=�`>W�(=�p��<ҽE�<%};W�>1�>��
?p/^>e�=4R��� ��UI?X⠾���R����7Ͼ'V$� �>�&:>��U5?WW�*�}������=�xw�>�>�?��?��d?�B�I����[>�WU>��>��<�_>��`�7(x��/>�h�=viv�ᬕ�Z��;i[>_x>��ɽ�9ʾ��l*M�s츿��}�C�ᙦ��l�?-����l�k�d��i�~��@U�M8��������	�.���^�J����i�������?w�?��}>[������d.�N��d��o����DK�(�¾	&U���Ҿ����UվL�&�k�X�������j�>,�Y��&���|�$�(�s펼��>>k�.?�vƾ�������wd=��$>�B�<Q��O���䦚�w�
���W?��9?p�뾙5������>;?�%�>�$>����S�뽀,�>�3?ǜ-?ͦ�����+���i���h�?7��?��??��O�j�A�>�J���5?\�?��>�Ŋ���̾�`�?��9?���>�&�9g���3���>F�[?�8N��mb>U��>V:�>���g���w&�)@���l����9>��
�����Lh� 0>�K�=j�>h�x>�"]��	���*�>�X����?�R�/�g6����������V>#�=a��<�#���oD���������K�z�9?>�?�_?p�-? LȾ3 ¾���:<��=,>�q�>��#>k�,�+5�=��t>�ɾ�]��r�W2 ?I��?#;�?��Q?���#�Ϳ���������N����A>y�=�^>���<�ڒ>��M>ŋ>�&I=�)5>7�>��%>6�>G�>�>08!>SĀ�i/%�Z���/��&G�����> �a� ��#�{Ⱦ#g ��/>��:��T�r/߽im��:����g�4Ѯ����=b��>���>ȧ�>�e�=X^R�K�����C~;�g�RX�������g�����l�0��_x=�O�=B�������)�>��|;,��;Z��>�{=��=//�>�3>E��=R#�<@~>��U>�`�>#+>��?>0-�=.�=���>'��>?���������B���V����<�(O?����d��
�Y〾�s*�H�>^�9?gf�>���ڝ��H���L�>g�1�}5���ؽb�<�)�>�?0��<�55���Ҽ�QϾ[8/�u�;<��>��=�^5<,���+��gQƽv� ?	���aF	� �>�%U?�y�? �s?�Q�>X%�>T�'>\2?Χ�>�o�>]ȗ>�Bk>�@?-b�?=5C?�]�>�>Q0�\�Q�ܫ=�o��ݭ�*��bɽ���=���=)�z�|��� !�#���J��^~
=T����A��-�<��>ֲ:?�ȕ>��X>�e����I�>#O���=���>`Z>Y�?��>�Z?�3�>z�?�f0>�D����䢾"��>��>��v��&����=�.�>�?>��c?�O+?�)/���O=���>�>?�?lWS?Xe�>�;}�Zg����޿��<�ב�>q�NRS=�6�=qVf��=S�?���q����<y�>�G�>�qq> Z�>�QO>C#>F��>-1e=�A�=&4�=y�]c$=l�;�󂻄���&��y�v\�����B��;v���|�����J�UO�H��>�G?�ܣ�Y��=Fi���쾠2�lĔ>��2=�e>X��>�`̽�����n�4
D�;�]����>PNg?���>�|$�;>3;������=<M0�>ܘ�>%�6>��=���Mf�ñP>:�>��E?�5�>V����h��	���37���A>�[�"z��#�?��N? ��/v�������*��S�r^)��/��du��O&�%J��2��,7�;5�D�#�^[>���>$��?����!X=���-��q���PR��1�=4m�>��>}�	>'F񽱴��i(�����7Q��B����M?�>�>�y@?��?a?q�?��/?;)˽<?r�>�e�>���>��?�V?�>��>�Q�>�ۢ=O4ļ���o���˽N��ek	>, />�H>�>���=��->%�6>^����Қ���=]$�=,8>��=dy>�)t>*�*?T�:?�	Q=��[��2���j��'�>�b=���=7��={n���0�>�v�>,�,?�,?�G?�y����"�#�R�S�������03?`?$��>3�S=+�=V���yL�ó+;��B>f���������Ҿ�OU�q��>�^�>Nb>X9_>q({?�8C?2#?�,�/�-�M�u�
Q+�9]Ѽ8�;���>n��>�`�=߾�3��t��a�L0�� !��k?��=uq�=)W>�+>6�=�`>W�(=�p��<ҽE�<%};W�>1�>��
?p/^>e�=4R��� ��UI?X⠾���R����7Ͼ'V$� �>�&:>��U5?WW�*�}������=�xw�>�>�?��?��d?�B�I����[>�WU>��>��<�_>��`�7(x��/>�h�=viv�ᬕ�Z��;i[>_x>��ɽ�9ʾ��l*M�s츿��}�C�ᙦ��l�?-����l�k�d��i�~��@U�M8��������	�.���^�J����i�������?w�?��}>[������d.�N��d��o����DK�(�¾	&U���Ҿ����UվL�&�k�X�������j�>,�Y��&���|�$�(�s펼��>>k�.?�vƾ�������wd=��$>�B�<Q��O���䦚�w�
���W?��9?p�뾙5������>;?�%�>�$>����S�뽀,�>�3?ǜ-?ͦ�����+���i���h�?7��?��??��O�j�A�>�J���5?\�?��>�Ŋ���̾�`�?��9?���>�&�9g���3���>F�[?�8N��mb>U��>V:�>���g���w&�)@���l����9>��
�����Lh� 0>�K�=j�>h�x>�"]��	�����>K�c�N��wH�W����U��<�Z?Le��>��h>&�>��(����|ǉ�����L?���?o�S?�\8?�=��������<;�=6��>���>q��=ג�J-�>���>�\�^jr������?�<�?p��?�WZ?)sm�lɿ����4_پ�_����= SC=u->C{�ph�+z�=�bP�n>��>5:c>uw>� V>�F|=)��=����"�Z.��y����H�(-�����Z
�i�J�l�վs(�Pa����q�_���\ۢ�P�C�ܩ��R4��x�-�����>�6?���>��?��p>hs�<g��3��2��;����;��*.������1,��,˾�'ݾ����0��hX5>�ݸ�A��=X]�>A>>q%>L$�>�s�=!��>M7�>Ђ>�\�>J��>��>$J=ه>�C>���>��B>ூ��c����F����%*�<�79?*�8�����$�Jꬾ�m���Y>Y�?�d*>�^2�?ƙ�����ᔳ>�õ�]�`���w�wȑ�Iq�>q�>��=��7��<it����]f�=�Ü>j3D>K��==*ƽBs>���$<�?A��Yͼ�^�;��>�e�?k0Q?��>�r�>\|�>��?���>�^�>�g�>�՝>�/G?�;?�[�>�/�>�}&>��D�<�z<>��A���G�0B@<��-�N�;��<�Q=��Z��G�vp��Ƴ�=��=�l\=^��=:�	?b]N?o��>4��>YOh�G�z�n�Z�>$�<T��>�3���>8�
?/�>��>jV�>�=�ߩ�U��[���;9�>��Z>�~��猿}���T,�>�j�>	1?�c?/��=�����;Ś�>H��>³%?%??�T�>`Z�<,Dɾ���*K��>cf��Q�x7���>���[>�l�=G��H>�m������>���>%\�>z��>�?aW>�2>�R�>�_>(c>e���G�m���}B=�b�=t�7>��=�T0=|��=�0�Si��~��7�^���<-�="Rۺ+?'5?2�T>a�>�E=n����'��eY�$2�>�A?:�;����M�R��XR�J/m�)9߾0�>
΋?��=?u-��'L=$x���4��8>�>3J�>^G*>lƼ�n��>�\?Y+?ot�>_�E��s"�5�a�p."���@>4O>��:�dy�?^X�?����C^��5�$��]l��/��˾M���G���.��a��
B�s2��4�Y`V>F|�>%��>��?�N�=��>k篽�XJ�c��y�
�����.�@>q�M��1žR����뀾/#���%�����p>���>���>���>D��>��>��P?��\?pl3?��=x�?7��>��'?��>@1?}$?M?ܫ?ظ>�:�g���'����q�Y쮻���=�A�>���>&Re>��:�j)>��6;�B��,�7�d��c>(A�;���=�-H>.~�=jN>g=?�-?����S�4ㆽ�@-��o|=��&>B8<=�=��C=��v> g�>}��>�@?���>�U�<���6�(���𾫖��E�)?(�B?��?C�t>|aP=)��J���s>�¬>��=T��]㢾%��Hc=Ӵ>�C�>�x�>�I�>ss?R�]?o!4?��n=>�{2d��V����<���X.>e7>m�2�IV��UG�s��q~�������=�\��D=k6=X|*>�*�=p#S��1�=�v�>�D��׷���@d>���>���>�_>��
?��]>T���� �����I?����i�L頾oоY���>��<>� ��?]��)�}�?
��XG=�Љ�>X��?V��?�>d?��C�!���\>�VV>>>�.<��>���{���X�3>/�=e{y���3؝;+�\>e@y>m�ɽ;�ʾ0��fH�|�J���O�U~ʾE׾�����`�᤻L��
�.�����m��㌾����&�߽��e�	��	u�Q������?��?g�>ˊP>�ּ��Q!����5��\���m��U����=��4� �Ů�8gI��?H�Q�,��Yľ��>��Y�Q���Z|���'�L����F@>�M/?܎ľ9��N<�)o=$%>�0�<n��O��RL������XV?��9?N]�����ݽK[>�
?�-�>�[#>Հ��x?����>3
5?��-?��!C��`E���Ԉ��u�?���?��??JP���A�B��Bv�?�?@��>�9��6;���??W�9?���>��`H�������>�c[?�M���`>���>��>3��:��c!%�r���#�z�"�9>������_0h��>��.�=v7�>:Gx>�!\�񊮾��>բ��[&��P?�)疾6׏���T�k�9>�^�g�~�R���:�z�V�t������3���:b?W�?��i?'?ܚ��`��Ϙ�(�>���>��.>2Z��H��=���>���=�oJ���Y�����#�>���?��@�:�?����T�ؿ���L��ux��E=��:=��6>sC��M!�=�,�;�=��G�;�b=��>`F�>�_k>I�k>�UI>x>�݅�@�%�V졿�č�p-��u�06�$(��E���������_��S͇���&=�=:-5�`N)�?�̽��=�9�� +I<�r�=��>l{�>ܬ?e�>.��37��h;�	Ԅ�ǹ���"�����f����[���z��>ɾ��&=�l��!?I�F>dID;gZ�>h����L>x��>�l
=g_<�����5=
�>>��>���jL>FZd>C�=u/8>�%>j
�����=�V�>4`��|V'?�x��q��P�羾#��)�Z���\=-}�>+��=ȢT�@@��6̍�^��>��<.���l8��\�=4��>� ?�>G�`��8�>�
�'b�� �=��>t��>��_=�:\��b�=ի$�L�>�վÖ�=Mpx>B�'?��v?��6?[m�=���>b}b>U+�>'��=v&N>�S>��>:?7M8?�70?�>~@�=�k_��O=W8=�>��xX�-=���"ۼfZ�V,�<�F1��B=9�q=z�<9�d=ýD=U���ܙ�;��=�?�1@?�>2�c>ʥɾL==���k�h���\>�C; ��>��>�?�)�>�U>�Q1�;�s�M6뾂������>n��>1�y�D���e��\+�>�v >�V?�0V?!~7>�
0�L��=���>^Q�>�j?�::?�n>r@����pN��翊-�5���m��q��߈;R�"������ʽ���҂L�Fߵ<�̩>M�>���>�6s>�la>�� ?���>m^�>��W�<�z�<e�m<E�Q�☫�"���� <��M��r��W�3���2���M�C�(��x���@"<$?��?� �;t(�=���;*��ވ�ꢓ>�l
>Į>��1>�:#�t9Ҿ�o��}B��]e��Y�>��^?�?�14�a�=+� =���	>́�>[s>�>Q���н'K!���x=�ݡ>q�?Fm�>K���1�l�삁��/����>Pn>>� P���l?\#^?����徼#�9���R�V���Y���¾���@�ݾf�O�>o�8O� ���Py���/>�'�>X��?W���\>������߲��ᡜ�L�k��`>>v o���?�7b>U"W�D}���%�����D�����=��>�>^��>��Y?]�?E��>8[�>Ռ(?3~>""X?޶�>��2?"�4?�5?��B?^��>_�^=����[�<v1�=�ҽܱ��LO�<zFJ��g�=��h=L<>��->�A�<?%��%��x[(�y*(=$ғ��cG=$�=��8=R�<^��=��(?pM?Q1���;��^���Xڽ���Jj����&>X�>�ʜ;HPu>=r�>�?n!?EcV>�餽�nR�w>پ����=��K?�u?�	�>2����>�<9�G^�X�*�̑�>'�t>�׾�ڿ��ī��S���>���>��R>��p>O�?+f??��%?|��3,���o���/��$� �c<�X�>漫>��=C�ľ�&1�Y�n��5[�V�)���y���X��[�<�	!>�(>ہb>��= � >�?T=+JD��*�`�<ގ��{��>'�>PZ?�V>���=����nu���B?���aþeq�����>gþ��۾eӾG�D�p��!���������ani�E�>�6�?6��?��?R�߾�E��P��``'>8��>���鍾�x>�_t>z���B�n>����=�;�>(%>���>U@$�r�qC���v=����a�􅚾�'˾�Td����h�s�+�����f��>�IϾ�\�����S0
��d���;�j(�������N�����?�~?II�=l U�����Wq��0㾪r<溾z����Q�����;ξ3{��龎�� �B�N�#-�賞> N�<���E-~��*�%g�;�5>�9/?pžM��Wo�uXb=�*(>��<�m�y���|z����~�S?�H8?��M���K׽��>�y
?0��>��>�叾�%޽���>4�6?d�+?�˼	ԍ�Ɋ��4w����?a_�?�A?8�;��TC���	��N$��?��?�u�>n:���x���
���?�9?�[�>�E����N,��B�>��X?\�S��]>v�>���>���zė��3��.���&o���,>�{;=�콡Lm���1�5^�=���>ζ>�R�8��<[\>U���" �HWj�dd���q۽m_���_�<"�ھD�q�c'�������f�Iz�G���ɫ�=�Y?���?� X?��'?�6Ͼ�E!������>��>J��=�ϼ=kl��8�>�M>����=�6�پ��>�>�?���?���?�q����ҿ!����P\��R��K��=��B>ܹ�>Eԝ=�<�={�ʼǈ��VP�M�=ߑ�> �>�K>'�>,{�=�� >�y���Y��x���{�@�+��Y�J���+���-�_5����+�G)��^ξ�)�āB�a��m�O�g����s������!>�y ?���>9)�>�e�="&_>�䞾e�
���D���¾�M)�������;�M���� ��2�va�<̢���ͼ?�4;�E=�>�/�<��>�c�>|a >�>R!>&JF>�C>��=n�H>���=tr>>���=n�>�y�>4Ρ�m���wM�)�)=q�Q��Z?��=:%;�v���N�>ɽ�\�>���>�UQ>N�?�ː���ǀ�Cܧ>�����x�Ck�J������>Aء>\�<��
���=<V��Q�]�]c�=��>m �>t3>����_������C��>��־�T�=�w>Y�(?Y�v?|6?WK�=���>O5b>\>�>E��=Z�L>v�Q>W�>��?��9?#s1?V�>�Ӿ=�\`��O=�::=נ>�غW�U����⼎�&�g�<_d0�#cG=}>r=Jw<��`=��B=�fƼ�֧;6 =w�
?�B?|F>�Io>ӄ����C�P
��/���݈>��=�w�>lǷ>,�?��>��K>Z#
�f�g������Q�Ӗ�>rk�>����i��Q����h?������|?��b?���~��f�>�{2=H� ?!��>J�?&�X>���_l���Q
��"ѿ�:��+�|h2�YI�P�6<��q���x�z���A���H��O'<�&I>�ق>�<>r�>��=�X>"��>��K>i+�=j�>Zϼ������c��:��q��=9d�:(�ʻ��!=o׽�]h�O��bc��J��d����d�>ES�>~��켋>�n��P��k=�s�m9�TS�>�L>c����ʾ������[���AZ�>�=^?�'?�Ax���U>�E��'��˺�˖=���>!ȭ�>;�=ݺ2>�W�<��C>%�R?P$�>77����@����ޓ���>4a½G��aj�?j�>?.��2о	���O�xs+�<����j����1;�2�DsK�o�0�11�*������>�\?B��?����c�/���ܽ�rs�&���Bо�}l>��.��>�>�Ѿ��|�GK<��`���Kq�t��>_��>\/<>(��<� 5?pq!?	�>�&?�[�>)'�>�p>?�F�>�Z?[�D?/?�3?(�.?3�<>���<�(:��ѽ�F��Q����>�#���v>Ì�=*#>Ģ�=i~�=T�<���=�Z)�$�����J�h=�H�;p��=��>��8>g,*?�!?
c��1�?�8���!�����q�=w��>�9L>�P���=���>�)?~K4?]G�>Z9μ�I��3�1�rW�"�d?f�R?�P�>U��9�=�پT_��X&��?�>ؤ>�l�|���Y���u��] �>22�>�
_>&�f>gY~? �A?��"?���0�-Su��+��Ƽ���#�>�۞>�=��ݾݩ6�Ks��!`��W0���-��E��=��=۲>U�<>���=�>�U=�����ѽ�B<��X�>g��>��?б[>���=O���gp� �?M������c&��]��=Z"=SG��f�=���Z3�=� ����[�ya���S��ٗ=���?8��?��?�l��so��L�:�G�=��>�芾�<���>�'>Pԏ���2=���<'$��k��펳<?�Y���˾S����#=�6ȿ$k���=	�]��&��xE�6������M�۾�X'��"оX�����:'�Q ��G����觾*t������?>�c?Gd>ձ����6��[ ��T��£���{龪uѽY����mA�����X���{�[�{�I���V��e��>
6Y�7���|���(�/��ڨ?>B/?�Rƾ0������ܩf=�W%>��<SY���� ������sW?j�9?`�!S���e��>��?� �>�&>̽�����m?�>1L4?f�-?�5缈���)��ڧ���\�?���?,�??�cN�2�A���1����?%�?[^�>R����w̾����
?�9?��>���8O����`��>Jm[?��M���b>���>�.�>Y��G����f!��'����u�;>A�%����"�e�`�=���=v�>�#w>��]���<[\>U���" �HWj�dd���q۽m_���_�<"�ھD�q�c'�������f�Iz�G���ɫ�=�Y?���?� X?��'?�6Ͼ�E!������>��>J��=�ϼ=kl��8�>�M>����=�6�پ��>�>�?���?���?�q����ҿ!����P\��R��K��=��B>ܹ�>Eԝ=�<�={�ʼǈ��VP�M�=ߑ�> �>�K>'�>,{�=�� >�y���Y��x���{�@�+��Y�J���+���-�_5����+�G)��^ξ�)�āB�a��m�O�g����s������!>�y ?���>9)�>�e�="&_>�䞾e�
���D���¾�M)�������;�M���� ��2�va�<̢���ͼ?�4;�E=�>�/�<��>�c�>|a >�>R!>&JF>�C>��=n�H>���=tr>>���=n�>�y�>4Ρ�m���wM�)�)=q�Q��Z?��=:%;�v���N�>ɽ�\�>���>�UQ>N�?�ː���ǀ�Cܧ>�����x�Ck�J������>Aء>\�<��
���=<V��Q�]�]c�=��>m �>t3>����_������C��>��־�T�=�w>Y�(?Y�v?|6?WK�=���>O5b>\>�>E��=Z�L>v�Q>W�>��?��9?#s1?V�>�Ӿ=�\`��O=�::=נ>�غW�U����⼎�&�g�<_d0�#cG=}>r=Jw<��`=��B=�fƼ�֧;6 =w�
?�B?|F>�Io>ӄ����C�P
��/���݈>��=�w�>lǷ>,�?��>��K>Z#
�f�g������Q�Ӗ�>rk�>����i��Q����h?������|?��b?���~��f�>�{2=H� ?!��>J�?&�X>���_l���Q
��"ѿ�:��+�|h2�YI�P�6<��q���x�z���A���H��O'<�&I>�ق>�<>r�>��=�X>"��>��K>i+�=j�>Zϼ������c��:��q��=9d�:(�ʻ��!=o׽�]h�O��bc��J��d����d�>ES�>~��켋>�n��P��k=�s�m9�TS�>�L>c����ʾ������[���AZ�>�=^?�'?�Ax���U>�E��'��˺�˖=���>!ȭ�>;�=ݺ2>�W�<��C>%�R?P$�>77����@����ޓ���>4a½G��aj�?j�>?.��2о	���O�xs+�<����j����1;�2�DsK�o�0�11�*������>�\?B��?����c�/���ܽ�rs�&���Bо�}l>��.��>�>�Ѿ��|�GK<��`���Kq�t��>_��>\/<>(��<� 5?pq!?	�>�&?�[�>)'�>�p>?�F�>�Z?[�D?/?�3?(�.?3�<>���<�(:��ѽ�F��Q����>�#���v>Ì�=*#>Ģ�=i~�=T�<���=�Z)�$�����J�h=�H�;p��=��>��8>g,*?�!?
c��1�?�8���!�����q�=w��>�9L>�P���=���>�)?~K4?]G�>Z9μ�I��3�1�rW�"�d?f�R?�P�>U��9�=�پT_��X&��?�>ؤ>�l�|���Y���u��] �>22�>�
_>&�f>gY~? �A?��"?���0�-Su��+��Ƽ���#�>�۞>�=��ݾݩ6�Ks��!`��W0���-��E��=��=۲>U�<>���=�>�U=�����ѽ�B<��X�>g��>��?б[>���=O���gp� �?M������c&��]��=Z"=SG��f�=���Z3�=� ����[�ya���S��ٗ=���?8��?��?�l��so��L�:�G�=��>�芾�<���>�'>Pԏ���2=���<'$��k��펳<?�Y���˾S����#=�6ȿ$k���=	�]��&��xE�6������M�۾�X'��"оX�����:'�Q ��G����觾*t������?>�c?Gd>ձ����6��[ ��T��£���{龪uѽY����mA�����X���{�[�{�I���V��e��>
6Y�7���|���(�/��ڨ?>B/?�Rƾ0������ܩf=�W%>��<SY���� ������sW?j�9?`�!S���e��>��?� �>�&>̽�����m?�>1L4?f�-?�5缈���)��ڧ���\�?���?,�??�cN�2�A���1����?%�?[^�>R����w̾����
?�9?��>���8O����`��>Jm[?��M���b>���>�.�>Y��G����f!��'����u�;>A�%����"�e�`�=���=v�>�#w>��]���<[\>U���" �HWj�dd���q۽m_���_�<"�ھD�q�c'�������f�Iz�G���ɫ�=�Y?���?� X?��'?�6Ͼ�E!������>��>J��=�ϼ=kl��8�>�M>����=�6�پ��>�>�?���?���?�q����ҿ!����P\��R��K��=��B>ܹ�>Eԝ=�<�={�ʼǈ��VP�M�=ߑ�> �>�K>'�>,{�=�� >�y���Y��x���{�@�+��Y�J���+���-�_5����+�G)��^ξ�)�āB�a��m�O�g����s������!>�y ?���>9)�>�e�="&_>�䞾e�
���D���¾�M)�������;�M���� ��2�va�<̢���ͼ?�4;�E=�>�/�<��>�c�>|a >�>R!>&JF>�C>��=n�H>���=tr>>���=n�>�y�>4Ρ�m���wM�)�)=q�Q��Z?��=:%;�v���N�>ɽ�\�>���>�UQ>N�?�ː���ǀ�Cܧ>�����x�Ck�J������>Aء>\�<��
���=<V��Q�]�]c�=��>m �>t3>����_������C��>��־�T�=�w>Y�(?Y�v?|6?WK�=���>O5b>\>�>E��=Z�L>v�Q>W�>��?��9?#s1?V�>�Ӿ=�\`��O=�::=נ>�غW�U����⼎�&�g�<_d0�#cG=}>r=Jw<��`=��B=�fƼ�֧;6 =w�
?�B?|F>�Io>ӄ����C�P
��/���݈>��=�w�>lǷ>,�?��>��K>Z#
�f�g������Q�Ӗ�>rk�>����i��Q����h?������|?��b?���~��f�>�{2=H� ?!��>J�?&�X>���_l���Q
��"ѿ�:��+�|h2�YI�P�6<��q���x�z���A���H��O'<�&I>�ق>�<>r�>��=�X>"��>��K>i+�=j�>Zϼ������c��:��q��=9d�:(�ʻ��!=o׽�]h�O��bc��J��d����d�>ES�>~��켋>�n��P��k=�s�m9�TS�>�L>c����ʾ������[���AZ�>�=^?�'?�Ax���U>�E��'��˺�˖=���>!ȭ�>;�=ݺ2>�W�<��C>%�R?P$�>77����@����ޓ���>4a½G��aj�?j�>?.��2о	���O�xs+�<����j����1;�2�DsK�o�0�11�*������>�\?B��?����c�/���ܽ�rs�&���Bо�}l>��.��>�>�Ѿ��|�GK<��`���Kq�t��>_��>\/<>(��<� 5?pq!?	�>�&?�[�>)'�>�p>?�F�>�Z?[�D?/?�3?(�.?3�<>���<�(:��ѽ�F��Q����>�#���v>Ì�=*#>Ģ�=i~�=T�<���=�Z)�$�����J�h=�H�;p��=��>��8>g,*?�!?
c��1�?�8���!�����q�=w��>�9L>�P���=���>�)?~K4?]G�>Z9μ�I��3�1�rW�"�d?f�R?�P�>U��9�=�پT_��X&��?�>ؤ>�l�|���Y���u��] �>22�>�
_>&�f>gY~? �A?��"?���0�-Su��+��Ƽ���#�>�۞>�=��ݾݩ6�Ks��!`��W0���-��E��=��=۲>U�<>���=�>�U=�����ѽ�B<��X�>g��>��?б[>���=O���gp� �?M������c&��]��=Z"=SG��f�=���Z3�=� ����[�ya���S��ٗ=���?8��?��?�l��so��L�:�G�=��>�芾�<���>�'>Pԏ���2=���<'$��k��펳<?�Y���˾S����#=�6ȿ$k���=	�]��&��xE�6������M�۾�X'��"оX�����:'�Q ��G����觾*t������?>�c?Gd>ձ����6��[ ��T��£���{龪uѽY����mA�����X���{�[�{�I���V��e��>
6Y�7���|���(�/��ڨ?>B/?�Rƾ0������ܩf=�W%>��<SY���� ������sW?j�9?`�!S���e��>��?� �>�&>̽�����m?�>1L4?f�-?�5缈���)��ڧ���\�?���?,�??�cN�2�A���1����?%�?[^�>R����w̾����
?�9?��>���8O����`��>Jm[?��M���b>���>�.�>Y��G����f!��'����u�;>A�%����"�e�`�=���=v�>�#w>��]���V=�ᙾd����j������4�*/��I5�=���#�����8�&�Z�5Á�h3����=�q�E?�R�?V `?4?��������켫XH>��>�@�=0'$>������>�}�>����2T���*&?nY�?9��?�Wz?��r��r������ W�?쓾r�>�l�=�z>�����=QI�<P����m�;���=x�>v�v>o�>�2>i?>Gq1>|݀���x��\ː���@��Z(�^U� �����Xr��g���ľ`�Ӿ\q���P�cK��/��S�<�&j�=$����i==��>�g�>d:}>�3� ��>�'���u%�`I5�K-�"C1��~̾�9�+�������n�X�!����Ԯ<r��ܼ>h�<i�T=<��>�w���X�>f׫>:x=u�w>4b>�ؼ=���>�Y>l�=7�J>�>�a�<���>�x>�4��t�u�&�?��-F�39?�o^��ǽ�� �ᖾ��4��)�>�?�-�>���p����)�>�l�<�͍�H�	���u=b��>���>�Dt<��:[��m����$���$>���>��|>ū=\b��"�ᬦ��j�>*���=��r> *?D�t?F?9?�>��>Vau>Q^�>E�>0Wa>屆>��>^�?5�)?<;?���>���=ϔK��w�=�|2=�]�CQ����V����ك�������q�=�5i=V��ܡ�<f��<�f=�`�=�j=M�!?	�?m�>��>U��8�-��$7��>��l>�>�u?|^�>�H�>�5�>>��>�*�=\�񽐑��|Ӿ�)�>�?�<j�hA����<���>���;r?J�W?�%�=�=c~�>�Q">�j?�9?�6?�`�>o,�=`>������jӿ�
$���!�Ԃ�e����;O�<���M��5����-������{�<W�\>_�>��p>��D>��>J 3>�N�>�,G>��==�=t�;5�;��E��7M=�+���F<rQ����'8Ƽ�^��쿋���H�r�>�$U���ؼ.a�>��>�y&�2�u�t�(�4W᾿ �K�>R�u>ZX�>o�>�1�,�#�5�i�x�/��U���?^�?:��>Fi��-'=NT���c>���=}
>)%�>	5�j���ϮL��6=v��>�,?��g>K�&�(}X���|�Z�X�>"�u��|?�i{?c��r� ���(�0��2L��B�=�T���׾����D�"�@�n��N
����3�>:c�>�;�?
�T���>���gv��Z#�J�|�g�=J�>��>	x>&(^=~d����ࢷ�&"ƾM��ZF�>.�s��T�=W�?�N�>`@?C%?5�>�^>�/?\BG<+�?��?�Y?��?�D�>��>�O>m��඾������Ri><u=t�=��==�>�?�=Nb����$z��K�Ὀ��*�潸���^<׊k=��=��>��?�j;?������;��ڈ�vc>\cB=ag��.�>�R>���=��>��>��)?�K?�@?ԇ>AAξ���9��x\�".K?+�?w�?]Cj�ܵ�=��̾�㕾��͓>y�ϼc���Cȱ�����|<���%>�Ui>u�.>�,g>��~?UB?�9"?B��I�.�WAw�4`+�����{@�x�>��>���=��۾6�6�+;s���`�F�1�CB<���F�}>=�	�=�">��@>���=�e>"=�P��"�ؽ��:<b��e�>��>J;?+W\> ��=�e���7�	�@?菣����5Q��sD��> �~��=�+>q��Ķ�>� ����*j���KA��J�> ��?՘�?
m?��6������I>^�P>&�<>��ռ�YB�\ݼ���>���=��a�������c<39@>?/�>�C��`Ⱦ�RL�[9��8�7���0�����S*��H�۾�Pwн`���܃.��)�1WN��ċ�k��3�Y�� ���h���u�v`d?��m?]Z3=�����-��q����C�%�����s�f���۾{�P�;=��
�վ�������{4��� ��¾��>�)4�<@{��;|�wJ��v��>�<?T�þ��ƿ*�E�5<��j=�n���&�:��^�������h?�-?ԛؾ���g�D�i$;>��?�2�>�-�=�SW�{�&�S�N>jB?Z�?�[��]������@��<'d�?D�?T@?[�N��A�g����?��
?4��>�M��(˾�%�6{?��9?� �>�����e�\�>��Z?�\M�Z�h>g�>�-�>�Z�ђ�8�-�@��6Aa�&�<>�G߻jV�gYe���;�9q�=�h�>x>Ի]��������>�@꾮�N���H�������F�<5�?ǎ�V8>�i>�B>��(����ω��,���L?���?��S?�k8?�]������	��=���> Ӭ>���=���8�>���>Qe��wr����?qJ�?T��?�[Z?��m��Wҿ�&���۾�	��ם=�n�=M�p>(=(=�&�=�	��	g��M�=�_�>�N�>�S.>"7�>�U�>�8�>o+>�P��&g#��ՙ��Ƒ�cJE�!����%��f��۾������G�p��Ǌ��@��)D�~%ؽ�&�����I?���j����=�"?�n�>7S�>��
>�.�=������,���$��0����診��b���Xž𕨾�q��ھ1޾�>�=޾�i!?��2�Ac�=��>g�-�%Y�>�>ϖk>��><\�>����"�j>��D=xVm>C�<���>!�=/"�>�=C���[��l�9�:JX�C�ú IC?�PX�����_h3�/�ؾb���wc�>I�?�V>>	'�Ȕ��7y�-��>P�=�M�_�#�ѽ���0�>���>ɶ=�3� ��Z�y�������=�U�>��>)~p��슾����q�=B�>HuѾ���=�9���/Z?���?�n?��>���>��m=z�>N�-�PM�>���>]�>Q�>��#?#L>?�J�>	�>ig��C�� �ｘT���9�=ll�#��	��h����8�~7>&��;TFL�#=������2f�=f�=��?,�G?�)>�)�>[����7G�<`�k����>�[�%f�>��2?R�?���>�U�>�dL>y��qp
����H�>f"�>:*O��ց�n�C=d�>D��>�?��[?����X��M̽7޲>�?��+?��h?(4?��=���	R	�^�ڿI�&�	/I��2��ꎍ<3��=5l]=�E��^��'��	蔾e�=�C�>�5<>�Tn>p�>�Zi>/!�=:�>*K>�$�=.��=�ZY<V�����lL<ؤ�tF�=���9�R�]k��o���+�<}@��]�0=�j
��T?;�?��f�򁚽	�{�"���?��$�>V��>��>U��>��=���Z���E��_����>y�a?��?�4�;��=4�k��^_<95�>�	�>�1&>�7����7і���P;w�>lh?�j�>7����X�xRj�k^����>%�3>F	 �X.�?�E?�9�(e�+�I��4���`�薩>tQT>����C ��}5��xb�A�$��"S���.�`�+>�?*ӡ?�پo����K��m���A���i�߅s>'V�>�KO?.O5>��ݾg��5<3�������þ�V>�V,?tWv=9�q>��F?��/?'0V?�/?w�<?3n�=1H�>��Q�
i�>�2��B	?W$?�E?�ޞ>�W�>A#�>�I����v�ʾW\}�@��Խ<qp>��~>�|�=��7� �a>Re�=Lܽ`B�=�i�<��iR�6D8�f�<�!_>0?�N?:$-��p=��=e���!/��hXa;=C�>C/�>Eþ<g�=�dt>��?&d?��N?v�>�Jy�f�����ㅼ]�S?�B`?`R?*�=~�> .;#{���2ڽPM>�ۀ�*j;^�Ͼ9Y��ؽ��>��?l�>з?��v?�r>�C�>k=	�ϐ`���~��)8�c�2>R��>�a?(?~A˾�^Q�h�U�x���x���P��?�>�\�h 3;�^�=�H>�#�>7�-��e�=�͟>Ŝʽ0�Ӿi ��ب�>�V?���>��?eڰ>��q>ދ\��i1��I?����a�8Р��_о��� �>��<>�����?i�Y�}����?=����>��?���?�@d?4�C��3���\>S�V>1>KO/<�r>��n�r���t�3>��=�Sy�j�����;r]>�8y>-�ɽX�ʾ來�H�(���_N�%�Gɳ�̯�������[��R�1�⾤�8惾�j��2���c������:��"�v^W���ľ�����?Q�?�cx>Q�p>�m�����#e
���v������F�z��7A��.B�����>�Ծ579��(T���h�� �B��>Y��6��p�|�a�(��D����>>�.?=&ƾ-]��c���g=��$>�7�<���`�������͊�-�W?D�9?{%�tQ���5�z�>��?4��>�%>�˓���콛�>�94?�-?��a���-���	���_�?���?0�??�&N�4�A�o��BY���?IF?��>�����˾w��&'?9?zz�>>��B���3�k��>�=[?fgM�b�a>�6�>�,�>8����p'��1������j7>_�E����g�C3=���=47�>j+x>� \�������?O>z�gxR�=�U��u$�����_�a�*�?��վ'z>�W�>c�
��#`��Ꮏ���~��R�/?#��?K-j?(�?�w�Z�����ő�=,�>�1?"f>��&={�>`�?!��,p��!�~�
?@V�?sr�?��J?�M��gҿ����ܒ�1Ӿ���=��N>�L[>�����R<����O=5̻=8�>ws>�"�>ja�>A>Q�->� >�"��� ��� ����.G�_r���	���i�=��f��y��!W��D���B�d�~���T��gl>���ɽ��	����6��={�F?��>��>���>>�>��=��ʾ��(���d|0�=Eؾ?i�%l�������y0���q�>�=7f��>��.=p��c	?�Xq���:>�N�>Yd̽��S>U��<e޽����=Ί5>t��<�i>r�>��=/t�>��>S��׍� �;���e��&E�^�?�*p�N�����%�8X���g�#R�>$� ?�S~>��E�io��$����f�>{ص=�$���K�s�=�v�>��>���<�Rd=��	���ӾD�A���
>$��>�!�>�L�>d50��/�������>dӾzz�=��y>�H*?�)u?�86?j�=c�>��a>i$�>Cɯ=�OT>��R>�>�h?�9?,�-?�S�>a��=Kd�a��<�1*=�9��J�M!��nԼ��1�tϑ<|�U�-=�t=��<��@=�-=� ؼOg��%=��?1�,?��q>���>�`����F��lT�$�Z��=�֣<�>> ?�k�>���>���>a��=�K��ݾ���>I�T>�K����|l��1߭>0�:>��+?��?ى�@���ơ@=RLX>��?؅(?b�^?}H�>6�y�]���=;	���ؿ�9�x���E�Y3o<�i<��?����]D*=�<�X�{�kH�='�k>6�>W�>>�@>�.%>��@>�=�>�&>S��=>(A>���<��!�@�/�u����˽~P�=�HI��(�O<u<'������^��H_���ƫ�v3��98?@?����oN��DƾXq*�����9?���>�&�>��8?�յ>)�3�9D���W�Gv־�8?*Rj?�=?ؽ
f﻽T����=���>1�9>bL�p0���\��8�������?�G?���>��=N�V�z쁿�*2��6r>3�=ɔ�>��?��d?R�U���l�L�@�j�O�$�3�7��TF�ƛ��S������OK��t�@cM�����0>�[+?=`�?��վ���oϾ�ߵ�Ջ��\�]��CԽ�=�N	?���>fj��Hܮ���K���� ,;��(>[��>�˽j�5>ͫ?5�>�k?�ޮ>B�'?�d��e�>'E�=��>�hL�W�8?�J�>�.,?�&�>V]�>�i��f�ǽȯ�5l���&@��P<��R�;L>m�=#B�=���]��=�)>z���Ï�ʃ���p���#=(�0=w�j>��?�g?� ����2��h�=�6a�S�Ƚ,���>��=����ȿ�=��G>�}=?��S?�d??W�=�.��K�%�	���
>��E?O�v?m�?+i�S�>�¾G)�"��=kx>���a�½6b�΢�}���w�>}��>�+1>�s>!r|?i"<?u?�����1�K~w�*(�S�{��������>��>�S�=޾67��2v���a�6�/�*��r.B����<M��=��>�1>��=�a>	�<팶���νN�<ҕ�c�>;��>L�
?�#l>�8b=�L��Y�	���I?�`��=z�Y���о!���>�R=>�����?:�k�}�'��~S=�3�>�m�?x��?�`d?�rC����\>�V>5I>{//<ܢ>�j��!����3>5��=��x�{��� �;��\>Q�y>l�Ƚ��ʾ#7�H����_�~����<O���f� X�k����Y��}��2<;=ǝ*��\M�'����m񽯾0�2J��"�*�þ�R��M��?�||?�o�>��>X��[�HG��|��<����QJ�:㾂�]�x������9���u ���?�'�_U���>�R��Z��M�y��+��F���=j.?�=о8"��ɉ��2=���=0�t� �����&ɜ��Ƚ�u\?��8?��о���R��7@>��?	�>�45> A~�w���f|�>��.?�,?K�4��N�������=г�?���?�}F? ];�4J�[q��>��k�>yI�>���>��r�=s���!�?�(?���>��	��*��P�$�;b�>��\?7�8�d�L>�r�>�ov>�&)��l��>f�pȫ�󥜽 B>Y��75����x��y>���>�9>�_�������>C1پ�QI���I�Y�/�4�̾�~6��I??�D��{u>Kd�>>��O��Q������^I�_>?!C�?��u?)>%?�᪾@f����*�=A6�=�?�Jb>k|���A=��>��ž}�p��(!�!��>�9�?2��?y�0?�=F��ȿ
 �<0���T��K�=D�>}v�>��΄���I����<�<�_U>cJ�>�݁>�)�>��Y>�U(>�=n>m�{�"��m������m�_�a@������2U�C�
�
�9���ɾ�|��sx��6�0��?�D�����S�z'?��Ř�����RZ>O|?:��>�i>7_&>�K>$\s�ӝ���;���ľ�n#�4U���rо=a�����p��Lx�����"^�= ��M�>��=υ#>4 ?�~S���>�K:>�t>�J>oG@>�N>�`/>i�.=y}>Mf�=�07>xݱ=Kً>��=�����,���0���?��r-��M6?�2�M���A0��q��YR�����>�Q?N�>�/�N���f�~�qk�>ya+��W��$���Kr>0�>y��= �=-���j-����}�=�u�>��@>�%4=��^����@��<�I�>־���=�7x>A�(?�w?�s6?���='��>@Wa>~�>��=��M>>�Q>*�>a�?j�9?�M1?���>���=,*a�aj=E�8=#�?���U��ﲽb��"^-�1��<(�+�HFE=>Pt=CT<t�^=�@@=c˼���;z =�4?��)?ϚF>LHr>+�2�����lU�@�2hZ>%؝�tI�>�^	?�� ?\�?�H�>�N>N���3����P�>�S�>B��Mw�Pe�=��>M�*>�?��$?�������Lޑ>�+1>�?k2?��Y?��>� ��NȾ"��mӿ�$�;�!���P�t�;��<���M��С76�-�����.��<�\>N�>~�p>�E>��>�<3>�R�>�HG>�ф=S�=�;�;ܕ;_�E��M=H
��FG<e�P�_���P$Ƽ򟗽����I���>�#:��8ټM;,?���>���L���|���� ��⾣��>a�V>��?m�?،��DUF�V�t��ML�e���ә>��S?��5?0&�S�=>�:�.�=���>�Ӳ>��2�W�~�>|Y��/��㳾>��-?�&?C����B�zH��j/��|>�Y�=hľz]�?�B?Ψ'��ս��N����A�7�2y>��,<HS4�����s����<�r���%'�е��zP	>�?�j�?}ۿ�;�W���Q��Ͱw�Z�j��,>1DC>u?���=?r�p>ݾ)
M��߾��S�6D�>��?_�K�#3�>H?�HN?�|�?�;?� F?��R�m1#?�?��w.@=%��=[�C?
�?��3?Nԥ>k/�>�����.�(��}���`*>i2�bf�=�jz>oO<>zo�=�g�J^�=���==���XR��)����X�t�^���o�Ê8�&��>�B�> �U?vё����n>t�,�;X��'�p�f?J�3�U�9\�>��>�P*?CK0?$�:?���=�h��+D �,N����=� 6?"�m?���>��ʽ䃠>	��!J���h<��=(!ɾ�Q��<�澎���E�-�T��><�>zt>�t>މz?�u;?�? 
���-�i	w��f(������i;ᔹ>���>0S�=ڑܾ��8��js�4�b��o0�Z����A�y�=i��=4�
>�t?>`��=�y>�vc<1pu�<}��jR�;�<,e�>n8�>��?|cv>��^=����3��\N?���7��2Ŭ�W�9�	�>�/�>Di)�kM�>��ϼ+�y�|����P�PB�>�?��?AOq?��.��AJ[>�04>�2>�ɘ=����墽!��Y4N>'8�=
H����� ����?>��>�u�Ihľ�Eؾw������s�J�Z'J=�������T���䆆���<�@Dľ}�s������8���(�5��{�b�}��5ɾ�j���r�?0h�?-�f>۴�=�UF��N��v����">�4վ��8<��u�y%o��ׂ�;Z���V������i��k��>u?[�7����0|�f�)����r�8>�D/?�AǾQ��N1���]=�!>2��<����΋��Ě����ͺW?�9?��#��c��D�>�@	?Wd�>�Y*>㳐����>Lu2?�Y+?� �x���؋�p�g��i�?�'�?�A?6�M�;bC��8��S��|�>�?�?�>������
짽�K?�
1?bm�>�	��ͅ��� �c��>_U\? hD��f>�o�>�(�>�p꽒҂�m>�����Nz<�>�q��s׽�-��+	�Cǹ=�*�>P4]>�dz�����_��>%&�]�N�
�H�������힏<��?ۇ�6>		i>�^>�(�&��ZΉ�Yj�8�L?H��?n�S? o8?�w��L�O��,7�=^��>���>N��=e���>$��>Qk�*er�:�#�?�C�?���?<CZ?@�m�:�ʿo���Y���+1)>���=�nJ>�ӽw��=�"=�H@��kZ<R�
>f�>F`a>=e>.�p>�l9> f>Y$��X%������׎�-�E�v����
�;�i��v��������Բ�!���ky���J�vO����2�+���Ւ�������>�;8?vW�>��9>~*b>��Z>>�<���bR�\V �����%�Ѿ+V
�T��p|ξ��T�-���d5�z��=�}�5��>mEB=,���:?��a=�0>g}�>�
�=R��>2�w>���=6��=��Q>�?�=�>�t>wL�=K��>g\u>�J��s�b�,�/���Pm���z?[Rn�,� �	�S��b@�М�u�>��>���>��:������p����>��=�y�	�������`_�>�l>�9G>"��>�%�+'d�Z+
�g (>�?=�=k�>�������=��&=-4�>��龳��=�S���7?7ρ?�GH?�m&>�e�>� >�խ>�}�<i̟>�/�>�.�>9��>3�?`E>?rW?���=v8O�����&�������v�j�=t��<U�� �<�_�8~A;*�ٽD!��ή=����H����α� *?��E?U�r=w��>�ʕ���l�3_��P�t�����>y�>�9!?ur�>��2>�>O�ż�e��ZZ�St��̓�>���=5M��Q�Rtv>V>~�>��?R�(?.?�����Z%c�KR�> �?��>ثl?��#?}�ۼ0�����ӿL��^�Ж�d��=�S�=&�s�a?� )���Ͼ�m�B�Խ���<��>�9v>��>���>�Ґ>���>�v>��=X90=�> �������0������W���#�	=�
=��ͽ2�L��������ࡻ��=��?��? z�e��(��U���þ��>:��>�]?�A?�<->S� ��b���E�zf�l�>p�W?dN?��8����=)���PQǼ�]�>�.�>mb>"y��W���~��4�H=�>�>�y?R-�>F;�P2b���l��W��ϴ>�2j>� �rf�?�u�?D�w�(���=H�p_�8�?�tJ�>�B�(�ɼ}����;�)䂿���}=�0g�Af=�(?=�?_ ���@ :�ӷ�<^�������(�'&��1P�>mG-?�I�>%����1���Z���a��~�e��>�Q<��2<d!?�>l�K?�=,?��3?�[��s`�>Q��;nM?1��=�P/?� 1?���>���=$��>2��=��=�5��u�������l����<f5>Ĝ�=�#�<�^<�!<2G��<׼�Ʃ<e�B=R��ԧ���8�=y�=	N/>�{?�[?i������=z�=�o����M���2>F�#?���=�L�o��q�= 8�>�jF?v�K?��>�ע�F�9��?�5=7�`?)P?�|�>���=#�>�k��pm�7�=~��>t)�C�N��˾i臽����{�>��>��=NϷ>��~?�
?�?�r����S���{���p��9:��>9o?�V'?[���_5��{7�����;k��r8�j�T>��:��J�=|^��?�=�ck>��!<y�>Lñ=8���OT������<�W?}Y�>bM@?�0�=W$>�������_L?MIh��
.�΀���lx���7�^Gʼ>�X>�?����x��;����1��S�>���?���?�`?pb���}b���>$��>��>��=-et�q��=��
�(�<���\����������[<9�>����&����.��`q8=���O9�����ĉ������X��%���ԋ��㟾3Y�����$��zLG��S-���n�t��TA��Xzs���_�D��?ay�?w�>�j^>��(�c�z龯�>>�銾��F@��ݵJ�i�o��������S��;'2�rCE��o���>A�X�f2��;�|��)��z��K>>\�.?�ƾ�ӳ�Y�_�m=�">�c�<���5����њ�?���W?��9?a��ى�����;�>�?(��>�%><򓾭-��p�>8a4?�|-?���ʎ�_B��혼�P�?���?]e??ixQ�cA��~�$7�o�?��?��>�M̾8��϶
?��9?�M�>o�����a��	��>E�[?\RM�l�a>���>�Ɩ>�H�а���"��ݒ��
����8>޷	����(i�E�?��¨=���>Nx>�]��z��lN?^ڮ�,�`�ݢN�;'��aܾ�(���&?��������>N�>��d��a������s���+?+U�?��w?��?��޾[��7C��|�=�#�>>^�>��=¤>*�a>#�?(���A�}��U���X?.�?o��?�B?�(�n�ʿ�哿wI��V�Ծ�A>��U>{q>�D�w�:��=N�e=o1�<+&>�Ϙ>��>�a>@�G>�H>e�=>_�����!�@9��5����kE�0{��	�������_wz�#��:���󿾹��࠮���Ž?�8����r�D���Ⱦ�t>�1?�d�>���>��>�(�>�1� Qʾ3ȼ��޾[�־펾��ž4{��֟�.Jy�t"8�SR_�'�%=�|�
��>��8=`P���!�>n�N�K��>���>*P����G<8�~>������>v���w�=��=�|�>�q>���>��>���a����6�m�*��S��4?�n*>�k�(��Ǣ�"kq���>+s�>�/w>�42�a��ߓ���ѕ>La�;!�P���A��:-��G�>�o�>H�L<���=�M�� ��%��\�>���>v��>�V>�j��Η|�-jH��_�>�h��� >#S�>;B0?{f?�u4?��=]x�>Pp�=�)w>�0>�y}>�#�>(ځ>|A?�y5?8�)?#��>8��=b^����'�D��=:9R��厽�3�<�&�{�<Mv�</�,�1��<I"g=��"<�<��<boI<s���9=�X?z�4?�b�>G��>G{O�jC6�ҟK�y����!>"��<���>y>�>�?ޡ�>�O�>Ϯ)>������Ҿ��ཱྀշ>[�H>��U�ghz���D�3��>4ih>sE<?��-?{�9�$ܟ�HR � �!>=��>%�?�l9?.d�>U��=��U��l���ܿԇ��˾�)U���G>�>?��������\>�5F� �C��<+>hy<>N�a>!|>sP>T19<��=.?$%�=�3E>&}>�("���}ĽJ�`=�`�<��=.��=�M�>�<~��U�	�����%�c�n��=�V=��2?,�>�������N��\���m���K?c��>���=m�B?��>�"J���o�ƴJ�7��sL�>wpY?U<?0*#���=R
�<�ś<x	�>��>�E>����I�������}��>�@8?��>h�6��@��tr�@�(��Y�=�-�=�5��Ȗ?ˀf?m�@���d���2��U*���/�!��=lt��1K3=繮�'��*F���"��i?��$����=�,?"�?/m��}�<%�پ|���M��1`�����y��=�S?�X=R����\��G=��e������"�<�}�>Ż���#�>��2?�N?/�x?�/?�;G?\���x_�>��<R�z>®5�R4?�&#?w=?T&�>���>���I;�`�g���߾�π<03����=?jj>�p�>�SE>�Tͽ��>oZ>f�m�/�a�.�/=��#�I9"�,�ü��j<<��=�
?�H?8�Y��ޔ��WP=~G��� ��ٝ��	?��l>��-��5���>�'?��J?NcC?T��>Κ��ʢ-��!��>��)?�<S?õ?��3=���>�Y����A�ν���=6E���
�T�׾����2T�)��>��>s/�>�j>p�}?��@?]� ?�����`.���v�o
*��3��C;�N�>Ir�>:��=�A۾�6��r��>a�b1�{�4�<�E��/=���=�R>Vb;>Ue�=�>5;= ���t�ѽ]:4Y���ų>a�>}B?�+a>�&=����+��I?.1��mr�!���Rо�t!�&>)�<>����?n����}����q"=�~��>u��? ��?�9d?��C����&�\>~�V>r�>s8<�>�I�#J��3>/{�=Y�y�Aϕ�uY�;�\>4�y>�qɽ�ʾ��㾙�E�欯��kA��f�� ���as�3�y�̨����♾�"�(�
��3�U�ʽ�>���ޞ��s.���p�3ķ��%��f��?���?�Z>&ཆ�(����!�VUw�Hꁾ�1������G��\��&⾄)��R7	���7�6�7�z%�Lq�>¾E�A�����p��1���=��5?��׾�Z���j�ҟ4=|�=7Ƣ�����
��{H���K��Ν\?��6?�(ξ���$�N� �8>���>�E�>��w>��P���)�Ow�>��?ki?m���*G��.݅��e=O�?��?.rC?��>�<�C��M	�+�#��*�>��?���>�����������+�?��0?_ܮ>��	�W��* ���>��Y?kwI�ťb>X`�>�~>��?~u�b��C���Hg�F�S>�i��sB��*%��뽠��=+"�>�dW>О���NϾ'%�>aѥ�;[��������������&?٨����.\>P��=@�8�S뎿�_�2 �=��X?�>�?՛H?�~??9��h�*R���Vؽ#��>�d�>*&�>����G�>?�޾�g�m�+Cھ
�?��?��?�у?/
{��տ�ٟ��o��`Ҿ���>.H�>5,?�vt���q���=x5���6�^z�>���>��>��]>��>��=���=�����������M�I�Wd�����ou���r&�%���L&����\�þ�C	��md��g����<�MG���a�s���`g޽D~I?�S?�?>`]�>j�f�M5�>0�jT��K�t�6�=�]d+�<��dk�@�T�������b��n��=�W���>`W>Z;�>��$?_�F=?�>xH�>��<�D}>��p>=�1i>�<�>��>Ã�>O�>���=�{>�و=q'��$����:���Q�5�;g�C?C]�9*��y�3��b߾e���̴�>�M?o&S>U�'�����x���>8�E��Fc�p�̽�����>���>�M�=�����)�9x��b�++�=���>\�
>S�b�O폾���r��=��>���(Yw>0��>��%?�E�?�.?l=Y/�>T�2>G�>��5=�>C�>��>��?�I*?"8?%�>�!>��^�2������=d�W�����c��l�÷��34輩���-�=��t= ���4��`cV:,��,:=Z�Ƽg��>��9?k4�>��>C�^KL�VX�h���W�?>r\ֽ�I�>�§>P(�>x��>!s�>��.>pȽ.Y������u��>}2>��q�B1p��F�m�>�+>3vc?FD?ҽ�=���='>�>�>��?6�8?m·>IF�>��9�����mӿ�$�:�!�tւ���Zq�;�<��UN��!δ��-�����IG�<��\>?�>�p>�E>��>
#3>�Q�>�XG>���=��=�e�;�	;esF��?M=.���F<ҬP��Z�� qƼ`ė��L��0�I���>��|�Z�ټ~0?�?�e-���^�ꦼ�B���v���?]Q?�?q��>���=���GH��
E��Q�ͪ>��f?W�?�@e��&�>`�>T��c?�>)b>� �>�I��'s��]q7�L�>zL�>"o?�g�>D�&��Ne���� ���f�>��=;\��I�?AD�?�M ����W{���]��\&��a�<<d�z���jⱾ�*���0K��R<�Ժ�W<������	?N��?	���B�뾉���d�}�a�Խ��>��`>�Ѧ>Nɹ<�q���9��7����zK���k�=ݬ?� ��Mn>���>R�=��\?���>�0?L���t��>�8:>���>˒�>K�?���>T2.?1�>�}r>�e<�3轖7��缾�XT�!.p<��(>��>�Չ>q����X�=9e�=S�轼y\���=���=�tr=K�>�K�=֣l�64�=�?��<?�Nx�q���cʼVN��o=�Hc>�>�ߤ�T(<�p>B3>|��>�[?�O�>�k=��}�����	�@K-=���>�*?uC?|=�TI=J辑�u��N��U��=e<:׶��U��.��$��y.l>��x>������z>?]�?��=?qk?���~1���l��6�݋ἵ"�;8�>��>�B�=,ž��2�۴p��[�6�&�M#��U��/=� �=�/>}�G>K��=_�
>C�<`�ܽ����;��'�i0�>���>��?QvP>!��=$F��w���8b?��9���2�����ۮ�<섾`m���+�>�B=Xj�=2���G�,�xT���]�c/�>�d�??��?��?����˪���>FH�>E/3=���q轺�]��'\=6�L>P��=Q4����c'��7>�ML=���<�K��r�����d<��ɿ�)`�w������������bm���H����۾E)��k2	��� =���5_���ꆾ(��4?��vƋ?�9�?bt?j�>��=�;�&�Ueg��ߊ�ɞ���t���2��ф���X�uC��]a]�ۈ�}�P�~A��p�}3�>�B��H���9y�lI��_y�E��A�C?�����QU�i��T>V�=T��?�5��M���џ�,�����?�#0??���T�����*>�Q#?��>�s�>����h)��?2�__?��I?�h�F+x�}�b�g�u{�?�۳?��O?L�>|S^��2����&�f>���>��>��=a.H�6�Ǿ�3 ?��>8��=�(2��ꇿ��'�?\�?�R��{\>T%�>�y�>4�~��ƻ�c�$>bp
��ޤ��\5�
`�=����һ����8D>�d>��>���������>������F��Y2���-Ua����I�>&��}�P>�>����BV��]��y~���Y׽�%M?nؤ?��d?�8?��^���%�'ž�!>6��>k��>���>}��=�V�>���>{�Ծu[<��ܾ9�?֐�?��?��x?�N��ҿ�֙�����#���h$>gF>�ߨ>?L���o=�~;�X+����ܗn>?�>U�>�)�>ڎ�>��D>�-Q>4�������ϕ��3��E�Z��K%���-������#�r�6��'���
|��-9�L˽U����x�J��𽰗��.��1`>?��$?H�꽸�?;��>F7����ZI��a��$hs�硤<0H��x�'��Շ���+��= ����=* 4��
?��2>��> )?-�7>��P>�q�>+��=%��=w����摽	�><�T>_&�>(%>�<O>�i>�a�>���=�����ҁ�Q�6�h�[��x�uwD?��b�=���hG,���Ǿ�9��5z�>�6?��c>i�-��Г�4�y����>yI;�?;V�4ԩ�"���+�>7�>c��=0�ż$��������!����=
A�>C<7>,߽;�D��v� ��N�<��>��ھ�R	>T�>�3+?:�v?c47?#}�=�i�>$�[>BX�>'��=��=>-�a>Yo�>%_?fm0?�Y*?�m�>�Z�=��Z���>=���<2�T��B�#3����*��{��/U<D���[�<ͮ�<�,�3@8<�U�<�`���Jh�qb�<Of?��:?���>h�F>�<�w�8�>�<�V�7<cr
>��>�@?b�?K��>`�?�/�>�%�=�[��l���㲾%��>��:>��9���t�o���M>R[=a"K?ֹ?�������P�<��^>BZ�>�a7?�YQ?ڐe>��.=���>��%mӿ6$���!�I킽t2�z��;��<��M����6-�-��������<�\>��>��p>�	E>��>';3>}K�>�EG>Մ=��=%��;-�;�'F�t]M=�>�t\G<��P��c��O�żl���%���I�t�>��b���ټ�9?[6*?�f�Ҧ���d�<�M�<+C�r�?)1?�n�>���>F݆���G���44J�T��=Kf4?�%~?�B?�飽c�K<BE�<�x�=s]>�~)>:��>�X	�����W���e=� ?[�?�z�>�.�;T�%��E�����:>ɜ�<�����*�?���?/8,�G�ݽ,m���Y���⾧�ӽ����3��
�Ӿ��r�R���#�JG��F�m�>�)?.��?��#���\�!N������Ԡ������;��=�P>��>b8[�~���̾\rF��׾�A�ֹo>,*?�ɰ���>0s?N}�>��x?�"�>[�#?��,����>�=B?�-I>�)�>k��>�
?�멺�z1>���=&���%�5v����=��ٽ�pl��O>��7>������=-&�;?|ݼ`�����< ��\���Kͽտ�=͏���`>��?[y4?X��	�4[�>.�پ�R�dm�>;4㼇Ц�YYٻ�9_>�{>�j$?�z?�?В��%��p*�`W����<$�?K=6?�)?�|Z=n�q>���c2�½*=�> �f�jJžDQоR��8C��{:�>O��>�DX><�n>�L~?$�??S?@���ͣ.��t���'��N���q��Is�> �>��=��վ�-5�@=r��a�}U0�8'4�U�D���<z��=�]>�{<>�Ĵ=�5>��,=)���t�ܽp\<2�i�q�>���>܀?Ƚi>�Tg=⻬��R���L?��n�5�������>ľeJ���=�y�>���;�A?�ŝ�<��u����C�U&�>�w�?�;�?�Uo?�[���߽gYM>��>_s�=]l�<
r���<X�ü�xa>�x>_E��OZ�+X�=��)>�)�>�J����?���]�g��	ÿ�qX�H�=�@���gپf���}���۾1����׽�����j�>f=�=�
T:�xs���9�(/��и羻G�?$9�?I5�>59>c�V�-D
���6B��$�ھTcD��ܑ�ߔs��g��&����Ҿ$(
��,G���>�ӷ� Л>CY��=��i�|��(��5����?>�(/?[ƾ�ش�d��N�g=[%>l�<�K�Ӳ��E���u��fW?��9?�J��������cU>��?vj�>�&>���
�Em�>�J4?H�-?F��	��I7������_�?���?C?��!�֧>���������>�?vy�>Ѓ������2�Sm?�N5?N+�>Cy�߽���?"�*��>�DV?�Y?�.UQ>�R�>�/q>���kx��hϽG�q�""��f9>���9�ͽ0��շ�H�'>��>�L2>�?v��WϾ<F�>M/��|�>�A�����)Z��訾�`�>Қ���UF>��<�у</D��Q���"���b��IE?��?L4j? �I?���!G�ˤ��N;>X�>U�x>]��>��,>�ι>
��>����[��/׾~?��?���?�E�?ym�oFӿ�	��ϴ�����Z��=�#�=��>>��޽�˭=ќK=�I���<=�֊>B��>wo>`8x>_�T>Ǜ<>M�.>褄���#��ɤ��ؒ�3\B�!����vg��y	�zy�>���ɴ��񽾛���⥷�@ߓ�/�G�����R>����4L��B?F�?�#`>���>n�J=��g�(��/���^�������P�	���=�\�������V�!�Cd>J���?�==��>���>lc޼����툑>� �@RQ>�h�>�)Y>� O><�.�CT#>c&�=�q>>��/9V�{>.�=�!����e:���Q����;��C?+�]��]��#�3�S߾�N���j�>͘?crS>(�'�������x���>��F�f>b�Nzʽ,1�P�>b��>~P�=�λC)��w����Z;�=���>_�>��d��ُ�)�~��=��>`[Ҿ���=X�i>��*?�<v?�)7?�[�=�2�>�d>C��>���=6�P>ʩR>'9�>��?t�6?��/?���>4g�=�:i�A�<�8=K8<�*!*������H�N-+�'g{<P�5��mp=�|�=Q�<�a_=��=~ɼ3��;9�=�A�>�08?�r�>�S�>�)?�e�>�i&O�%=��->�r�w��>M��>u?v��>��>��3>�Z�.�¾U�ݾ���>�1G>�a�y��$��<cw>��j>�)Q?�2?�b�!�f�ĩ�<��=ԥ�>�s?�"+?iL�>Y'>�Q�����`ӿy#�y� ��z���r�����;�_B���b��s��O93��������<'\>���>z�r>?�E>�Q>�X2>o��>�^G>t�=�.�=@1d;re	;�$Y�y�H=�U��$<D=_�����mԼ�6�����hL��9���7�м�)?D�?����5���N�c��N־��>+�?�@�>�t�>����#��T�7U:�i�I�\��>od?��?�}�/�;>�os�^���^���>F�>�*���̾���<KЅ>r�?��Z?B��>{қ���t�%q���.N���>���{�Ծ�t�?���?�*����f�.l�&�ݾ�gԻ �8�P`ӽ���� �K��w'����@��#��=@"?K7�?8^��<��l���9��^ h��xM���O>�[>?K>X��,���'�Y,��x��.#<�[x>�B?h�E���? �?4�">h�?	S�>	L?<Ym=/�>�\T>!<#?�
�>�:�>���>��"?�Q�<�;�aZ�<�p�;�P־�t�� \�H��t��
�w>���=j ɽ�L>���=���N��H�=8�"���<=��|���>�=R?_>LL�>�L?u����$� j[>'ž6a>���>o��mO���>X�>#�>"�O?��C?�p�>�r�[Tоȡ��M=��{�:�
?��N?A�*?�s>\Ә>B�ݾ��c��F�n�>�R�(���������{=�=�>�^�>C�<��k>lG?��??�?o����/�.�u�k)���ʼ�^�=��>��>Ƴ�=ևоn�4���r��Jb��:2�++���M���=���=Zk!>v�D>J�=~�>@�&=�ǡ�g�ٽqU@<5S�����>���>G�?ފf>뫌=ꔩ�W��pb?��$�Pb�w󻾒����֦�S\!�,9 ?�m�>
�?�z���y��W_����K�S�����?4
�?�Њ?Ή���U��=
=��=&�>d�C>����">�����W��w���W+�J���k�_��"">�M�>�;?�)�^;)��8�4�п����=OX���_�����=�ޖ�/���U�Gݾd�F��k��y>z���T�D>�eu��~9��d��D���ؤ�?PB?��> I>A��DH;�,3��>K̑�A���0y�<YQ�������
UR��������8�<������>�zY�*@��`�|�e�(������?>H3/?8\ƾǴ�ӗ��g=�l%>�̱<�<ﾑ���������gW?��9?8I��&��R3ὠ�>j�?�l�>�%>�3��_[� �>"=4?��-?d(뼪���8��9����g�?���?�C?3�=)�>�5�F� �&��B�>9��>D��>�����ڳ���4=��1?BE?�R
?&��l����J�{2o>'�m?����X��>2�?^#�>w$�<�-Ծ������L����+y�<o$�&כ�Y����"N>�f�>��>2��=�d��G��>�4��?\�xm�n���If/���K��?��|�Ĵ�=^~">� �<�+�q4��?p���'� �M?��?:bQ?�?�K�����>l��=`f�=ri�>��>cR�_�z>7�A?�f>��F^�ԥ��F!? 1�?�`�?��5?��L���ο�������թ�����>}Ě>Y�g>&�w����<���=Է�̗J�k:�=�~�>��>EiR>��>�_>���=����5&��������w�A���U�E�*� c(��g?��9��7 �ڽ��;=��<�΄��N��D罱������\�h�ȗ7?��#?cq��y�>�a�� �����B�N>�4��,!�sŽy׍:�R�Q�x�;�{�����g��Q�=~�0�
?���=�R!>���>�~>�bd>��>��ڽ�2�:V=S>�>2�>L��=��>�:>O^=<�3>݋{>��=������w:�pQ�DR�;��C?[�]��E��s�3�k߾�x��	�>��?�zS>ݕ'�(�����x����>�%G�(|b�<u˽$� ��U�>��>�ϼ=ߚɻq�E�w�4�-d�=&��>�A>S�h��돾�o��%�=���>[�վ3%�=p�z>"*?
�r?��6?D��=��>R�]>2��>�%�=}�K>�K>\n�>��?|5?n*?�>�g�=�}`��@+=3aW=~kE�v�r� ʽou���w��!=�����Q=��8=||���_N=�(4=L+�����;&v�<���>�F7?^��>���>cKw���D���S�v+Ľ8@>�-�{l�>8�>?��>���>���>C�>Gy���V��Ԇ�����>~�Z>�$d��~�s�#�.�>#Yd>:HX?�U>?Q�����k�smr=�}>�ϭ>9�>3�%?|	�>��_>�aA�f��8mӿ�$�b�!�肽���;^�<���M���8ǧ-��������<ӓ\>��>σp>��D>^�>�53>%S�>�EG>~ׄ=�=�R�;��;�F�/�M=���UG<��P� ׮�E9Ƽ������U�I���>��>�->ټT�0?��"?6Nپ�����)U��� ���I��!?��?���=�D?�e�>d��B�Q���V�Q�]=�+?hue?��#?����A�=�4��N7����>��>3>>��^�/�*����<9G�;�>b(G?��?�í<�`��Q{��y`��>Ȣ���zΑ?�d?���C����?�x�-�'�ھ���=6Th����<���|P ����5���&�)�~ՙ=?��?;����m����������u����=?FO>&l�=�8?�ؕ=u���!9��a�$����0L>�%?ٳ���S>�,?���>�P^?�b�>��M?��*���=*�3>�/�>F��>���>MP�>���>�r�>��=o[�`h��_����.�ϻ�4�9g%>�8>��3=C:�� �>��=�`D�7� ��\�e�����<p=��/=OO=W[F>��?R:/?_��B�����F���.�@>ŉZ=0�e��迻�x�=��J>�2�>ѐ?[v)?T��>�h<�d��_!����L1�=�?~�,?��?1��=���=�����*���E$���>1�<e ������+�A�@��-|�>��>��2���k>�l~?�DA?� ?����/�+�s�Χ*��(༠�/�nd�>���>r�=��վl�4��q�.
`���1�7^W��5K��=Ɣ�=�a>�>>X�=M$>���<-���MEн�c<
����>���>��	?c�`>�Ė=���������[?�B��cJ�j����i �`u��F�8=��>��?>��e��fP�@����\=����>��?�7�?��?�D �naF;p�A=�q]>�9��_���幑<�>=�]�=�>��o��������Ã�>�k�=E�ƻ�q���'���Tҽ�;̿��y��쎼�$�$p&���<�>	��W�9��^{�=���B0۾kd ���%>��N>�����Jv��ܾ��y?P�~?�@�>S��=x�G�e=2�LH��>������6="�:�̻�5־_���#��1��0#�!g��K�>�����&�w���I�a}޽M���G?���읾d��~��=M��=��ٽ��D��!��?ۯ�kw|?a%8?f�� �������`>(2?v�>�Z>�]� �0�T<>��/?�lH?r�(=�!��ln��䔼���??��H?���=��5��I�X�9�&�>�z�>U~�>%m�K��#��ـ
?&5;?��p>,���s�.���� ?K�Y?[�6���S>�Y�>F��>�ď�"��er�=R�
��۾$�b>H2=a�>�E�G�VE<QG�>(K�>�ڠ>?Kž�'�'%�>aѥ�;[��������������&?٨����.\>P��=@�8�S뎿�_�2 �=��X?�>�?՛H?�~??9��h�*R���Vؽ#��>�d�>*&�>����G�>?�޾�g�m�+Cھ
�?��?��?�у?/
{��տ�ٟ��o��`Ҿ���>.H�>5,?�vt���q���=x5���6�^z�>���>��>��]>��>��=���=�����������M�I�Wd�����ou���r&�%���L&����\�þ�C	��md��g����<�MG���a�s���`g޽D~I?�S?�?>`]�>j�f�M5�>0�jT��K�t�6�=�]d+�<��dk�@�T�������b��n��=�W���>`W>Z;�>��$?_�F=?�>xH�>��<�D}>��p>=�1i>�<�>��>Ã�>O�>���=�{>�و=q'��$����:���Q�5�;g�C?C]�9*��y�3��b߾e���̴�>�M?o&S>U�'�����x���>8�E��Fc�p�̽�����>���>�M�=�����)�9x��b�++�=���>\�
>S�b�O폾���r��=��>���(Yw>0��>��%?�E�?�.?l=Y/�>T�2>G�>��5=�>C�>��>��?�I*?"8?%�>�!>��^�2������=d�W�����c��l�÷��34輩���-�=��t= ���4��`cV:,��,:=Z�Ƽg��>��9?k4�>��>C�^KL�VX�h���W�?>r\ֽ�I�>�§>P(�>x��>!s�>��.>pȽ.Y������u��>}2>��q�B1p��F�m�>�+>3vc?FD?ҽ�=���='>�>�>��?6�8?m·>IF�>��9�����mӿ�$�:�!�tւ���Zq�;�<��UN��!δ��-�����IG�<��\>?�>�p>�E>��>
#3>�Q�>�XG>���=��=�e�;�	;esF��?M=.���F<ҬP��Z�� qƼ`ė��L��0�I���>��|�Z�ټ~0?�?�e-���^�ꦼ�B���v���?]Q?�?q��>���=���GH��
E��Q�ͪ>��f?W�?�@e��&�>`�>T��c?�>)b>� �>�I��'s��]q7�L�>zL�>"o?�g�>D�&��Ne���� ���f�>��=;\��I�?AD�?�M ����W{���]��\&��a�<<d�z���jⱾ�*���0K��R<�Ժ�W<������	?N��?	���B�뾉���d�}�a�Խ��>��`>�Ѧ>Nɹ<�q���9��7����zK���k�=ݬ?� ��Mn>���>R�=��\?���>�0?L���t��>�8:>���>˒�>K�?���>T2.?1�>�}r>�e<�3轖7��缾�XT�!.p<��(>��>�Չ>q����X�=9e�=S�轼y\���=���=�tr=K�>�K�=֣l�64�=�?��<?�Nx�q���cʼVN��o=�Hc>�>�ߤ�T(<�p>B3>|��>�[?�O�>�k=��}�����	�@K-=���>�*?uC?|=�TI=J辑�u��N��U��=e<:׶��U��.��$��y.l>��x>������z>?]�?��=?qk?���~1���l��6�݋ἵ"�;8�>��>�B�=,ž��2�۴p��[�6�&�M#��U��/=� �=�/>}�G>K��=_�
>C�<`�ܽ����;��'�i0�>���>��?QvP>!��=$F��w���8b?��9���2�����ۮ�<섾`m���+�>�B=Xj�=2���G�,�xT���]�c/�>�d�??��?��?����˪���>FH�>E/3=���q轺�]��'\=6�L>P��=Q4����c'��7>�ML=���<�K��r�����d<��ɿ�)`�w������������bm���H����۾E)��k2	��� =���5_���ꆾ(��4?��vƋ?�9�?bt?j�>��=�;�&�Ueg��ߊ�ɞ���t���2��ф���X�uC��]a]�ۈ�}�P�~A��p�}3�>�B��H���9y�lI��_y�E��A�C?�����QU�i��T>V�=T��?�5��M���џ�,�����?�#0??���T�����*>�Q#?��>�s�>����h)��?2�__?��I?�h�F+x�}�b�g�u{�?�۳?��O?L�>|S^��2����&�f>���>��>��=a.H�6�Ǿ�3 ?��>8��=�(2��ꇿ��'�?\�?�R��{\>T%�>�y�>4�~��ƻ�c�$>bp
��ޤ��\5�
`�=����һ����8D>�d>��>������
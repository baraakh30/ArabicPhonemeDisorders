�   �   lG�=�㥾,O�D� ��!��q�����>q4�>��	�`<{��=�:%߾��S�ɼ=>������= �@���=�i>�>��5>���<:ټ��YT���/;��.=����Mt����=��#>NY�=�pj��^�=��=�ff�|�׽5;�=��U?�A?�K.?�)q>�b��K���&���׽����%�:ͽ=���>i�۾�.g�B�¾�$�C<��3��N� I>j�>>�>{�>C]q>�B���@&����=/<Ž�I >Fk>�:>��x=u�>�UJ>E��a�w�f�յ��&b�] ׾y ޾a3��Li��s�=p5�>'����
>	:����;�З�-�>�Mh>]�c��>Q�=���]yȾH��A� ��Ӿѷ��L���a�;�r��X�=��������n��C�5���T�]]{��O��Z5���|�>���<ޮ�>�WK>��?(�?T�=��B/?���=$?ی->6i&>jH�>?Y�y��>T��>�S�>=���7Zw=V@}��-��@f�j'��Zu<�%[>�++>�K3=�>�=�ǌ=t�O��������� ��i��f�a>U$:>@s�>ӷ�>�*>,���s�����%�>]��X��>���>/Ծ=J�=].���J`��h����F=WX=�̀ɾﻥ�ս��>؞=��=A5>���<�.�:�Ƚ[V�jm�=�N:<���_����2���5> �	;g���rQX����	��<gּ���=K�1?zM?K=3?�� >��S��b��\�n�/��@g��X>��>k{?��C�㾬���{��������<Kζ��̽P=�mm>ʧ�>�">��==�,�퉈=�;����=�;>	��<[D>X'�>ҍ%>���� X]=n%��X/�Zѿ�h�����+7�H��=p�.���0>-A�>�N�R۾¼d��^�E�н�� <U��>���>�g>��=���=8��=�q{��h�2K��'P��$U�<��q>�a�"m�����[�,��x��E���2�v�w��P ���j�����%�?�~K>��=%o�=#�?��>3�>>� �^a>��>�Z>�cx>Ů��%a�>��?�j?��>X�\�1��d�������jl�D0�����%>���<`�뽀�"<��>�z`=?j>�l�:�P��L�>���=O> 1=\�>t�0>S >���@�n��;�3�;�>O�>\A��0i>��p����ዲ��]>C����ľ��vѽ��lO>���=e9����Խ�Z�<�N�<�彩�ѻ&1�=���=�-�=��>!���p�߽x8���	�Ow^�w]�=��;~p�>�MR?_!?{�b?(�U>RþU8��[�����	�Ȼ^��>�v>���>�"�a�h�x������M_���������]�>�/�=�Ê>�.�=��=���=��f����=�=�>=�9=x��>O=�>$r>o�Z>$-�;/�������h-��#T�7�&�x������c��=�yb��ƾL��aQ���8�d��k8�ZB+�웽#�7>=�'=y	��鉾w�(��<���<��ɷ��-5����'=껋�0�=C^�'���,�g��y��
�W��b~�?�8�
��������>$aȽ��">�4���>qy�>�>�q>���>�|'�ω~��P�>y@>�[)�RV�>�?�2�>2c�>��l>�+���-��Ϧ;��۽�EB<a��=��p<Z�>q�?�l_�����n�����F���W�=z��S�=]M�=���=A,�=Jh<��<�y�Ծ�\N�+¾�d�>�Z�>O����˾V�)����2��bɽ+h˾�v˾\-�=9O�D��Wp�>�>�O=i�.>��=[e<�8���iB=���<��a�������� �=,a���t�=�Ľ�\�8N�����c�>X�!?���>и6?ݱ>c�zz��ɾ����s�V>��l>-�<;�>�@½Y�߾��B�c������ƹ�:G3z>~*�>��w��Ԅ;���=h�d��|�XaѼ��=.zq>T��>��>·�=
>�cq<JD��\z�*�ͽ�]��ܖӿ����� ���O��I�=0�<�?�� �Ӽ'�O=��x<h�d�=���D2�>�>g]�=�/>�7b>;��p��5\���������/��!ӽÝg>k�ͽ�����o��?g���j����磩�V����=h�<?n)�կ>��=�:�>_$�<�		?l�?�V�=�b<�z�>��=K�>�,�>��,>�>���>��>���>���>v�`>H�	�)�	9���H��\4�<>z�>|�=���<>�L �}2��n(���ü��Վ�=SL>�9�>���=t�0>S >���@�n��;�3�;�>O�>\A��0i>��p����ዲ��]>C����ľ��vѽ��lO>���=e9����Խ�Z�<�N�<�彩�ѻ&1�=���=�-�=��>!���p�߽x8���	�Ow^�w]�=��;~p�>�MR?_!?{�b?(�U>RþU8��[�����	�Ȼ^��>�v>���>�"�a�h�x������M_���������]�>�/�=�Ê>�.�=��=���=��f����=�=�>=�9=x��>O=�>$r>o�Z>$-�;/�������h-��#T�7�&�x������c��=�yb��ƾL��aQ���8�d��k8�ZB+�웽#�7>=�'=y	��鉾w�(��<���<��ɷ��-5����'=껋�0�=C^�'���,�g��y��
�W��b~�?�8�
��������>$aȽ��">�4���>qy�>�>�q>���>�|'�ω~��P�>y@>�[)�RV�>�?�2�>2c�>��l>�+���-��Ϧ;��۽�EB<a��=��p<Z�>q�?�l_�����n�����F���W�=z��S�=]M�=���=��==q���*��������1 ��i�r?9+j�wH0�fָ=������y��\n�>^=�=��T�%k��Z>T��=>=O�N��Pq=B=b?�����Y��%0>�O=��g���=�2=�jѽ��J>2Ʊ���#����<��>�9Y?��b?Xy?Ӡ�>�=��\P-��FW��V�;O�r>Q[>��>ħ>�c��x-ϼ<bA��/1�"_�]Ъ���a����>�N�=�q!=��=Et�M�g=�ש=��V���U>�<�ʊ>�R�>�]�=�X2>(p�=�6�=��=\Ҽ�ÿJS��ˠ�Yj�v����|��F��#o���S��Y��%=���$d��>����<���g��{��=3�=@��[�Ľ2v�~�`��Ⱦ�Ὡ�X�"�=�3���ھ� �!O>����(�%�rpS>���� Gh��T���m���>�<1>��a>±�<�D?mC?��/?�7���G>��>5�������Gx�>"��>��3>���ܯ�>@5�>�Q ?V	ܻo�W�_�j���
>)5�=
s=ۆ�=�l��8>�>�Wd�1Ӫ����~I ������ǽ#��=��=RdD=��w=����׾ �	��.�)���>׽U
?32@���a�uZP���������r��۾ҿ4=��$>t�y;�~ɾNs�>�LK=߱;�wj����=e'>�D}=O~~�u�3;��>�3�["��k�}�a���=�ք���r�q깽ƞ�=��z?��?��??�
y>x��/{R��|�P8<���<\f>�)?��>�q��sQ>�A5�x7��0��8�+�p=�4�>u#>�Y�<�U>~a˽����A�=�=���F>��I>���=�5!>���>ӡ?>�%>���<�(+=8D��OSv��پu[�������������%�=�C��&��*�s�D�g��O�?^�1q�=�
=��=��>m0m�n�����žr�����=���~;�طe���#>H�k�(�վP�=�r�����f�P����﷾��"��̽Θ���>��ݽ���<��>� ?�I?`?��[�3�#>=N�>�&�=�x�=1��>���>��R>b^��|�.>�ԕ> ?g�콛U�&�=�N�ء�=4ҍ��>��׼̲=�罩���V=�p=�%<��>����<�R�>�A~>&T�=<W���Ͼ��A����')]��B������<?ԻѾ����Y��۞����%�t�������[D:���(���%��J�>!����[X��꘽'@�<Ѥ�=��>
n޻�ڃ�ڰ<	��=�<>���Iɻ�u�� E9�=Fܽ��=b�*>Gr�>/q?ߛ0?�h
?+b�=Mn��V4��{C�_6���O=R^�>�#?^��>*�\>�֟='���F� �Of��}���P|K�>T��>��>|/>�a��
�ҽ�8=9�>�O<�#��#�w�=E�R>�Ci>$`�=�m�=O���5�����R�p�%���d��P �Ȏ���\8�]��nӛ=�{޽ʀ?�X>����t���G�0q\>��=�cͼW���*J�UO���Lֽ2�ܽ������ƾ���=)�;@��_�.�g���]���&� �K�&�f��X����cDs�:+�>�>�>�>N��>ٟM?�=9?`<�>[��Ez�>4?�[���,<S;�>�p�>���>��u=Dy�>�x?�?�S}�A���E<ٽ�=� >�x�<2����>���={۷�:ཟ�p=�O�Q���7o=�	�=��X;��=�@>qR�������ܾ/� ���꾰�ؾ(�?O�C�y�N�;�*>?���8d��9(��Ծ��6>*�f>]&¾_�
���>����ҽI�
>T�>Q�?>��1>g9�Y򦾨� <�>�o���-��=4a =��l����<���<HuF;1
e>6�3?�8?4��>$�>������þ�p �OS�6$>K|=q�>�S�>R�=W!��W��:A��B�������&��?P�d>b����=�r`��͜�,� ��c�� �Nؽ>�0\>�=>���>_Zl="4q=�s.=(oa��G�ڿ�Ѝ��SѾU��6���������n�r���8=&?��h��jBb�Ĳh�_��<?lJ�����xa�e9�=~�=:~�>ԋ�>q�ٻ��=�"�ӈ�k�Y�=c0>e#�=��޽[�$���>�&Ȼ7�d��"���P�R:2�Kuk�͸
��*�>�n�>r9�>G!�>��0?�7D?2�(?p���@�Q>�/l>;�Ľ�̂>ES�>"?]�?%���
�<%��>
?ʭ��ta��0�K��2���'�=��,>Ā>=Y輭��>�Ii=�\��O����b��=��=أ>�K�<`V4>�T�=Q;�=�C��N������c�8a���3?b���{7�5�>Ӷ��s��Z�þ�/���=-��8��>��=�y��4��>4}�=�K�����[��L
>Fd]<9n��mW��o>�`q=��<^��=!��<�e�=��=�����X=���=�Cd>ow?ӄ"?6�%?�os���c�Ŋ�Ƥ�0��=+�*>��=�w>f>N����L���o�N�p���
�����=��4>!��=LJI>��$>�z�#���:ؽx�=jsռ��P>-2�<m�>G;�=Q!>߬=^'];W�W��?�]'��J1��ڿ��H�+�X�����(����w��<��n��`��
諭�4����b�<%��ؗ��1������*B>��>}���q��V��%��Mm���|�g̑��<�JZ��D�L�x�^�o�5��_��!�0��Z���͇���¾_��>��9>��=�r%>-��>\:?y�?�[�Ρ>�{������]>��>B��>�Y�>\�>~[�>!�W>�Y�>���� 2��O�=7d�%�<�˝=�|9>j��=��=�X��rѽ�y�=�n�D�~=��ǽ�S��D'>��U=�#Q>��>��>���P �F���叾/�=��$?�Z=>2o��K߾�< ��ξh ������g������E���{\e>/L>�I�=B'z;I�m��F�����M���.ܼ�?>�R���3�=�E�==@L���	�s<O+��:�<L=�I�>JY?��Q?�%?�酾�V�
�i��p��q�<�>l>i�^��@_��>>y&�W,�e�8�ʁ�����+��=��¼�J>��.���;���	>z��_~M���=}(>a��L�=9V�<��>F+�>�>8��=K��=t�J�����T��Irۿu�����*������H.�$��G�<��4�������a�>��?�V�>��>Gm�=�u�>�.6�=W��po��ď��s˾�"Q�ʃK��)B=<&�d����uE�1�Y�ʏ��@7���������H���]P�ܨϽ��>�
`>WI�=�L�>jE?uJ1?L��=G	>�L(>�匽mt?w��=m�P>�!�>$�(>��>3�?�]�>4D��ٷ�Z�m��.|=���>� >��^>��j>�������+qм���=����kI����/<ҩ�G����H�=/[>��s>��>��>���P �F���叾/�=��$?�Z=>2o��K߾�< ��ξh ������g������E���{\e>/L>�I�=B'z;I�m��F�����M���.ܼ�?>�R���3�=�E�==@L���	�s<O+��:�<L=�I�>JY?��Q?�%?�酾�V�
�i��p��q�<�>l>i�^��@_��>>y&�W,�e�8�ʁ�����+��=��¼�J>��.���;���	>z��_~M���=}(>a��L�=9V�<��>F+�>�>8��=K��=t�J�����T��Irۿu�����*������H.�$��G�<��4�������a�>��?�V�>��>Gm�=�u�>�.6�=W��po��ď��s˾�"Q�ʃK��)B=<&�d����uE�1�Y�ʏ��@7���������H���]P�ܨϽ��>�
`>WI�=�L�>jE?uJ1?L��=G	>�L(>�匽mt?w��=m�P>�!�>$�(>��>3�?�]�>4D��ٷ�Z�m��.|=���>� >��^>��j>�������+qм���=����kI����/<ҩ�G����H�=/[>��s>l)�>����w⌾(����F�߳�Y��>��ݾ��=H�v�/��՝�������x��D�-0�Ӟ>,�>9e�>%wU>N)����gG���= �>E��<Q�=�v=3���,��������=8�Y=��o=zVj�)z������Ϸ�>t�"?�xY?��@?;$�=���1���뾢G�=�F��`�F>�>��
>Z޵����~��:!�`�q�'��n����>���>w��>�~>ǈ��ƀ�����v��=�!=J�<F����a�>;B	�𾟽G,<�,R>���@ڽ,s�o��Oi4��&޾7�����k޽�<�
����=(���W0> �n>�7����>Z��>�?$7]>�=l�����j��.�'r����C8S�%mt��c+>.?�R�A���;��<Ox_��U������	��~�䩯<�+����>���>�C=��<�D�>��>j��>U�>�<3?R�ƽ#$�>^?��"�=�b?�&�>2$?���<�A��\y���:�
���h�:���=�$��\�=�{+>�X�<�?�=�q=]"�<�D<.{����=(=^=3&�<a >���==��>��>���P �F���叾/�=��$?�Z=>2o��K߾�< ��ξh ������g������E���{\e>/L>�I�=B'z;I�m��F�����M���.ܼ�?>�R���3�=�E�==@L���	�s<O+��:�<L=�I�>JY?��Q?�%?�酾�V�
�i��p��q�<�>l>i�^��@_��>>y&�W,�e�8�ʁ�����+��=��¼�J>��.���;���	>z��_~M���=}(>a��L�=9V�<��>F+�>�>8��=K��=t�J�����T��Irۿu�����*������H.�$��G�<��4�������a�>��?�V�>��>Gm�=�u�>�.6�=W��po��ď��s˾�"Q�ʃK��)B=<&�d����uE�1�Y�ʏ��@7���������H���]P�ܨϽ��>�
`>WI�=�L�>jE?uJ1?L��=G	>�L(>�匽mt?w��=m�P>�!�>$�(>��>3�?�]�>4D��ٷ�Z�m��.|=���>� >��^>��j>�������+qм���=����kI����/<ҩ�G����H�=/[>��s>l)�>����w⌾(����F�߳�Y��>��ݾ��=H�v�/��՝�������x��D�-0�Ӟ>,�>9e�>%wU>N)����gG���= �>E��<Q�=�v=3���,��������=8�Y=��o=zVj�)z������Ϸ�>t�"?�xY?��@?;$�=���1���뾢G�=�F��`�F>�>��
>Z޵����~��:!�`�q�'��n����>���>w��>�~>ǈ��ƀ�����v��=�!=J�<F����a�>;B	�𾟽G,<�,R>���@ڽ,s�o��Oi4��&޾7�����k޽�<�
����=(���W0> �n>�7����>Z��>�?$7]>�=l�����j��.�'r����C8S�%mt��c+>.?�R�A���;��<Ox_��U������	��~�䩯<�+����>���>�C=��<�D�>��>j��>U�>�<3?R�ƽ#$�>^?��"�=�b?�&�>2$?���<�A��\y���:�
���h�:���=�$��\�=�{+>�X�<�?�=�q=]"�<�D<.{����=(=^=3&�<a >���==n��>\�����=���_��=��uټTZ.?���C�>��p>8)��ľ)d��++���+��w>�?F?-�?V�@>֊༃tc�A�=桶�9$=�@�=+��@��U�<�Z�	=_K_=�^ ���/��aI�U!�=���=\=�9�=�>�)?��?�*?}�G<�;��U-�D]%�y:���˾Â�>�d3>�h�=>���IS��󺾺y׾o�!���4��=+r>�􌽌���p�=Ѩ�����k��=ܒe>�~��X��9F�C=��>I�>Z�
>��>c��<��%��}�����<���i��Ǻ����_-�\����پ/N�FU-��_���jl���6>��q>Ơ>�d>Pd��N�=Ǳ"�n�;�?C�����9g�s�8��΅����<,���ީ���V���x�Z�!��.�?`h�'J�⎍��m:���.��ʭ>-��>Bԧ>��>[%B?��B?��?%+f����>1\;7n��fq>R�>c?�C?��n>+Nr=��������k%���=� �>�ڱ;S�	>��&>0#">Z�+;߆�=���>��=0z�=�g�:e�=j��=�*���6=�I><�N>� �J���!�{S?����c���k=��>������=���I�=�������r�?���N���?��%?�S�>�w�����<��{<UԳ<�����=��H������X�'�����>p�	=*�=�-������Ƽ���=�n=�]�=-�?�?̣?x�"�k>㾥g���Q�4���G��ZA⽎6�<q� �W�	>�T[=:����� :%��W�E�D�Ps�>���=��&>�|>��n��+"����=��h>>W�kY7=�6�uy�=�3`>��>�>�&�<̩,�1n1�����f�+�1=پ^c�C%B=�Yy=��"=�	�h���a�� �� 4!��G���r(�r�ѽ�Q㽩�����=i]'�%!b<{'��"Q߾�f�گ����}�T��k��3��0ž�݃�Ĭо<��̖���Pz���h��� ͞�t�>�m�>�X�>�'?��,?�Q�>�U�>�R�=�r?���>z��>�P�Ǖ�>��>"B?;2?<�>&�C�o���<܆<\��;5�<��C=Z��=�g�>�̎=%#=؎(>>> �= |�gV�=jb ���Ѽ�Q�=s�=�><L,>�z�>�|>�H8��z'�O��;���є/>�1?��:�*��=����S���� ��P_���Q���O�-M=�iOe>Ӷ?�5d>ـ.>��=S��djI��
<=��[=��>"VĻ�0��>L�o�l����=�X�<KS ��O?�%���>��>H�>��?�>Z�?��������,�f�����dj���DE>���=�h=+o>\�<����6Ѿ��	�pZ쾈Qͽ/Z>'�t�9�=��b> &��Ŵ��Ww=��%>��v�@��<Q��J�G�R�m>h��>��>��6���>�o]�)��N9翧���� ����5{����׾��r���D�p���'¾H�5�	Zq>�_�>E�a>k$�>iT@>���=��->���d�%�x����#�o�� ��%k�b� ���8<�y2��6��$���?���!SY�����-	�C*�?F���hb>Pf�>\?��>�y&?CY?p��>zF��,?A�>��>��b�D��>����n
??�ʎ>�^y=��q��m�v���j��ܕ=�bI����=�&�<�U �� �e�C>��>耐=֙�=b��kۓ�p<)<;�=p=��=R��>�������)־����>��>�9�>Ԍ��ɯ��^��T���5����^z<�9��`��R�����R?5�;>uN�ܻ/<v�=�q��㽂؄<Sw�=�z�*���$��$�=�q=�u�>�P����4�#Z�==!�=�p>APb>��B?�3�>,7�>�O�E��v��c-����^U ����=PD>ގ�=`κ���%p�^/���4��������t>a9���ݼ5#�><��<8J��J���i%>d�����>�h>;!m=�c��(�?��>Z��<�3���O��|ſ���z;�1~��� �����G�8�X=#x�#xؾ3�ϾZ�:�<������=�ه>�|�=v� ��Nּ(��==Ji>�ʽ<����W��bX������97�����G�-@��_�1�s�$�l�Kڂ�~=�i��"�K����.�>�6>6$�>��>o?\?�j>�>���=Rr?!y>j��>m#�>�T>��<P?'?a�2?1'�>�H���W,�%�p��!>��{��=� Q>ƿ�>��>yN(>��=x$2��F�;�̚<��Ƚᢺ�AZ>""	>w�:>���=��w�Z$پ6��������=@:�=�x>�P��	y=A���s��W�=���D}ʾD�l�4����U>��G>c��>�s����u�e�<�p��QA��}�>߽�։�1�h>>0���X=҇�=��=�g=�!���3�@��]�>yM>6��=�
'?_/�>Ȫ�>`�)>�p�e�����cսȭ=�2����9���� ����m>ʽ3iY�킲��tо\���R�O�Y�#>17>�����=&�=��H->*�>��\rj>wqѻ�t�<#���da�>?6�>6 >�t��<'� ��ڤ��p	оk��됈������:��72��7����@�=�އ���g�VL��hM%='A�=���=�؞�g��-�*�r��=�~��[n=/Î�uWs��9��,\Z�Щ���¾\���FԠ��:���"��@o����ݾ�kѾ�J���e����>��>�I7> ��>O?�Û>�.�>�P>���>���=k�+>4�y>j&�=@S?�0�>� �>-�>�>͋���j:��r��,�=�y�<�Qa=(�*=���=w����,H>��8=` ���=�@��޻��8=17�<�U>��;�;m:�$�>U�<>Ջ;��`�k�Q���ɾ�ũ>`��>�ϾY�(��3�Ȣֽ����Y>h�|��O4�L_��\, �����>�~f=��b�30�����<��=B��=�k>��*=0�==��H=K|d=�ע=���=��=$ƹ=X��=>�<v�ǽ�(�>�_?��?��>ʆ-=�v�L��M�۾r�ھ]��=KW.>��*>���>�\����"���쾆9_��
��j���=�W�>f>>@��_������i�S��rT;�;��pA=���=O)�=�3�%^�=6ӷ�=?��,ؽ`F��(򿖊�� LӾ!�M��4&����{8������1����<ܘ��>'���<��F
><�(>3G�>��>(�>rS�>�q��AQ��1u��㟽�P������2�G�I��;��6�WH���͝����`�Q�ڴ��7����8�H2c�C,���W��1m�>ȮV>d��>��>f +?�f7?��=q�=�Y?̚9����>�<�<Q��>�:��Q(�>�e$?SU?5��>�(J>SrB�������=S=���=C��=!�>QX2=��>�|�<��=��M��O�1����<E툻a�=Z��=-�O>Ox>��������Q=P�� �u�N�>
��=��W�~ǻ��ȾQ�Q<�����(���=�p �z�ͽj���Y[��ޙ�>���>���
�����c=(��=���=�*�=;B���	Y>V��Տ;ݞP�����yf������\��)�>��!?�?SR?��'>�/�G��^���K��6@�=a:b>��N=D�>]WR�Y�]����I*�`�W��G-�����n#>X��>�ov����>��y��Kʾ6ʧ�&L��d>D�>d<�A�>��>^_#>vlO=
�=�������p{�Fr���?��ɷ<���Z��Iѽ�:�<�Lӽ����I�������⾵a��4�,��S>�x�>��<uؾ=z~>��������xq�W����J���P�@��o�C� ����� ���л ��uS.�!?�=;��a�����®����>�Ҁ>��>dБ��I�>l!?@�>��$>+�?u��=:�>��2>�(h>.!�>1HL>�c�>| ?�ҥ>)�Y>Ӗ���4w�J�ڼ�Jq>J+�=<��=mv>8��=N��>�jd=#��<5z��s�۽ Y��Z<R7�=ɢ	>J�>�ɋ><�=��@>��{����_����>���>�_ʾ�G_��߾�Ӿ�޾��D��,	�𧖾?����A����=�ш>)Ɓ>��ɼ�*�D�<�p#>\H>a�S�8�ڽ����j��=��I>h]�_O����;�؊����+��+>l�>,�;?��L?��?1�>q�*���+��u4�y����D�<~�>rf�>\}>�\�����m`�sϾ������<�l۽�e.�d
>1>�s>l�<�k��BҸ��[>1�:>:�S>u�T>��>��>��8>F�>�c�>T�r��o���ɬ��ӽ�V��x���&�����3��Mwｐ,)��o=�s���P=}ة��K�<�X�=B�>��D��Mn��G[���� �5�<�W��G��`�ۂ���谾�:��ֆ��� ���������Qգ�G �2ý�䒾�w��Ъ�Zc���'?H'B>�.>��`>ޏ?�~=?*|#>�?;>ŧ/?��T>�2j>&��=�9�>��>���>�?�0?yv�>Z�{Å;9��Lg�=��^:>zl����>��">��=�����w�=��G�s�M��z�=��=���f�=.�Q>�+<Ox>��������Q=P�� �u�N�>
��=��W�~ǻ��ȾQ�Q<�����(���=�p �z�ͽj���Y[��ޙ�>���>���
�����c=(��=���=�*�=;B���	Y>V��Տ;ݞP�����yf������\��)�>��!?�?SR?��'>�/�G��^���K��6@�=a:b>��N=D�>]WR�Y�]����I*�`�W��G-�����n#>X��>�ov����>��y��Kʾ6ʧ�&L��d>D�>d<�A�>��>^_#>vlO=
�=�������p{�Fr���?��ɷ<���Z��Iѽ�:�<�Lӽ����I�������⾵a��4�,��S>�x�>��<uؾ=z~>��������xq�W����J���P�@��o�C� ����� ���л ��uS.�!?�=;��a�����®����>�Ҁ>��>dБ��I�>l!?@�>��$>+�?u��=:�>��2>�(h>.!�>1HL>�c�>| ?�ҥ>)�Y>Ӗ���4w�J�ڼ�Jq>J+�=<��=mv>8��=N��>�jd=#��<5z��s�۽ Y��Z<R7�=ɢ	>J�>�ɋ>x�u>�_>���H����[�^�u��?�;;��>S\.��s���]�R��7�zPǽh����,��]���ώؾ�����>F�>)�2�(�=�#�<�`�����b���$>��:�m!>�>�(�=�T�=�:C=�Y��F>�껜&���J>�Z(?���><=?h]�=����)Y��6,��׾�_�>BL�>��g>=�>��g<�׽W-����O�����p>����=R��=��s���=�?���Y=G��������=�W�=I�=�=�> �^�xR�>
�y>ؿ^��l�OHнi�ſ�4���,߾7��y�=��,����=Ԡ��=A��νZٍ�|Ȫ����{(A�}1�=�>�=��h=��<>+%־���h�ڽ��S�e�Ծ7E��7�E��ƽ�*��#܉��ƾ{�)����8�����ξ,�=
績I��e�-��><��<�h�>�L�>f�?��?�պ>�3�= ��>���=���>��>ql�>za!>�s=R�>_~�>0��>ٹ�>��H����f�>F�=P��=v�k>M9>���=�u>��=���<�Te�'��)�:C�;�z#��$�=��>�{1>�X�>�g��,�>���"�,�A���P>40�>�g?o��8�o��gQp�2y��8�����?���k
����>>��=�|>�,
>Q	��)D�=`V���?�&cٽL ����p<l|�=".�z%����+��V+�:�'�W����������=81�;�-Y?G�T?��5?,"$>y�o���j�~5A����>�>-��>8��퐻j�Ҿq��ƻ�n�nE ���<}E%��	�=�"�
#={����MĻ��e�g>��=\��,�#>���=�4�>#L�>�F�>�8>�<\;��M�e�\5뿊c������ ��>�D�=��>�c��̚�ya#�؂�{������<�A>��,>�z�>��>��>�Z=`��>��<m�3=�נ���Ͼ�2��Ԧ�ʼ�>���E^��|�s�Z�.>����ć��
���D��*о�O��H���g>NB>��0>i�>�0 ?�H�>��>2�y;�E>��D>��>��=��>!՘>�d�>{�>��>��= ��3=����M��_>a�(=��W>`>�� >۴Q;�;?>�W�=�=���U�=��=����H%��,V>?5>h]>���=6�>���=�&̾s�������%��s�>Kd>������Ur�W1�>��z>���	խ��{���>Cu1>:Z�=&��>b�%=���5V�%03<�*<��P>�:���>�0��w�`�7Z�<8y�J��=�"̾9���(��@�e>���>$&�='e?�@�?�QM?� ?$Q5���u�r5Q�g��7>qD�>4�̾���.Q��d'�Pw�"2���`<rRѼƲ����5=Ix�=~>�0A='�;:�ｚ��=����"�&�>^�*>)u�=��n=qe�> �=r|�=�*��Cw��@ؿ=��^�����a��=�gͽ��K�.�V�i��='�Ž�ʣ�e�5��i�@�h>��D>@ՠ>x-�>��=	 J��x(�s��E���-$������k{�9�P=Ykz��⪽�6����5���}���: �c��p������1�ƛ?�*<�3�Weξ�,;�"�G?8�?x?b>J<A9�=M�f�>> �M�?7��>K�>�f��ʥ������Iq��H�p�=�~�=��J>;�>��G�o7��o����J>�&�=3��U»C�����<��_>|&>¯	;\�j�o+�>�~����R���*��->��>��>�<�=�.��ڬ�L�ƽ)�9��(�=�]�<��/��۽t_=,6�=�3x>�q��4�=A��:M)<�`����=Ob1��=@Zܼ;�`�I��=�:l��s=�-ξ�H��O�<�'�=:s�>���0T?��L?![?���>�G4��/V�b�K�W�����>��?����t��VyA�s!��m>>�H�W�欿�^B۽ۧ���A�=6(A>��p>��޼������L;k��Nڽ���=l�%>�o?=N!�=���=/C��Pu�=AM���Ͻ�b̿S���D�~"���Y��ؼq�&>�:�<^�;{�=��L�����^�ϜC>,c�>o�~>�����ܼ�zŽ�ܩ�I�=����߮ƾ�*������#��w>sd�����1־d����C_�I����=��ν�c��N���`U���ؾ>��B(���dW��>iG�>��>���>�~�=F����w<ɍ�>�v ?��?8c���&���=�c�>�ݔ>�,�����<ظ�=܋=��<��>�K=ɗ<�qG>�n2>�f�=��4�O�=�錽KC>�g>�}�<��=f��6�>���=�&̾s�������%��s�>Kd>������Ur�W1�>��z>���	խ��{���>Cu1>:Z�=&��>b�%=���5V�%03<�*<��P>�:���>�0��w�`�7Z�<8y�J��=�"̾9���(��@�e>���>$&�='e?�@�?�QM?� ?$Q5���u�r5Q�g��7>qD�>4�̾���.Q��d'�Pw�"2���`<rRѼƲ����5=Ix�=~>�0A='�;:�ｚ��=����"�&�>^�*>)u�=��n=qe�> �=r|�=�*��Cw��@ؿ=��^�����a��=�gͽ��K�.�V�i��='�Ž�ʣ�e�5��i�@�h>��D>@ՠ>x-�>��=	 J��x(�s��E���-$������k{�9�P=Ykz��⪽�6����5���}���: �c��p������1�ƛ?�*<�3�Weξ�,;�"�G?8�?x?b>J<A9�=M�f�>> �M�?7��>K�>�f��ʥ������Iq��H�p�=�~�=��J>;�>��G�o7��o����J>�&�=3��U»C�����<��_>|&>¯	;\�j�o+�>�~����R���*��->��>��>�<�=�.��ڬ�L�ƽ)�9��(�=�]�<��/��۽t_=,6�=�3x>�q��4�=A��:M)<�`����=Ob1��=@Zܼ;�`�I��=�:l��s=�-ξ�H��O�<�'�=:s�>���0T?��L?![?���>�G4��/V�b�K�W�����>��?����t��VyA�s!��m>>�H�W�欿�^B۽ۧ���A�=6(A>��p>��޼������L;k��Nڽ���=l�%>�o?=N!�=���=/C��Pu�=AM���Ͻ�b̿S���D�~"���Y��ؼq�&>�:�<^�;{�=��L�����^�ϜC>,c�>o�~>�����ܼ�zŽ�ܩ�I�=����߮ƾ�*������#��w>sd�����1־d����C_�I����=��ν�c��N���`U���ؾ>��B(���dW��>iG�>��>���>�~�=F����w<ɍ�>�v ?��?8c���&���=�c�>�ݔ>�,�����<ظ�=܋=��<��>�K=ɗ<�qG>�n2>�f�=��4�O�=�錽KC>�g>�}�<��=f��f��>�ߴ�sc����<�����y=b�Z>Ua�>W0��C<�2T�� $� ����򍾝G���=Q�> p�>�2�>�i$>������ >�K�>[��R��=�|^>��^�!�a��+�������a�8�0ҁ<���A�x���v�>���=XH=��d?�y?m3U?��/�F��D��Wؾ[Ү�:�����>��3�W�)��毈�q�v�h��T ��<��,���n�=qbu�$w9���>�ݖ<c��=7�0>�<v"ܼ��>#_�>/�>��7>�ĝ=����������Z� ��?��G���a�m�.>11�=�����2n�����/���8ξa'>w��=I �>.u]>���o&���>��� =��<b��=��s��In�^��}�����]>^OS�����!�aؼ}����e��	���+��S��"�+�6LŽ���>z��=l�|�ݞ��nf?՟?��?	��"K)?v�?�Z'<�>�[>�?%u>76+>"=�;��6:>�g��.�;l�=���)�O=���Y�X=n��=�܃8��5>�@�=E���#������m^=��=hf�<�v�������>/ꉾ֦��CϾ����^���T/q>$�>9�˾篽�����pY��ԭ��l<�?>��>d�>K�>i��>I=�HW=fh��y�����=���=J���� =�G=G����G�=�����i�uO��}<޾l=�?>�g>�T�=~M3?��4?�A5?����=����#���=�%>��> �=���=�x��۾ϭ���n;�Q��?
���H/�X>�t�<]e��I�=���o�½9�	=x>�Q�=f� >b�#=tF+=�L9>�t���LM� ��}����7�c�2ؿj	��g�;��弞v�<�/N�i��mG
�8Xu=s�����IZ=��f>��>Q�X>a{�=���=Ś�=�����Ƕ�*0پ���'8-��k�T���]�=t{�����Ր�B݊�<� ��9ϾC�ý����y�D���[[��c>��~>xo�����T?/	?���>�Cj=wص>��������>�_>�v�>�/>O��<XQ=�� �܇o�1Q��s����=��n>|�� V�=�U8>^:>�~�U�ս�缏� ��i�=iL�=�\>���=s�=cm�<��&��>5�>>�r.��S��_:E��F���-�>1� ?N�z>9���R������齺}��B�=�=�>AF�=��a��$��*�r=κ-�܉�=.&�=p����������=�ı��5����=�߮��ؚ=".���C���<,�o=kj�<�q�<�A�>#,�>��Q?�:?UTо;���'H�P��!�h�;���L�>t��>���=���iUC�f@ʾV񮾻�m�����=#>�{�=o���>{>$��=�d�&���t8�>�~�֪<��E>
0Y��<>4z>|(>]��=������Խ9�ѿzԠ��0_�n(��K����\>Iή>v>?x�=D> �%�L�#��n�>��>��>>M�|>�>?=K˼#�>�W>�@��B�<�j!J�VU#�g�?=@�@=�6~�3'¼_ ��.�<O�Tr��-�T;��k�bѲ�u��q��>��>-om>�fU��K0?w�?�}�<Bj��x���=+4�=>��J>Ya>������|��	?�C�>=�ʽ7���e=�p�=�}O=)/�<a�>���֪�=�>� �B<]��R����y>u�B��(���ʸ�=]�>�_�>Qꀾ��½
ǣ�����ֈ��8�s�p>;�ϾUV�>:�H=�n��Q7��}��Xe��>x�_>�	�>��>s�f>��,=R<D�ý��!�r�>0�<�󽽹��#M�=�g��8>h >$��n~��7/����w=�ڒ>�~�>�<)?!&N?!W??䫾�$��a ��9��>�.����>Y�R�$���q�=�ꦾ��O�<9x��,��x
���!�J]$>yi> ��=�	ûh%��-����8�!К>�T����=��=�B����=S'�=�ߠ=)��=��x$�p���2��� �߾פ������X��j�?=�� �=FD���ھx>���4����>�Đ>䥪=����G�����:ھc���q���,k߾�\����I�׭�"f=�#��DѾ>	;��!�蘚��H	����6�,�L|���վQ�Z�$�>���>����y�=���
?D�?���>,�Y>�	�>��T�jJ��J�>���>!�>��>c���>�@�_=�Y>�:%�-����U>�>�����=��>Ƴ��F��=m��=eA��(�f�~=�>��=y�{��6��>d�->??'���[¾����Q�g_��{�Ǿ���>({ ���e�r�,�*��)��qWپ��y�~�@<�t>>�M�>)�=(�C>�-=�68�l�o�������>�J�����5�i�<�>�槼�U潭��=E0���CW�,vr�ip9>�D>��=�|&?J�6?�x=?�ƽ�lܾ���=Pv_�!�����Ⱦ$)�>=��4�e���Ž�xȾ���*Q���Ӿw��í½#��=B�<�;=+J>�Ұ=���	=��i>�?����ZDJ>�h>u��=�S�=��=w�X=I����	�����ne翡׼�ڑ־j9���L��y�<��T�~��:=��޾$W+����<a��>��9?Z.�>f�+>d�8�ы=$�B�j[�<�*��	��Ô{���W�цV�x`#>�(O�Ԇ��@;����L��[��V��`��r��)��V����r�Q�1>\��>�/=4񕽵:'?�?��o>oP>>��>*�>C�#>�}?^��>�>��>��z���}ֽ���>#�0��� �@~>�>�C�li����=�=+�=�I�=D#<���n5��q���ĺ=>�ҭ=��'<c�����>�0���̾-���_����)\��� ?�����ǚ�MĹ>q{�;e������<��ଽʉ���ӻ/M�=9�>�ZC>������K��rڼ!a�<�*>�7�=E��;�=��C���f�;ޔ��Ђb�����|U���&��݄>�x>l1?��?[?U3=,yL�ՕɾB��x���4��>e�[�g����O>��޾0(`���E� %��΀���������p>yj�>�"�>m��>'��=Ig�?듽t�> ��$��<q�����;�n�=�>���>�k\>{WӼ��ҙտ�Qf{������."�WAr�`*>-e�
 ��U>�t|���<=DO���0>g?e>�
F>��>+ �<�B����>�d>@=�=?(k=����
����ٴ8���20�=�[L�9\��?�� $����d�ӽ@�����C>E��}ӽ�F�>g>��r\8?H�=?F?�>�ˈ�>�K=l� ��@U>[�y>�9`>��>���=��>��!>P�ü]U@���Ӿ��i=uI���]��7z�=<�>��=�ؽ���=ci�=Z��=��=��^=�*h=U�G�ʧ,>�U�<'B<���>Ƿ_�t.�[_���㾄<���g�����=���n�/�?I;>H������QQ��۱�/f��-��;��>:qS>���>�*>^۾�.Z����;�'=��o=��>�B>OÞ�u�C>�8n��s�=�Y>���9\ټ�hv=��=��l>��>���>�>Y�?X���<�Z�ھ������e�d*=ylC=����_�_ ᾶ1�������������[���J ��A>�*�>s�6=ң9>x��=��c�.��CB>@n=n��KO>#��<� �=uUo>%с>�Q/�LC�9�z����Ǒ���z��S;���ٜ�u�7<A�>����t�=��>�M��[>��9>Py�=xҨ=fը<G��<�t���X������gϾ�꽲J�=�#�+���沾g��|ھo>�2Y�-8�<�4�w����K��2�n���TQ��h��.��=�:?�f�<3$I��?R��>��>3�>z ?����~��Q�>�?62?�?D�>~'V>W�m���"��P��:۽L";>U;> *>��=�m�>�
�c�n8j>ʁ��CH���3�����m�>=���6��=�u=S�=�M�>�ֽ��<b ���V��F���o�=�4�>��������g	=V�Z�Y����9�=������7�1>�?P|}>uu�>��u<m␾�Tʽ��f==0%W>@}z>(��R�t��:�=�$���<�D��J��3߼�g�=�$>;��=4�E>��'?���>��?-�U=����;!��%���s>��"���>2;x����Q��?��re�����~�}��Ľ�0��X
>1�4>�T�`�>�d>T2����P����>�ZZ>�컽12>��j=3Ĩ>���>v�g=�P-���Z��ٽd⿋޸�+ž�|Ծ��(�2�>�$��	���������>��w��Z.���=��5>�>�d>�f�=����$#>�Ҍ�I�F��g <������! ��������^=� ��j�w=@�޼qc��4�@Iٽ�m8�HM��\��F|��&��n�>�a?��/���(6�>�?s[?��P>��?�=Gda��0�>>@#?��$?0�=?P)�>=�պ���cֽ�m�U��#
<�>M�y>U�*����<�x7> ���苽��*���	��=h�ݽ�{=�
=�X>��a=Kc�=3H�>I';�% ��u*��	=�U�(��Zp=��>M�]�ඛ�4�o=\Cҽ�]�������I����<�%�<|4�>��<6�>1�=u�r�L����^>8U��� �=���>˼�=@{=���>��}>�A=�^>E���mS<UAP= 4>�,>�)�=���>��?�?Qr�W]���������ޓ��@=,��>Y�D���]�,��ibX�^k��֞���f����Y���eQ>�C>�e>B�Ƽ��<W�ؽ����T_>!��q4�@��J��=Lak>�Д>BB6>;@=����u ��Ph�-������g����<�n<g#<����}�q+��C{��ռ$락�2>>>��<��W<�/=x"�<Xҭ�P햾���ٱ���!1��7������>V�˾d#�`U�`ǟ��(f��ٽs:���d?��ċ�[�4��n��i3>�/�>��9��C��D ?��>>��>O]>b0?�=j�H�W�>d;�>�*�>��>�*>��_>�̽��2� d轞����R>Qi=,�=pN>ɺ�=�>:�R�ǽc�n=�����U���ľu�ٽY9&�0�<P[,>R�\>Dx?ST��u����u��󭾱�p�|����s3>�b���/=z,n==���=�㾲d��݅N��F=%E�=�m�>As�=��>��;��$��h���|��=��>�9>"p>T����*=�;Q�߽E�!>VUz<J��d4���=��;o��=��.=q�5??�>�d(?��(������v%�-rоb�u=�@��c=>T>��E�_�t<P$'����O��Q���NG����ɾ�<U>T�>���>�>�=;�+=��ν�r��/e�=�/@��/��%>V�h�ĵ�=�05>9k+<��M=0�U��G����է��;^��/w׾l�!�L'�?�'���+�����b,>�
��b?�X��=E[�=4�>Iv,>���Dݼ���?�>>��>�a�Z���*0���ɾ����Or�=ze���8��p������M�$�*)ν�=D�����d)'���l��U�=�|/>%"D>����	?(?�?��4>��>(O�T�9����>Õ�>s��>Π�> �R�e<>g���EJ>�N���E$�bUY=��c��D�=^M0�@������)mh>�^><�4=��>��m��φ���ʻ|9=����	V>�=�O�>�i�>OU$��s��'�z�>{F^<��*?�VX� �����;�V5>�پ���^T:@ͳ���"��㰾c�q>��>���KdȽ�9�=tEn�c�=��=?>�U��$X��wZX>��m�S�-��<�]k=��D�ތ��0>���=�x�> "?�t*?�EB?5��=4� ����}sǾx�f��䥼Ƹ,?�� >�\�B�?=Sl�{���j$�]�]��^Q�������>��)����<�#?�Q��5X����T#T<T,ϼWb��Ɇ��=��>�C�>$ �>�B=孾��j�O�鿪ȿ�C޾��þ�H���۾X�>�St�UF��AJ?��0�FL >\Q>������>�>��ѽ��u=�W�O!>�p9��q�U\������;��p��'�"t�,{r�#�=Th�<uZ���D=������ž!���>DNT>N��>���=�w�>+�
?���>nsC���>?�=�GὣZ<>8��>�-w>ڷ�>��>�{?*2�>eƽ9X(��@����}>�v��=���0>�ݜ>��[=��>X� >�펼x�Y=�=qΆ�˩2�����Y>9��>��E>��1>Q@c=U��~$ľ*2�M{��u\��g�>��-�?3�=����(R����=p��-�Ҽ�r��?�z���s=Ŗ{>��?=}����̽l*ڽ���=A�=���=��w�A�=j��=_M=>_�A�t1��|��X�F��yԽ�=>3��>�ԧ>	�	?W$~>�:�>�G���.Ц�s���q��ۈ>  �>I�2�U�R�nb�Ƃ߾Q������I��ӭw��P�3��=�%/>�Vk>���=�e� 0L�G�&�i��?T����={I��牉<Z4>��I>q/{>�B >�O��_U�{��뫿h7k�NA������%Ƚ^4�=�n���
I��	Z��=̾��=��>9�b=9��=�9>M��=���#���G�֛^>l�˾�C�BX�U־����O�;�x�;��?6=&W�Ve���^<0E���D���:�Z^������;��%9.>�]�W��>�>)C8?h?��>�(=�H>��b����>��>"\9��N�>�ŉ>���>J� ?�?�������F�M�='�5��4s=�l	>�ji=��;q��=�>����"<�'üG>^�=�m�4�$=���=��>�E�<c��>���>SG�/���o*���>�m�=��>0��=]ξ`���>�����U��x3���	��.M����>m�z>c��ϵϽYP�G�˼�=F=�*>�>/P��=������G=��=��=�<��l{���C����om>k��>�?� ?,�#?�n�T�*x �B�޾������>:��>��=�s��IR�)����ֽz����� �����͠Խ�GH>X�n>��>~U�>Z���c�s�U��J>\�ܽ�7><��=���<>/>���>��k>TJ�<��ɽ$��ii��oʿ~����߾ �����S�Y�,=�-=]�� l��q.��-�ܾ��>`+�=�;�8��=�����f�*=�T�Poh=�iQ�`�l<6OѾ����O���ƹ�<�Z�~��轵Ѭ=�<��ۙ��~�N=d�=�H��Vq���n�,mI>��d���?�l>@<?���>y�>?I���A=�G>�=�>���4̇>&|?]\�>�D�>�1<?��?�����"���#;�L���>Q>��>>z�����:��>��0���5����̼�2�b�<A>>L]>f�D>�=�>�����@�s���!�ʋ�>뎵=�?`�>du
�eȾ�|;�Ի�ܚ���X���꾍� ����=���>e��>:����X��)����|��=�q\>�5A>���٭���<�j5;�$=�]8�C�����H�)�D�{�H>�U>��%>��?�"+?&�;?��$�!65���-O�D���#x�>��?����l">�n���|��j�'�`����,����1��A%��s(>tي<�J>�>,�=�w���9<&O>(���z=�[�=Tw�=cZ=~L>_}1>>��= ����	�#��$e��T�Ѿ=��5��z� �_2��"�J=�\��峾�vI�<R�=���W �=�t�=zּ��=Y��b�4=�i>Mv:�gq�u헾k績��]=������^�����3~�ZR�5&�<������>�������־�.񾁁N>�s>���>Q؊>�(%?�X~>�*�>a��3�+��y�>��+>��=�O>���>�?��>vl3?�p>�=��}E�����wA�=�Xj�E(J����<��q=���u��=Š>�s=�<ܚN�=�=�����>B©>9^�=[j�=�O�>�i�>OU$��s��'�z�>{F^<��*?�VX� �����;�V5>�پ���^T:@ͳ���"��㰾c�q>��>���KdȽ�9�=tEn�c�=��=?>�U��$X��wZX>��m�S�-��<�]k=��D�ތ��0>���=�x�> "?�t*?�EB?5��=4� ����}sǾx�f��䥼Ƹ,?�� >�\�B�?=Sl�{���j$�]�]��^Q�������>��)����<�#?�Q��5X����T#T<T,ϼWb��Ɇ��=��>�C�>$ �>�B=孾��j�O�鿪ȿ�C޾��þ�H���۾X�>�St�UF��AJ?��0�FL >\Q>������>�>��ѽ��u=�W�O!>�p9��q�U\������;��p��'�"t�,{r�#�=Th�<uZ���D=������ž!���>DNT>N��>���=�w�>+�
?���>nsC���>?�=�GὣZ<>8��>�-w>ڷ�>��>�{?*2�>eƽ9X(��@����}>�v��=���0>�ݜ>��[=��>X� >�펼x�Y=�=qΆ�˩2�����Y>9��>��E>GZ~>�B��R0���%���L=oj�>|��<��
?y���C[>���N3L>�뫾dþ<
�^�
���S>���>��>x��>��>]񛾴����̽^�����=��V>7��=���=��&>m�:=I���齀�A�g��=��R>J�>�=gߨ>���>�mp?F3l?������p\*���K��>lI>�����ƾ���>�Y�<�IX>��㾱_<�uv9��9��5����4=��i>���=�NM>�b��S��	b��G�����rz��e���=��>�֥>�>!b.�C���~�C��6�͉��>���
��%��i�þ�zz�C�< &��#/O�y��6�>�I>~�>=m�<&{���1m��}��K�d���T��Pݼ��}�GW>��mn�,Σ������s ���q���;��Ǌ�d��������a��	<%T�>R��>�傽 �޽�� ?"�;>�>|x�>��>���JJ?��>WB1��^>,�d>s$�>2E�>��>>�rҽ��ٽ�j�r��=�=r6�X��=�6�=I�u��=U��<�6>��=P*�=��e=�.ѽ�,��P��=V�ռE\k=!���(2m��S �*	�cI:�đ_���q�f��> S��\D=>q3��#��^��������汾�ź=9@>�b�>�o�>�8�>�-�=�l��0��=-Y̽3�>j��>g+�������>��d=�@�=� ��jD�W��=�1>wK>���=�W�<�˷=�#?8}?X�V?�Q��Ӑ�ޗ��O�L�n�?Gֆ��w����>>��3?f�=�9����E���T�}cO�B��o����=ZR>px�<_�=�����1{ڼ�R><�����S�=\�?>��>~�x>�E=�X���?k�8qL��ǿT��b_��(G޾0�Ի�K�;����ݲ�g(a�>+��ug�E�F���r�K=�7<�A="�w<�����/X>Mi1�Hy�;-q��Ǿ��ƾ1�mG�l����gS�~I�<��}Z{�<�Ľ�l��T��݈ž�7ξ��;���=>��>�[�<�o����z?���>a&	?���><Z(�W�=��>���<	����?>@��>��>��>�t�>(ڜ��#ּrt���-%>�K=0\�=�>��B���i=��=�hK�2�^>�Z!�K�ݼ�%��xk��\�>==C�>�Y�=GZ~>�B��R0���%���L=oj�>|��<��
?y���C[>���N3L>�뫾dþ<
�^�
���S>���>��>x��>��>]񛾴����̽^�����=��V>7��=���=��&>m�:=I���齀�A�g��=��R>J�>�=gߨ>���>�mp?F3l?������p\*���K��>lI>�����ƾ���>�Y�<�IX>��㾱_<�uv9��9��5����4=��i>���=�NM>�b��S��	b��G�����rz��e���=��>�֥>�>!b.�C���~�C��6�͉��>���
��%��i�þ�zz�C�< &��#/O�y��6�>�I>~�>=m�<&{���1m��}��K�d���T��Pݼ��}�GW>��mn�,Σ������s ���q���;��Ǌ�d��������a��	<%T�>R��>�傽 �޽�� ?"�;>�>|x�>��>���JJ?��>WB1��^>,�d>s$�>2E�>��>>�rҽ��ٽ�j�r��=�=r6�X��=�6�=I�u��=U��<�6>��=P*�=��e=�.ѽ�,��P��=V�ռE\k=�\>�8�����ݽ��U��Ú>�t(<�Z>������e>��վD�6�̐;���>Z!�G�=���>��?
O>��>�5�<�y=��(>(ut�wp^>�{��S��3
>9׍>I{3����=3E�}��mļ[8�=�}H=��<I)¼B�4>�N�>��`?�B?��8L6��5������:�>����FT�>�#?��(?��=�?�@jB�ӮO�ߣ�hCO���0�<��ؽ�QH���>b�N�TOU=�s:>+����R�Y �=�>j�w�u>,S�>+\>��=�V�����G������嶿�Mо�.ؾ�V�����Y�=����%˾���A�>G�=w_�<��=�y��3�T��@W=��=�7J�f����{�8�<����$������Y)�=�P�b= �)���Ԝ�8�.�o]/��������G��N�=,(m=��>s��>����@��+?�j�=�����$>JD�<�>�2A��^ľ(�����>h�1?��?[��>�uh�紪����a��,��=��=����=;��=�̒�� 7=�����H=y�ݼJۆ;^Z�t4��:%�P��=G2)>��=!���(2m��S �*	�cI:�đ_���q�f��> S��\D=>q3��#��^��������汾�ź=9@>�b�>�o�>�8�>�-�=�l��0��=-Y̽3�>j��>g+�������>��d=�@�=� ��jD�W��=�1>wK>���=�W�<�˷=�#?8}?X�V?�Q��Ӑ�ޗ��O�L�n�?Gֆ��w����>>��3?f�=�9����E���T�}cO�B��o����=ZR>px�<_�=�����1{ڼ�R><�����S�=\�?>��>~�x>�E=�X���?k�8qL��ǿT��b_��(G޾0�Ի�K�;����ݲ�g(a�>+��ug�E�F���r�K=�7<�A="�w<�����/X>Mi1�Hy�;-q��Ǿ��ƾ1�mG�l����gS�~I�<��}Z{�<�Ľ�l��T��݈ž�7ξ��;���=>��>�[�<�o����z?���>a&	?���><Z(�W�=��>���<	����?>@��>��>��>�t�>(ڜ��#ּrt���-%>�K=0\�=�>��B���i=��=�hK�2�^>�Z!�K�ݼ�%��xk��\�>==C�>�Y�=�fS><Ɖ�������:��rt�����=Gc?U���&U=
Ώ��Z��e�� �� &�=�b>^H!��Aڼa�I�nv�>V�>�8��\�l��!b>�~��J>b�����3�=��	�:x�=�Ȣ�n���R��W�/��!�Ta�>*�>rܵ=g��>4?�P:?��J>��о�A�̚X��Bt5�RA?���>���5������"0�so�Ln��h��=`���@�P>Q׌=��>�&�=�茽X�S���=gB>>I���=
4>��=5��=5�>f��=�=+j�i�C�=���LR��*�}9�.C����=z;ܽx���	㒾m������辍�,����>�{�>쿧��:5�$���������¾D�9�8����Y�%9��k��B������𼑎���B�_��g�#6�=;/�����Ǥ�Q�⾠ӣ>��>.&>�p<Ԅ�>�?�,?;�0>E�w>��j<]i�A*:>|��>�>dac>���>h��>���>��M�R�DW7�7��=�C ��j-<��]>��&>�AH=dۮ=��=��r=� )�7C=�
�=*�m������<>����4��fS><Ɖ�������:��rt�����=Gc?U���&U=
Ώ��Z��e�� �� &�=�b>^H!��Aڼa�I�nv�>V�>�8��\�l��!b>�~��J>b�����3�=��	�:x�=�Ȣ�n���R��W�/��!�Ta�>*�>rܵ=g��>4?�P:?��J>��о�A�̚X��Bt5�RA?���>���5������"0�so�Ln��h��=`���@�P>Q׌=��>�&�=�茽X�S���=gB>>I���=
4>��=5��=5�>f��=�=+j�i�C�=���LR��*�}9�.C����=z;ܽx���	㒾m������辍�,����>�{�>쿧��:5�$���������¾D�9�8����Y�%9��k��B������𼑎���B�_��g�#6�=;/�����Ǥ�Q�⾠ӣ>��>.&>�p<Ԅ�>�?�,?;�0>E�w>��j<]i�A*:>|��>�>dac>���>h��>���>��M�R�DW7�7��=�C ��j-<��]>��&>�AH=dۮ=��=��r=� )�7C=�
�=*�m������<>����4��fS><Ɖ�������:��rt�����=Gc?U���&U=
Ώ��Z��e�� �� &�=�b>^H!��Aڼa�I�nv�>V�>�8��\�l��!b>�~��J>b�����3�=��	�:x�=�Ȣ�n���R��W�/��!�Ta�>*�>rܵ=g��>4?�P:?��J>��о�A�̚X��Bt5�RA?���>���5������"0�so�Ln��h��=`���@�P>Q׌=��>�&�=�茽X�S���=gB>>I���=
4>��=5��=5�>f��=�=+j�i�C�=���LR��*�}9�.C����=z;ܽx���	㒾m������辍�,����>�{�>쿧��:5�$���������¾D�9�8����Y�%9��k��B������𼑎���B�_��g�#6�=;/�����Ǥ�Q�⾠ӣ>��>.&>�p<Ԅ�>�?�,?;�0>E�w>��j<]i�A*:>|��>�>dac>���>h��>���>��M�R�DW7�7��=�C ��j-<��]>��&>�AH=dۮ=��=��r=� )�7C=�
�=*�m������<>����4�(l)�c[㾠�1��/�+jM�B��=�A�G�&?<&�; ƾ���0~9���.d-��6�>���Z1��������ξ��G>
�6;z��]\��w�|���>ޘ=?)��y�=�� >�fI�Ν�=E�1�@1)��O�w��=���:C��=�v/>��*�	] ?��P?��C?��Q=��'��"�u�h�M�A��~�?~?�>�6>v5`>�$��B/�6=��h0���E��ּ�Ջ>�P�C�V>&�<��:��F=ʀ]=:��� 6J>��=�3>�ß>�>r�=�3�>G۶=���:����c�_���N����5�=��&����>��%����ƬB>�|b��E�<"��=y��<&�N=����o�:��)�Kz��!��^i�::ま�����܁�`��
ཱ�;����K���E�x�'�"�<ӹ���T�������¾F��z?Խ�>��!>���=��?��>��>�	=np�>  �>�/>rϙ<uP5>�F��WȻL	?X�?3�?w��>j���^/�Y�>�>b�)>�>>[��=�!=��
�g�.��e�<K�����=�ý�s�����\���0<�IǼ�fS><Ɖ�������:��rt�����=Gc?U���&U=
Ώ��Z��e�� �� &�=�b>^H!��Aڼa�I�nv�>V�>�8��\�l��!b>�~��J>b�����3�=��	�:x�=�Ȣ�n���R��W�/��!�Ta�>*�>rܵ=g��>4?�P:?��J>��о�A�̚X��Bt5�RA?���>���5������"0�so�Ln��h��=`���@�P>Q׌=��>�&�=�茽X�S���=gB>>I���=
4>��=5��=5�>f��=�=+j�i�C�=���LR��*�}9�.C����=z;ܽx���	㒾m������辍�,����>�{�>쿧��:5�$���������¾D�9�8����Y�%9��k��B������𼑎���B�_��g�#6�=;/�����Ǥ�Q�⾠ӣ>��>.&>�p<Ԅ�>�?�,?;�0>E�w>��j<]i�A*:>|��>�>dac>���>h��>���>��M�R�DW7�7��=�C ��j-<��]>��&>�AH=dۮ=��=��r=� )�7C=�
�=*�m������<>����4�W��>s¶�0��ب��1�V��=�3;���>#���	Ľ��y��?{�1���ߐ�2��h� ��M ��dǾ���>�F1>� ��˝�7>�=��<�>B1�>��轘|F�2]&�"���W�b��s�>�s�;f[��;�=i@S�R`׽�>LG�=�g?dAO?R?��=.��-��u�����g]>+�>>�x>G�8>��:�&�4�=Cٽ�Dk�:����o��<'�Y~�=E��=�[�=�.ѽv�����>�6B�<�I�;J�]>ʛH>�A�<6ב=\����^�L�>��a��M ���տ�a���-��.p�/�+�S '==�s��<�(�-�~	�=�!�3~�=Β>���=��>W!k>B%:>|��:��>ֿ�>���y8���*��é���0��>��~���<����I�[��zg�
���v�y���e���� �Y'��А�>T��>ܓ=%t�>��&?~�>w8�>nm�Fx ?�5ܻ��<�>��/>rR�>���>zY?[`�>��>��Z�l���՘=����[�=�`=����UZ[�ҕ5=i�>Q"����=�t;��#�RS>${�:�[>O�Z>�>b�>S�X���龒g��ʟ���=�[<> �P>����|��2���v�o >_N��	(��B���߸�%�>#��>Ab�>�:�CE�����5�K��=��k>bB>=�䢽D�м�N�=�Ƹ="� ��f���՜<Jw���ۘ���g=�F>���<&F!?yV?'B0?e�)>�M��B&�.�L�6K��Y��>/�>q)��UJJ����0Z�=��>҄F��
7��6!�\
��H=>��뻗C>aY�=/�>�m7�/�s=Z�!>T6=.�>#�=�ګ>�>M�>T�b>�h�>-�x��.P�6^�z;ƿ5v��L�ɾ�Fj��T��\h�8"��P�cT�3]����2�}�佟�D��.>�g
>�V>�=�7[;�¾�꽎��<�cQ�bh�����Xp�|l)>ѫE��鏽ä��2���0�9�Ǿ�M꽦q���ݾ����PD�G��>Td�>����><��>v8v>�\�>��>�p�>� ӽ�+��4��>$�8=���>mM�>��>"=�>�c>Z������6��� >D��<�>��؜$������<tS�<��/�Ά&�o%��9��u���<	a=��x=��>:t7>P���$�?N��O��Ĩ&��V�=o��>T�����>�1��V��$������4��!򓾌���K���w>-�>�w�=w����U�<�M=�/	���ν�;�=O�.=��>%�=re�<��&��T��d��]e��f=�+>�9�=.�<��/?PB?(W ?��>J��Yx%����f�<*���V�>�Z�����@����=���<�����ȾF��L����a�=�lv�o�9�2=<�n^�\�=�5���=E:r>��=�;=n��=���>Ppq>��ýPǩ��v��t�������"������虾ޱ�AǛ=���Ș1�JѾ��ʾ���<9��>0��>��C>�_�=^��;���=t>G�龘Z��Fc�q<o��r̾�ζ�����s%9n�:�H��eޛ�^��]�����R�Q��!�:���龗P���_�(��>�Ʒ>n�=�'>���>��>��?>��>b��>
E
=�`�=)�:>��o>���>�1�>�FP>�\�>�>�[�=6�^�%�~_>���=�!2=�4
>�;(>3��,W�=|f���jܽ:�8��J[=W%>{�K=��>�>��E����ގ>?�=c�ʾ^���ؾѰI���˽��?{w��ƌ��D���<���M���y���{�zz���Y�ap=P"�>�h�=�(1����<�ð=�8>8K�=F�G�p�>�헾٫�=L�f>xf��혩�pd��.s�:��W<��p>�>��"?t?g?�)'>%$�(��J����;DW.>r��>��`>}ʽ"dS������+���B���gӱ�A����=�=�=��>Ў>�i|��M���=g� �80>��>~� >�6=Kt	=�4>�1�=��=/�I>7
���1�a_y�J� ����4>�� ;*¾:<e=��\E��˾������<�Z�=g�n=�8>�{]>��/>=8-��;=�՘=����ꚾ�鄾��j�_�оF����4�E'<�t�0w��z޽+������!�,����Ƕ>��]>��Z=�>疊>�Y�>(��>�Լ�)/>��><��h<*1�>���=�~ʼw>�=4>��=Ɛ�=r/�3!��EM=Q~=<��=�h�=��0���ؽ�U}>I��<��8�����O��=��R>���=d�=�W(�N[�W��>s¶�0��ب��1�V��=�3;���>#���	Ľ��y��?{�1���ߐ�2��h� ��M ��dǾ���>�F1>� ��˝�7>�=��<�>B1�>��轘|F�2]&�"���W�b��s�>�s�;f[��;�=i@S�R`׽�>LG�=�g?dAO?R?��=.��-��u�����g]>+�>>�x>G�8>��:�&�4�=Cٽ�Dk�:����o��<'�Y~�=E��=�[�=�.ѽv�����>�6B�<�I�;J�]>ʛH>�A�<6ב=\����^�L�>��a��M ���տ�a���-��.p�/�+�S '==�s��<�(�-�~	�=�!�3~�=Β>���=��>W!k>B%:>|��:��>ֿ�>���y8���*��é���0��>��~���<����I�[��zg�
���v�y���e���� �Y'��А�>T��>ܓ=%t�>��&?~�>w8�>nm�Fx ?�5ܻ��<�>��/>rR�>���>zY?[`�>��>��Z�l���՘=����[�=�`=����UZ[�ҕ5=i�>Q"����=�t;��#�RS>${�:�[>O�Z>�>&�?�	 =`��+�˾����0�>��=��c>Yû����<+��>�!����j3�7?�R��=G�={��>iaD>�8K>&�u�Jy�����6kW>��6> �=����Z�#��5<Q��<��E=�
(��&��Z���>4�(>��>��<��{>��F?TU?��?��B>%�?�9�U���ྱm����B>3���r`Ͼ Ӿ��/����.����
��0�!_��Z�&>�fy:�hy���O��a6�Ƃ�D�F>B�>�פ<=�Q9ϧ=t+�>=�>�E�=Q����Y��Q:��0�fm��>�Ŀ�8�~F��(�Գ�d*��������*�4�HzW�
�>US�>X]B>a*�=�}@>�ɾ=��=��=sC,>~�u�	���I#龽��v:�BE�=@���%�<YD\���k�H�f����q�Ƚ�T8�@Cs�|�-�@'}�c�g>,�>$ր=V_�>	��>���>��>�D>w^�>�ν�'(=`}�>t�?��?�ʗ>���n�M�z\�N�#>T8S�A��X>h_�=��=q��=\C�|J�=R��<  >�{���&��<bC�<���Ǹ�=^G輬N=�r=5T�=��>�{	>{S�/���PH��4g>�sj>���> {�����L��<�pZ�1j¾���Gλ���=+͎��#�=�HG>a�>�i�=O�&��^ϽCEC>�R7>(p�=g'/�z�<J\�<:뢽H�;'���)����<<�>p�=5i�=�����>kv?s�B?׀?,��<b8��b�L$�h5�c8s>��w�6�����U�x����Ms��ݽN����L��Ol��$>�>���=�>�<�չ�Y �1T<p��=�\K�K��=Do��z�F>�=���=ZoS=������AW\�ğ�nҹ�A���@��Doe=+@@�lbo��9K�'�׽�t���)��貧�Ď=��0>��<>��==�=��=�w����>
��>���n��N���9��ƢO��g$>�(��w���H��?�s����,����v����K�7���P����'>Z�><2>���>l�<?�wn>]>pL�<d"�>pZ5=D=>m��>��>�?d\>c/�T �:�3=4����.��i�����=�>��Ҽ=���N�=N�$�t;@��Y=#�=-��=]���^�=AV��#��jns=��=%E+>��>�o��;��ks���8���>� r>i����Sʾ�i#>}a;>�{h��c���Ͼ��>"�>4�>8�>�vV>$�>U2=��s���$����=H��>$��>�� �u�׽���<��=�8�=S�h�4��`���6=6��=��=�p�=Cc�=�?gJ?yN?����mL�{q-��uȾ�g�=�
�=����^��'ս#��?���+7S�h����Z��g���_��4�d>��M�gh����>݌F��ӽ+%>���>��"��(�����=�qF>�Ԃ>�:p>i!�=Zg�.>��� �Ϝ�
Oǿ̘S�dϔ�"/�=�~��������ʾd�����D���7��@b��!>c�]>��=o�=�2q�oΆ�&�f������Sq�������I�����v��=�G� �<�+��H��m��Wͦ��Uv�(��`ި������i�L��>��>�L2�>\#�U?�?UԲ>5�>�P�>��O��(�</��>�P?�?��<�/�������8>ޡ>fE��DB���t>��S>2y=���<.H�<7`��V=���=�	�=�ײ��f����=��
=�7���
>�		><��=�>�>EbJ>���;J�ID��R�P�>4s?����r=C>��ᾐYǾxu޾2�>E�!=i�� Q>{5�����>S >tu1�rh��%�$�5>6�#>*ܚ<8k��LA�<bef=���`��<�H=��u�)���Y��=�#�@1=�>��/?�"I?pP?s��ÔA�?U�lv���>����>E�=�Ӿe���QھQhP���W��k�ݴ1���R�]�#>�/f=�B=�4�=$������Y��{��>Y�*�e��� >��=�*�=В>�">�Wܽ����i.����`%ڿC�����?�=� ����6�X�վ��<������e�-�d�}�
����>
��><=>�R>�=�=�Y�=Ƚ��eȽ+�2���Խ>y���N�����o�r%~�`����,����(�I{��}��{e������E�ʚ���a�b[�>�ٞ=�G ><��=v�?�F!?9�P>�u���>��j>�<�;Kh�>�r#?N,?RH��bｼ��=\�*=��=9��W�M��O>Į�=h�=�0�vE��8������=�Į=D�a=v�=S���bJ���$=��޼z�w=>|��=���>�K_>$�Vž��z>z��>u��>�:�%>ϐ���S�םN���Nh��1�C��x��w\�>��>'9d>���=@���s���=��>0��=�[�=pLǽ-B���e�˼zJ =}$�����<].C>��W> x�=
�=�^U>���>��.?��@?��E�����#��|��w�q��;V�ƫw=`]���݂����'���S���E�Vt���c�)�e����=�o�=M3b���=�_��;=V����>/�K����=$!I>�#a>/��>Hf�<#�V��P���[g����<�P��S�п=Ѿ &� ���m���K���2��ދ����=!=�r�һ�m�=�9k>�a>ᢎ=�N=H�_=����e���e=�Rq��0���� ��忾�}=���1�ѾR{=�:_���\��Jo�!�󥽓�/��~���
Ģ�?qp>B�O>Iē>M>��)?B��>8��� :>�EC?4�$�>���>;��>g�?2��>�u>���=�g���-�5�?�c���=>f�=*��=Tg��=��2 =�H�=�F>]u�=��������ս�<<⭬�-?�=���=+=f��>� ����i���Dؾ�	�����t�>���f�o=�ך>���<֧�����U���!��b���dվV��<`w�>�aH:˶�aؽ��D�Jd};��>�HI>��=
�'�焘>Uܧ=� ޼�q��GoJ���P�/�=@��>�l^>Ƒ�>���>��??��?5	о��*�D�žC���3^�W�>��j�5�>S�>El�����ӆ����c�r�Ľ�I�=�>���?>�U���{>Q<F>񼮽-忽��$�qp%�X눽FQ��i�˽��침.�>O��=޾3>�=�;�ǃ� V���̿�ĉ�}�%��c���Ǿ���4�/�K=�����r���I�Gfҽ��S>�<>���>�>�����<���r��*+�m����M���&��ܾ(=[i���!�U%����>!��=�Á�3h����G���V�������e�/Ҷ=Ҥ�>�8ӽ��_=�2?��?%�?�����(�>xE�ĢR�f��E��>�>�"�>2=>l�>u�>%��8��bN����>.<�8]:��=d�z=
ڕ����=��=�Jc�Tl^���ټ���=��=7�=�;�[r���+==>P)�����;��f��v�y���"5v>���\����a���B>ǋ�+t>�J�j�"$����"�EQ��"6�����>p_=��
=�U�=���u<+��>��=?�>=R�>�B'>���E�Y�r��]���G��B��>���>�>�z?�GR?�L?��)��6�h�Ǿ����C��[�>�u@�k�>.h�<��{�|���>���<�!�����\������,2!>Nt�>.��='sZ>�w�!$���j��,̚��j����4>��>b�A=|`p>���=Mse�e6a�2��7�0��`n!��1s�͂��/��2&��A�<�އ������
��d�=���>h�>�y>c/>4�<���륯>VY�>a0O�>��\����߾�Ӿ��	�86�?�;�i���fA�=e�w�.�x�KO����3�KO ��侾���>��f>ȱk=��8� "�>&?�Ȭ>��T>��@>or<��u>������!>C�I>=^�>�6�>I�u<�N}=}�&>WB�+����G=U� �b|��ʆ=:��=b�=i�t<~�>p>-= '=��<�w�=��8=B��=Ol>�����
=>�>�F���ɾ�Ѿ6*ľ�[���u���?-@��>���R�=�n>��;��侵�̼� ���q��W��#'�� �>3V��n3>�ڍ������K�r�(�6�Z>2,��`0>�ԗ>��>E�=����=2V�����>�>�;�>6r�>;60?юN?_���Nɾ�׾(���|�؂_>}�I��͎>�~>c�k�x"��>T���}��(>��d¼=�NG����>]E>[2>��=��$�<0���Gu��cZ���=>�T�>�5g<Y��>�k{>��&���3�ֿf��]�쾺'پ#�A��=�F�ޚ�������i��I��AĽ���=�f>�?t=��>��m>g�T�����>�L>%�����+�Q�=����,ö��ʅ=*c�������~��������3���tӽ8���o�m�%��_���D��>�}�= x:��E!?��@?���>�Mx��� ?Ɍ�hmi=/M���>:?���>���>��>UB\>]��0h��d9��A�e B��/=� �>���>������=��i�KR�<`���j�
��=���AqO��Sƽ�+x=�^A>���>���=�q���:���vо�j�������>ܼ��g����Ř=>>����q���?����̽7͏�㶽������>���;=��n����<*)�<�8��S�>�3����w�l�HP�r*ټT����r�!WH���eo�=�a>���>��
?\�?I@?{��.�P�L���N� ���7M@>�2[���>`�=�K���Ҝ�Q����d'=�<>��{���d>����"5>Z��>���< C�>�?�����;��置Ϲ=Z5l���=|�Y>��>dL�>�>�R������n���οi,Ӿs�J��E�=�~�>�� >�r׾�t��b�����C�q�Ǿ��ƼAF�>eX> ��>SC?�p>�ԍ���qʆ=�C+����)A���=���:lƽR&���P���}߽��=㊤;��u�2%G����n_�y����d����>�ן>��>4���3�>3q?e&�>P���==�8>��M>8������=�O�>+0�>���>(��<h����=�M>��}��_C�=i���@o�Ws�=T��>*� ���5�TI>�>G>���<�nz����=�F�=��I�1jL>f�=��n>f��>� ����i���Dؾ�	�����t�>���f�o=�ך>���<֧�����U���!��b���dվV��<`w�>�aH:˶�aؽ��D�Jd};��>�HI>��=
�'�焘>Uܧ=� ޼�q��GoJ���P�/�=@��>�l^>Ƒ�>���>��??��?5	о��*�D�žC���3^�W�>��j�5�>S�>El�����ӆ����c�r�Ľ�I�=�>���?>�U���{>Q<F>񼮽-忽��$�qp%�X눽FQ��i�˽��침.�>O��=޾3>�=�;�ǃ� V���̿�ĉ�}�%��c���Ǿ���4�/�K=�����r���I�Gfҽ��S>�<>���>�>�����<���r��*+�m����M���&��ܾ(=[i���!�U%����>!��=�Á�3h����G���V�������e�/Ҷ=Ҥ�>�8ӽ��_=�2?��?%�?�����(�>xE�ĢR�f��E��>�>�"�>2=>l�>u�>%��8��bN����>.<�8]:��=d�z=
ڕ����=��=�Jc�Tl^���ټ���=��=7�=�;�[r���+=_�=����A��iM"�-ľ�=H����h?	����"ɾ@\��s��^�v䢾�!Ҿz���Ȥ�����|¾Gw>��3>0,�=�#l�[&�i�=F��<R���E�	<ppd>����@�������!��f�	��X�<b��c�i}(�G/�=�H8?��!?�f�>����K0��KﾩR?�{o���=�G>�T콵��=$���;���o�ƾv����!�W7��(�ͽR�>7J> �[>2]�>�[�;r�\���Ž�&�AJ>o?�>��.=�L/>
�>m]�>,k)>�&�=qA4=i�=���׸��^]��	˾��۽���H�<`r>���=hX;��ླྀ!1>mH��<�9���>�=�<��u���>�y>�i�#�p��L���d���w��L�e�خ���;>�����䋾�2=�c�=�d�k�ེV���bB�7����Z�� ����>�f�=�W�>@��>��?<m�>�*�>���^�>���>���>Q��>�9?�D�>��>5.�>��?�(?R2?=2\=�5 ��ϽԹ�<�;���==s�>��S>�5>��G�yD�/� >F�+=C$����g.<�b��(>�>���>�pF>�Y�����0�z4|�H��-c?��= \�ۣ��7x�kܾO�f�q�6����?��T�
�]N���>�ˠ=f;�����d=>W��<�o�=�>�(������=S>�">:5=@堽³@�I2b;��=g�=�HI>��!??'��>�Z�>�
���+��I�ܶ��F>�:">%��=�_k=��-�D�E���r����: �����p���[>DTr>$Ɣ>o$K=P���q���Q�����8=��e> =�>�B�>$a">���>Zr�>�H=+oսbdľ��0�ʿK ���/�=Y>����|��W�p->>~��=Z�������$��˕=��8>�L�>J�U>��>L��>q�����&��$���.���(��F�Q����V@������>lT�*ɽ�T�����TU7�sO�����i��U����u���L�>�!:>!4@>�>��>{�?Q�P>7+��n$��=��>��>��>��E>��+>A}=�(�>��{>=�9=���wG�E�< ��=1%���>�̓>�x=��>6��=��P�,�����M�$�7�{�v�=���=�=���>�}�>���=�־������ƾ[�<Qk���>~�9�����yܾ� =�>K���s#��>�$@�O��"E���9w���>�Q�=�P��������=�	w>AjϽ�.��N�֤5=��=�w���`�V��H���X/=��}�ߖf�c!k�'�T>_1?�q?�j�>\뽘��ğ��}�1��?�,�#>a�;>��x>+��x�T�{��#��������u
=��>�k.>W8>>Q=�_����Ϙ�<�_z�,�[�1Zb���;>�gi>�ϼ�M>CU>�?>Opr����R���ÿ�s���q���o��,Gr�d�t>�3��V�,>�?���ʶ��c�^��P�>C^�>�(�>y�>�l�>�-?�\Ѿ�a4���Z��5����������t�b��=b%��^b�t���XE��KX��!������sy��Ɏq������T����>�=�>�ϋ>v9 ?��%?\�>����a6>	?��'��>ȑb>B�D>F�=�?`�Q��>n�>�u�>��=��bڭ���=04�=`oƼ
U�=��j>�io�ה�>��>u=�=�K@���!>�.>�:E�;�/�`=43�>��>�>��>$�7�~�i#�I�����L��>ŋ���M��!Ƕ=����ٔ���@��h��ψ=�/Ծ+���Y¾�gy>���=�\I�Ev��G�{>>�>���>%��<�P�+o�=�|O����=��w=�%��ṽ)X�<�f<>5=�=AHH=FvY>�e5?��Y?o:?�# ��QT��ɾ'.8�s�;���>-ў���<����a�+>��j��}�cZ˽�8پ��Ҿ̑�}I�=�?�=��>+9�>�-��&\�j�;�uo=>1)=g-�=�0�=9�=ʉ�>Kب>R&�����^<����N�șʿsJ��GĬ�$-�P��#7:>�.>�,�>�T�9���x�[=3H����>~��>�N?�k�>wJ�>x��>Q��D��X� �Sn������ ���p��jl�=�*e=�Q�� ��Z����?���
� r�VB�!i�aay�\�x��7�>�k�=+�0>� o>��'?g�3?�?��j�\U�=��>I(Q>
oq=��>�R�>-��=ԉ���L>�~�>B��>_r�M=���:�=���=B��*�=�ڱ=}��Me�=�7�+̘��3ܽ�z���6����1�T�>"�Y<Xf,�Z�>���>�pF>�Y�����0�z4|�H��-c?��= \�ۣ��7x�kܾO�f�q�6����?��T�
�]N���>�ˠ=f;�����d=>W��<�o�=�>�(������=S>�">:5=@堽³@�I2b;��=g�=�HI>��!??'��>�Z�>�
���+��I�ܶ��F>�:">%��=�_k=��-�D�E���r����: �����p���[>DTr>$Ɣ>o$K=P���q���Q�����8=��e> =�>�B�>$a">���>Zr�>�H=+oսbdľ��0�ʿK ���/�=Y>����|��W�p->>~��=Z�������$��˕=��8>�L�>J�U>��>L��>q�����&��$���.���(��F�Q����V@������>lT�*ɽ�T�����TU7�sO�����i��U����u���L�>�!:>!4@>�>��>{�?Q�P>7+��n$��=��>��>��>��E>��+>A}=�(�>��{>=�9=���wG�E�< ��=1%���>�̓>�x=��>6��=��P�,�����M�$�7�{�v�=���=�=���>���>�9=,ݾ�˽��K��^���@���?�k]���<���="Ev��zֽa���MEٽmk<���6���X�Nb�>�z$=��C�+L���S���XN>��Z\����ǩ>���Ehü��=1�f��^'d�#�Ǽ]�9�vg>��ּ��K?�)^?K�4?��>�k¾��ܾh�&���q<,ɩ��ǽ`��>t?�>�Ǌ=��#�6���o�,�+�
�@�= �	��&r>�O/>lk�>�x�=��5z��2'��'>i[H�6">m��=��z>�Q(>5I�>�s�>���>wn��-|����@����Ɩ��P/������z+�T�x�XG_�����S�{����5�"ʈ�󄐼���=�v��k+�VP>��������q�����Ͼ!\�������%��=��+�o�_�����6�=�1��?��*lY��n~�Xì�yB߽��.�"B�> �����C��s>3Z?��>���>.t���ɐ>�>_�&>g���/F��3�>I >�TP>e�>a��>���<������=	�v=R��=^�>��N>��^���h<����=L`��=l
�]�(=�2���=��On&>D��d��>v��=�O���h��,�/���彣�@>l&?�л=w����g�=�:���\<��>�轸F�5�+>ޥQ=��P>n�V>�����c�T�ҽ$)�y�v�a�L��'=��D>�e�l����TČ�a�����Z��>�p=ÚG>�]�<U/A?�(i?Q?��>�׾�k��H_��Y��Ԝ=��W��D=7O��j�Vy�Z������C ���a���޽���=�]>��=�L>8���㏽�\=/�=�)��>�<8j뼒;�>�H�>��>SQ�>ܯ��{�N�e������l;Ŀ����]*��Jf��!i��0E�<p���n��?������aL�p�޽/U4�v����%�>ց�=yS�<"��{��7�C��W���b�����ێ���n�E�=�c�s��9�4�,Zq��>;�T���������x��7��G����>��>��H�%��>j��>g�?i�4>�&4>ǭ�=�9�>�}�=Ч�=�i>@��>���>6��>�ϵ>ኙ>�m�=Ϻ����:�j#�=��>���=�&'>_�w>��۽�����]*�g �=s�5=h�Z�Ck�<��u=	�x=�A�<M��=�A�=*D�>K�=ֽ���ž���vW�=�95>��
?��(����/<V����Ԉ`�e��#k��2��!��dM�	1>P�=��ýFS���K��y>J�=Æi�%��������!�?{�=Om=$L�<��{�q���P|㼠)Ž.�d>K4�=��*?�td?���>��>=��W���|�r���!��=���=�?��U����\+�(�Ǿl�˾�P��v�.=���_{9><X�>d1�=q�>�xս,,����X�o҂>R=S������=�4>���=�S�>e3�>�3K>^�-=�f¾�,ٿ�뫿�ܾif��E�a[+;}�>{%��M���Β<ݑľ5K���"�R�!=s�t>�zZ>��;>�˕>��k��%��<۽����m����¾i�#�)LB��5>�ks�p�S��"��a�+��ƽ0�~�s�FAƽ��Y�j ��%e���>C��>��B�Y<?�"?�u�=�e��JQ>���>�Nx>�*!>X�/�>,��>��>�I�>��>Z��>������&�f���z=���>�6>�t5; !z>o$��F��=��>]Rd>�.W���*�c������
轤߻�q%>�B>1��>͞���i�X�\��I󾡦X>ŗh>���>��-9U���qv=i�=�V>��=hJ���P��o��3_t>��$>�ǒ>�)>@�ɽꛨ�T��
+��4�U�0>�}���]�=:�G�����?<6�	�ɽ�� �e��o�=H޽d�>"�o=ɢ8?�t?^j?�T%>��˾��!��4�����/��`�<��>�����5���	� �]��	V{���=�ӽ��=|z=hi>f� >����꺛=#��=o�>��k=�^���>��>�/�>�?�'�>Bx�=4�v��f���ٿ�ɩ�b���F�4���G�X��2�����=)��s=<n�3���Ⱦ���.�)�Q^�=4w>J
�=��W=j�T�iܽ�H~��l۽a�f����	TN��>!U����ƾI=½6��<�+ۼ\5�[J���K�7̀�Ը=~��y^?I=�>$�2��y����>�N�>He>�6>�%�>��=�	<�c�>�A�>�?Uv�>��=�	)�0��=��o��7��=B=�>U��=��>|���
�Y��M�=�%�>
�#>�6�:�U;&�3��P�EJ��NH?>�9�=̨�>pUD�A�l"�����_���U/��	?�>7;�.����2<�>���=>��<%Q�5M�ˌ�+ؕ>;�=XF�>s�x<���^����a}=�">s}�=E%u<@�J>}�~A��7���&�������<��Q=RJ�=K��= q=}�]?x?��a?�2|="�⾺����D�u��=�[=�Ȧ�-9��sܧ�"�"��v.�X�>�]z�q�N�t����Ӿ�=�"�= t�>*@>~�Q�I����E�=d�>Jⱽ2Xz>D>ҩ�>;xL>Eߨ>��<>��l�ҽG�����G�������%��i=�IO���R��q��Y�f�e�=N�z�}���R�-7�=�F�=��>�Z>jSw=�u���i�i��<�y�}����-�X��唾W2W=c�&�$_��b�����)����ʽ�U��X��iU0�Nî�����I�>#����D���>�ۊ�>�>+?��?�l>�=�y>�?s>����XZN>�A�>!�	?WV%?~w�>n���Լ�]2��7�9�=���=�r��F��=��=;7�o.I��?k��d��
�&=�&U�Sk�<;P��	��
=}��;��=��>��>\_t�	ڠ�� ���V��`H>9>DG���r�Z\��L�<�<`��� ��Jr;�Aa>t�v<�d�qqž��>�FL>?�������X)>���=����?׽� ������%����Q:���ͽ�Ǿ�"���Q���(��?�=��w>N:[?��u?��#?��{=���q.�	;q���i=`>y?6�̾�@>6q=�Oξ]yX��X�v{�}��=���Rd��,/>��3>Gt�=�M�<�7��A`=:�L>�(C>ө>���=�'�>���=-��>�J�>>��P>����)����ɿ��:�AD���׾9�(=�U�=�n>r
���~�> �S�+�I3G>6�T>�Φ>��;B�=l>z%�>1_��ޱ�7[/�1߱����޾W�G��b>BV�X(y�iG����;=�0��l��b���(��͙��W�t����ڭ>�݈='�e�f>��?�*>�?#>`Ў>.el>�܉�^8N�e%�>ZAw��Ss>ZnX=�>��D>�T�>䪂=��J��Ѕ��b�<7�3>3:�=�=�8>!�м��=2�=���=��<%q����>��>gXw��*=͚�<Ya�>�'�>1=�<�����4˾c+�Ds����0>Q~>���w?�=���
N��>��ⴝ�M43��0�����h��kݟ���(>\>FA�<�m��{;=���=ty�<H$�	�ͽMG�=ʃ ���U�� ��e</��7⢽Kf�Az=�{[L=l\�=�J?�	P?׋!?1m|=���R�U��[�_�4���..>��\�<�)r����#�r��+���$��U]�2=k=��J��#z=��>�߻��p=c��=F�D>�/'��U�>0a>�>�.>h�>���>\�>G�=;�&�^����տ���~�*�G�ռ�`�=!���[�>RNŽ��ҽ9G��&l���>�bG=豶>���=�D>*[<�B�>��?�w����=+2�=�䊾뇗�����k>Fž�ֽx�
�'��>z��k���e/�������#r8�ā��,�>��>{�D�q�a>q� ?B�>���>%�>���>s��<iգ>[�2>�i8>�r�>I�y>�	?	L?I?��1>d*��5���1����!���<��M=VQ(����=�B=d�=v.ܽ���;3d�=!ѷ�v���݃�=�q>��>�1�>�E)>`��fU������p����n�>�HžP�n=����<����.����Y=�g��O־��y�������>ǅ>�Sݽ������=J�b>�o�s��
�>��VN��0���T�����<�P������_u��>�g��d�>��-?HE?��?H>�bE�:p��f�b��
��9V��B>:+�qi�>�:|>�O뾋���
����8����&�4�H2>��1>E�6>���=�����=����>J]���>?�>��+>;�>�`�=���=�{>3%=��=����ҿ����=^�X�B<q�2<��'>Ɠ�><�L��?����A���;*";����>f�>k66>�Χ>��>���{I*�gⅾB/M<�6����ݾ��3��d\>��9/?>S����ό=��x�,�m���>"+d����Ss�RIQ�pۿ>��e>�=t>?#>C͢>�$�>r��>�^>�p�>Q�S=���>��>��=�I�=�_�=��>��?zh?̠�>���g
�W�>!l>������=.u�=A�f<Vd�="l�=�t=)�н�Y4=��=<A+>��$=�߸=� ���>F��>���=���"z��C"��⫾�t}>���>`	[��e=�eʾ��>Jz澿�v�/$=�������.�D���~�>���=Nљ=��n���=��@>����ҽ.}y�l�:>;B`�%�)�Ll`��C�=Q�_�<-N=�z��C�k���^:���>��Q?z�2?=�?�>I�<�%�].D�|`�4��Z{>�[�U�>�>$	ǾQ��'�J�����Z=�63���=">�ˢ>�Zc<�m��$#>�b9����=!����r�>�ݼ={P�>�R>>�>�>�>F=�7R>���=0��4ܿb�K���%�)0���Ǽ�=�vD>���1��z��r���)��`>1G`>���<�&B>��}>�va>:�j�Z��/쌾�P�� ���Y�������=��ܽ ���v��T�=��>��s�b0w��*o���,���U�(�0�>��>��>H
�>��?��>�+'=Ż�=m?}�T>�X,>��>Y>�T�ݥ�=�7%?�R�>��>bۍ=���CŽ�^�����=CW�<֮>��^=E�S>kb��fN�P_�d	���	�q8��ī=P3>r0@>�E�='�>�{=|}��Ͽ��R�|��@�����>�3,��$�8d�	����姾_�4�ڑ��k�R�Id�0��K���2v�>}M�>���=��L���;�����Lg����4ڽ��̽z"۽4qY�6�������uN��?#u��o�=]��=W!�>��K?��U?�>�u�����<���U�f	�=����'��=��M� ��>���<%��C`���:�_�����=J����)��%E�7u>(,�>�ܱ=9�>@�>�|]��[g>�Jm>f��>Η�>�3�>�N?2�>N4�>5g�<����Z�z�¿J׾�\��~���4r��<�>y�>B�����?e��n C>��=+�V�+�a>"��=�[=�d>GI>|Ԍ���ĽqH��L����þ+i�u7i��w>8�|�B�彆萾�a����5���޽�	��8Bf�l��z`��#ƽ�K�>�0>t�G�2�\<n��>��>┢>��=��>�b�=�n�>*Oi=ɽty�>ǣ�>��?,�?i)?ߚ�=��,��5��\�v=�X���+�2>�~=/�=/�:>B ＇^!=;���c�<!�˽���9�ѹ=���=1��=� �=p��>N`~�{�߾�T��6�e�<!q�>�7�>��I=A�]���¾j�����`w�2H��R�y�e���<S�]B�=G�=gֽW��<w�a��>�,I�`�����������=�Ⱥ�<E=��$:��<������ξ�����>�k>)�v�- �?���?9�i?�?ՐL��`f�F�}����U�	�H�,>���>#\&?P�>��<�n�� �о5�1��,;A.��?̕=\�>f�>.�>9�;N�J�-EC=K�=я(=0�b>[F*�hqp<lJ/>���>��>�x�>�~ ���`�ֲ�
������-��Ѿ��>�>�U<����v<�a]��_��8��c��������t>�c>c��=�6>?�
u"?D��=`�ӁW�*U/��D�='B⽞�	>(�=�H�}U`��۽�c�aK��$� ��~{���K��)���M~�>Բ���Yd�"�S�d�=6*�>���>���>3$�>4�>��c> D�:���N��=q�>^3�>���>6��>Ɵ�e��M�ʼ���=f)�<�&q=��O=X)D>���=��=ׅ��aF��4�=��=PT���S=E�~=�[:�=�|�=k��>�8.=����w*_��&m�bI�>�$�>,0>O�=\
V� (��=�,�=��]ƾ�4�"�!��Ҳ>i��>UyH>��ŽFe>1��;'C�=C�M��`��R�Ǿ6�x��z>�3=�>~�����yݽ:U�ɻ�Qa>���=:*��SV?�P�?��x?V�>��+�m~����S��0�z�>��=�ӣ>�^k>,b`=�þ�n徥���wܾ���;�����=w�>�n�=&U>�O���;=uψ>����C���<Af�=ճR>�Y>�j�>�l�>{�i<�W��j�6�ÿ"�����4��(�Jq�=�{�'�:�0�F>~�$�r�>P�ھ����Sl��IR=}Ka���A>��>j�w��}>�Љ=�`�_`��l-˽�b��X{Խ�޽��>v�Y���$;� � -��f�(�h���T��On�j;�)�z�-Ѝ�\�>��>�Jݽ7���D|彻>Q��>7M�>ݘ�>0�~�ꭋ>���+�r��ǀ���	?���>)�U>5��<4�ݾ'�޽�Ğ=�7<�*b�J��<�k{=\�e=���<��>�Pн�I&�h�ѽ`���Ħ���ٽ?�>ҙ=Y*F>���>ʵg�%����z�������>���>@?Y>�/G�x"��=  >X�+>�z >��¾O�۾\s��HjV�8n?諹>��g>���OV>�.�=�H�;����`D�����P�<ߋ>�iý��>مQ<�m��Dž��g��A=���=~JἃGT�b��?}l�?��m?��?�B�+�>�Ƽv��au�&$�=
�2>�z�>���>��=���"9�������� �5>���=,|ͻ�Ud>C�$>����-���J�>L�=2b&���2>��=�&�>r}�>�4�>�إ>�Є>�|[��ˤ�&Lڿ����#��ؾ���؀,�oj��RNt=��=����4�e�o���ƪ��˩e��b�=�?v=Q�>��s>�C&� o������ DžY������Q��.<`>-��l�a�$�&��ێ<�o��ys�������Ǿj���s=)M��l�>LY���������\��>��>{�P>�l�>}[U>ɥ�>��J��p���n�G>P��>��?��u>��&6���"���l�<�;{=�N��%M�=�K;>�D3>ˀ=}b��}�<���=�ɽ*o�<I���M�+���=��׽I��;��>FT�>$��=��k�\�]� ݍ�8+��6�T>3��> �>�YԻ����������z�Ž�PF=�%W��ాP�1=�#1>�5�>����� ���>�2�'�|��*>�� =, �wr&��O!��X4>$�<&B��:��@�d��j>Q�=�R�<�@>�C?�{�?�9,?��>j�^���"�jX�L���_��>2��;1�>g�>���=�ɼ�8���0��,s׾�� >�߭�p��>7j?=W,>T >F����Ҡ���=܈�=��>eN>�4= ��>���>��d>NG>��D�L`��)�޿HC���#�T"�h/H>|��x	=s!*��b�<�O���q���9ľϜ��f�=g��������>�>̽�i�>�(����?���0�$���O����Z��_<v��;�<Phܼ���&�./��t�.��I���!��##����=H#�}��>@�>���K���XP�c�?Q��=�Q�>ؘ��j��:�>��u>�=�=P�Q�ũ>��-?��>uIo>�aɾj����<W�9>��_�=.�=��K> !>^�����[=�Nx�l���L����Ľ/��=HD�=s=Рս������=���>y9����.��V�S�G�Р>��u>|?���ʹ'<%�¾2(N�ƗϾ�熾V�>��b=����a�k�����=�!P>o,R>@4��)2��l��_p>!٢=���=2�$=�L�Ջý���=b-�=�;�=#��=����,��	���^׻�_O?�.�?ڥp?2�0?�QF������M�@���C��m%>qΊ>���>�8>m��	�����(��,=(���a�����<�O�>�e�>�0���{�������=mpa;�V�>o��<�l���N<��f>��ϻ�>1>b�.=!`�\3��º���������e��=]<��
�0J��P����P�eT1�ʑ��M_���w� 0p=���z��<u�>���>���>I5�ľ;��U)���_����b�A>����4��=dX��x �8{�� �_�D"�ӣ���W*�N^�<��]�Ss?wLZ>��7y�ij;5f?��>�K�>��>~��>��>a_�=���=��I><�<����>���>�ڷ>�bE>�����iսvX�<o-����=�qE=���=��/�(5���ٴ�����B�=�`�=��<�����p+=T�U���}�(�>\�:m2��=�7}վ�&��w��J>>
��>�ڭ���g.���� �_�u�������G=�������5�nrJ����>�:T>�����V �<�2�҈Z=�hn;�)�����=#v��o�� <3�i��>S��'�������$�p=O����>L�?��?I?oj->-c�x0�Q#�V\��.0@>�R�>p�c>:,l>�}���4����G���j���Z=02>�.�=Xh>1[=�/�>kn�=��7>a��4>6��<��>�4�=k͗=�d�=>;�>�U�>q�>�q�s�h���� ۧ�Pw���4׾�X��2>O�au���T*�Fr��.���R��`42���>��>>�K>�q�>Pv*=�P>�N>�������!V�Sf��^�-��(⾣�p��4>f�l�K�׾�UҾ�`d�ZV��Y�Y���=�{��ԓ�����'Y���M�>*T>�>Up>���>��>�\o>���=9t�>M>Sl>r·>�����s�{>��>��	?f�>��=�1����:�>-��=�C	��R>��=��A=<�_>I@�=�y�=�]�=�=�<�1;�J��.,�=�J>݄�>�>���=t!�,�(��Ra���V�V�K=Դ�>2���^�A5־ήȾ� >=���|���N�$�D�` ��tJI<���>[��>V����b�� >i���w�=��$>~��OX>J�K� E=� >����J��+��7i7>Qga=�I�	�>?��>��%?�?�S>
ʶ��55�\���:� ��"�>0|@�I�>��&>1���Yeݾ6|��Ϫ�*z��!���i;�uOO=	��>>}h� O�>�I;<\�^�y�	�Rg>}��<���>��$>7��=��]>��>�B�>[��=f��kW���u �	Ȕ��־����k_�)���8��;��6��'���`8��SV�oZD�#M>��Q>Б�=n!�m��滬�窳��U���dI��(۾�t9��q��-��4C>��1�C����ξ,W��2P�%�"�|M%>��"�/�� &��޾v�>��6>6ܪ=�V5=�L�>:-�>�_�>�ΐ=�j>1�����>�b.>0%Խv ,>F�H>�;�>u�>mXA>T�<cʼ��-��6����>[��<��9>NB>|Nս�*�=센e9�8�:JvM�W��i�9��O�;�oM<�؀>��>`Z�>�>�־��D�~��߽��_>{��>�$���ɼ0އ�)�u��B���9��K��d[]�,����/���t9�]�>ٵ�>{���]~w��n���0�Eļ=��=�#�;�I����=酄=7N��OU%��&��E�_�<��&�@��=��>��?n��>`י>j>���� �K�g��@G^<�r=��E��`=��b�ʄ���@�Hv��^	޾��O�r�+�I��hf�>�E�>Q��>\G���ֽ��k~!<cS���E>Fy>Z�>��I<�`q>��>:ڑ>�-z=����f�˿�_����׽��X)>�W`��k#����g����Y�=�T��P�>lY�=fD�>��>�+�>��>��.����_��5~������֮��yD����=�2J���y�&��l�-�t���5'ս�W�=y8�:��'���������>�>z>g�<>CN>9��>�_~>?[#>�^=�e�>e�J=���>�z}>�>�[.>	�>��r>���>e�p>�琼���=6���?>�]2�ÐŽ˳�>*,�=�����N>�>S)��bh��%>�Q)>�c��������= >`Z�>�>�־��D�~��߽��_>{��>�$���ɼ0އ�)�u��B���9��K��d[]�,����/���t9�]�>ٵ�>{���]~w��n���0�Eļ=��=�#�;�I����=酄=7N��OU%��&��E�_�<��&�@��=��>��?n��>`י>j>���� �K�g��@G^<�r=��E��`=��b�ʄ���@�Hv��^	޾��O�r�+�I��hf�>�E�>Q��>\G���ֽ��k~!<cS���E>Fy>Z�>��I<�`q>��>:ڑ>�-z=����f�˿�_����׽��X)>�W`��k#����g����Y�=�T��P�>lY�=fD�>��>�+�>��>��.����_��5~������֮��yD����=�2J���y�&��l�-�t���5'ս�W�=y8�:��'���������>�>z>g�<>CN>9��>�_~>?[#>�^=�e�>e�J=���>�z}>�>�[.>	�>��r>���>e�p>�琼���=6���?>�]2�ÐŽ˳�>*,�=�����N>�>S)��bh��%>�Q)>�c��������= >`Z�>�>�־��D�~��߽��_>{��>�$���ɼ0އ�)�u��B���9��K��d[]�,����/���t9�]�>ٵ�>{���]~w��n���0�Eļ=��=�#�;�I����=酄=7N��OU%��&��E�_�<��&�@��=��>��?n��>`י>j>���� �K�g��@G^<�r=��E��`=��b�ʄ���@�Hv��^	޾��O�r�+�I��hf�>�E�>Q��>\G���ֽ��k~!<cS���E>Fy>Z�>��I<�`q>��>:ڑ>�-z=����f�˿�_����׽��X)>�W`��k#����g����Y�=�T��P�>lY�=fD�>��>�+�>��>��.����_��5~������֮��yD����=�2J���y�&��l�-�t���5'ս�W�=y8�:��'���������>�>z>g�<>CN>9��>�_~>?[#>�^=�e�>e�J=���>�z}>�>�[.>	�>��r>���>e�p>�琼���=6���?>�]2�ÐŽ˳�>*,�=�����N>�>S)��bh��%>�Q)>�c��������= >��'��Qӽ���.��L��_��2K�=�ӻ>>������l��=�W=-�����f�4��=��v>��>fT>�S�>�|	?^�mоS⽯���`e�=�fN>�M>��Y<���]��C���4>��>�T�=@Ju���z����1u>��>�?D?��>�������羄f��xj�s�W=�tͽ&�>��>n�>�d��0���B�<E��¾�GJ<��A���>�u#>;>K�<7��B����")<�*>7	�=J&�=�>�;��k=5�=�J�9���<���=j]��n���r��G�⾷=���.< �����>�v!��a��I���W>�>�<�{�1�ҽa�Q�"c>YW>�AD>9�>�c&�ﱾ��_�=C���ɾZ����Ӿ*��=|�*�Ϳ����0�M�>�)=:x��w������4�P9@���>�G?��K>�	_>��>�l�>��,?�׿=u\K={�
?��=`8.���7��V�>K��>Q1�>.#>nT<�R��r�x�Q���Y��:5�=�{�>f�.>�Y>��)>��0[���k�<��=>��=MJ�=�\(�&���D9=P�=� /=�+>���=g#>yV�p�&�辟����=~��>_v��fCu�E��AS�>%�]p�v�
�BY��-1> ]�>��B>�k>��(>a�����[��Џ=�=S�!L�=��>V؝=�*:t�̽����=:�=<8b>�5���#��
�,>���=P��>�?>�g?w@$?x<ؾ'��4p
��2�ޠ��X;�>
��>%t-=X�?�R4=8'�<�h�Z�\[�Z�x�ۼ��\,�>��6>c<6>
d=��~S�3�F�)0>{��C?=�+>�i�=��>�O>�.C>>F=�<[��ñ��T�l�ֿ�c��n��cZ�><�;>D��~����Lz��򇾏��>ұ?��}���Š>�Rr>x�F>��'�E�T���/�/�+��>e=nM���^�ѮҾQG��Aō�ʙ�tާ�������!�Lǳ�]�c�Q;�i����K���3��M��8z��C�>p�p>F�^> >�f�>{m?}1�>y2>���>��:>�FT�:�o��^�>���>䟰>�I^=�>��=T�T=�޽�﴾�/7>$v>�'=�C�>�+�=���[l߼�:>ל0=
�<{�<Ak������=x��=|�J<E�z>��'��Qӽ���.��L��_��2K�=�ӻ>>������l��=�W=-�����f�4��=��v>��>fT>�S�>�|	?^�mоS⽯���`e�=�fN>�M>��Y<���]��C���4>��>�T�=@Ju���z����1u>��>�?D?��>�������羄f��xj�s�W=�tͽ&�>��>n�>�d��0���B�<E��¾�GJ<��A���>�u#>;>K�<7��B����")<�*>7	�=J&�=�>�;��k=5�=�J�9���<���=j]��n���r��G�⾷=���.< �����>�v!��a��I���W>�>�<�{�1�ҽa�Q�"c>YW>�AD>9�>�c&�ﱾ��_�=C���ɾZ����Ӿ*��=|�*�Ϳ����0�M�>�)=:x��w������4�P9@���>�G?��K>�	_>��>�l�>��,?�׿=u\K={�
?��=`8.���7��V�>K��>Q1�>.#>nT<�R��r�x�Q���Y��:5�=�{�>f�.>�Y>��)>��0[���k�<��=>��=MJ�=�\(�&���D9=P�=� /=�+>S�>�r�>�(Ͼ�U� M���߾�"=�?��C�����έԾ� ���7��s�)=i���𐳾2:��6^�=eL�=k��>7�=>��U�]L��	��=q�y�-�;���=Y��=6]=��?�8i����'��ʙ�c�����<���=�P=;���n�>b�>R,j?11P?@����RQ��4�y&B�>����*>�=>�>�>��>�^����������/þI�Z�����8�=D�>'M>$�/=�69���3�:E
����<Ϊ`��	m=�l�=��Z>.X>RU>��$>��̽ɮ �G���]���5ƿ��?�N��d>=ʂ�w�=1�=}����y��ͩ5>�Ͻc)-����>�|H>��=�4��~F=C�*��m6�P� ="j�O��!_��9߾b`���`#>��U�ڝ���y���=��g�.#�_���߽]���6u%�������>"E#=�w>��>�ݻ>`x�>�Q�>HS����'>N�>m�'>��c=%>��=/`^>�1�>�?	Z@>���=��뽄�c���)>Ǯ�=4�*���Q>Ȗ=>_)����k9�=5�L=���ρ<�(m�����ʁ��Q�=eH�='V>��'��Qӽ���.��L��_��2K�=�ӻ>>������l��=�W=-�����f�4��=��v>��>fT>�S�>�|	?^�mоS⽯���`e�=�fN>�M>��Y<���]��C���4>��>�T�=@Ju���z����1u>��>�?D?��>�������羄f��xj�s�W=�tͽ&�>��>n�>�d��0���B�<E��¾�GJ<��A���>�u#>;>K�<7��B����")<�*>7	�=J&�=�>�;��k=5�=�J�9���<���=j]��n���r��G�⾷=���.< �����>�v!��a��I���W>�>�<�{�1�ҽa�Q�"c>YW>�AD>9�>�c&�ﱾ��_�=C���ɾZ����Ӿ*��=|�*�Ϳ����0�M�>�)=:x��w������4�P9@���>�G?��K>�	_>��>�l�>��,?�׿=u\K={�
?��=`8.���7��V�>K��>Q1�>.#>nT<�R��r�x�Q���Y��:5�=�{�>f�.>�Y>��)>��0[���k�<��=>��=MJ�=�\(�&���D9=P�=� /=�+>ru�>{���/�*��ˠ�lG���*��d�=X����>�g�<�s��	t��Z���Ӿ2��<_�>�=�>��->`!�>4��=�&��]T��_�<y��=������<�#>��x>i���ь�?0�=�i���G��µ<c��=�e>(j�=. ����X?��>��>��b>k�M��BE��¾@5��]��c�>���<��=$�SLھ�W4��x/���뾓�=9��+��=8i>NH�=��>!�A�G<�x�<(����X�����=%�r>���!uk>�NI>��=]��`g����a��f�����������'���*��蚾;��XЇ>!"�M�C�x��j�>������<Q�=b�O�W�ȽY�x����;Bf��`���ï��1u�E1�:̾i�j��z>ãc��4��
���=*�t$v�#Ğ�*ٙ����w,��_����/->������<�o�<�MI>��,?K�0?W�;�>>z)���a�=��>��?,2?�j*?�
�>α�=��8���,���½���^�>� n>��>N=��(>�i�ЯU�j����>���<:=h6=�߳=��Ӽ`�Լ|4c=S�>Ӎ�>�A����־�}�w���cν��>:}>�N��j��=��<>���>��+	��v��$�R��9�>Z��>�UW>@ot>%��<�<�)�O1�Hh>�+�Yp�}Fؼ�Q7�ω�<��`�&i��� L���ڤ�%�(=�g�=���=��>S�)?�@?Ɗ�>��f='��R,F���.>��(���P>o�`>� ?���o��pþ��5����7�=Sd佻�`>"��d7���->���3(:"�D>�j>�>�<j$��E�=�C>�%�>])�>.47=��>x�B�����E��m촿�_}�����B�Ѹ:=�` �9�!�\���G�������־�B�WG�=0&�=�.�=�߂<�q���[d���u=�R�=�`�#�_� �+�H��0�x [>���=�5�<�|<�Ur�=oy�h.	�
�<�Ar=�g��A޽p&��3N>�-�>�̎��e���>�>�>��2>6>U(c=�i���y���o>��?%�?���>h��=�wQ�����@�O��j��G>Z�>?�6>�Ы=�[0>�%f����>��=<��=�=�����=T�;䁣�xơ=�*>l��>2x��+��/8%<_X����x�?�-�V�>�:�w>K��=�9��q)��-=����/@���z>��
?f�>��0>���=�X�=��/��a���|ɺ��D�`�� ��O�Խ�b�=Fq���5�"/��`��5���Dor�M�M=�L>Hp�=�J[?MQ?:�?�bE>��~a�IZ&���=%�ۜ�>��<g��>0�i���MJA��!A��rr�fX�>���c��=E�𺨁>�'4>h���&��=oV>�F�=� ����ɍ<�0>ׅ�>
��>�C�>�=g<"�� ��9�����������#��6��ف��S�;�o�;Ἃ�kP�=�Y��������a��<X�G>*��=p�=T�����}�C�>�=>y�����G�WG�b�����*<>(����>����Z����^����3�=u��K�rX\�ު���Ne>_��<3D/�ٯT�����?B ?p=�=�s?�a��2{��]=���>~?(?}��>��^>��w*���޽�?O���%<O��=>^�=1>���=�ܽb��=��=FM=v��=�;e=��b�����hhK��'c<h�==) >]	�>4'��)%��������<n;���>N�þ"Z�>6��=ח9�/.4��p����復+����<��@>\�@>�Ps>S��=�	O���:��M����=� �g6��2!=�%��w=��<�W�����>�����g���x��s�>�̗>0�(>�\@?��?��>��>4�@�2a����v<�:����x>�繼[>ړe�󱻾�7���F��緾��H>ӕ,�^��=��*�1�Z=��w>ҽso���<"e�8_ǽ�����ܸ=t�>D�T><T�>dU~>��=!
�ξ����(	���� �%��LT��&�t����)R>{����HY=�[�)H��}�:��=�w>�9 >̃P<w�
>�+<=�(>��V>�V�O{l�e�ž��3�7�-��M�=Jv޽JWO>��@� �K�>L�;��s��	:��2��\@�<1Ze������!>\�\:���=@S�=.��>H�!?��?�&�Ϧ>b�S���=�8 9>� �=�?%�?M,-?a��>����0��8�G���u�R"&>�g`>�Q<x}\<��>>�1�Ф<✺i��=�{���#>�T�=�'�- ���U��
=���=ru�>{���/�*��ˠ�lG���*��d�=X����>�g�<�s��	t��Z���Ӿ2��<_�>�=�>��->`!�>4��=�&��]T��_�<y��=������<�#>��x>i���ь�?0�=�i���G��µ<c��=�e>(j�=. ����X?��>��>��b>k�M��BE��¾@5��]��c�>���<��=$�SLھ�W4��x/���뾓�=9��+��=8i>NH�=��>!�A�G<�x�<(����X�����=%�r>���!uk>�NI>��=]��`g����a��f�����������'���*��蚾;��XЇ>!"�M�C�x��j�>������<Q�=b�O�W�ȽY�x����;Bf��`���ï��1u�E1�:̾i�j��z>ãc��4��
���=*�t$v�#Ğ�*ٙ����w,��_����/->������<�o�<�MI>��,?K�0?W�;�>>z)���a�=��>��?,2?�j*?�
�>α�=��8���,���½���^�>� n>��>N=��(>�i�ЯU�j����>���<:=h6=�߳=��Ӽ`�Լ|4c=S�>Ė>����󬃾�z�� ����\��?�<�Mp> J����2�Dt8���E��o��K��ME������ٸt>�>�̕=Ypp>���(!��# �>	>�<�x�=]:m=j�Խ����
�Q=�[d=�J��0σ��֛�9b8��)Y�r�E�1m>'Qz>�Q>)�*?�$B?WA?���>�E!����>)�{�->y�=��=���>tډ�������=��/��s��h��.Ne�ǈ�<Z�>�?T���1>+�o>n7�=�%��4�<��L>��6�D�R=��=�9>pA�>?u���Nr=���=ҝ=�Р����ÿ�_���zپ�k��F펾��8�?%�/Rپ	��r=�6�������NҒ<�Ϋ=�3�=0	;>k�=i���qf�A�E�8J6�hx��-���zs�uZ�:�=w9��A���Å�/_��ڊ�٫=`��ǎo�ʉG�T]i��#��u�>z�c>~�ν�h��a>���>z@�>�hN>�">�>��>AG>�h�>���>7�$>��=bO��
ܽ3��=6��o/y=;�>�A����+��QL=#^O=��>�P�=^��<V<�̢�����ڶ_>bo>C�>�7����ڽ��c>����!��C'�S|�w����,>�G�>����>Z���d�}C5�����ZpV>���>�qJ>"਼��a>n��<�ے=�:e>�ν1�>��z=1�8���<3�=B(>��ͼh�8>רl��t���*��S���k�=�� >�0>q�&?ǟ ?w�?�bμCB�Rod���Ƕ7��j����>�=�>��=>��f�o�Լ羌.�$�о���'���n >��=PZ��w>�����:�+=7�?I{���H�=7]w>�������>Z"�=|	>-
>	�d�M� �����q����]޾ӥ!�ˡ2������\��"�`�b�u�Ì���R�`,���o>�5�=�0=<����J�ߘ��X�����=���������ᾌ�`�f����3��K����9����^�ƾpИ���U�ʗ���Sh���� ���3��CX>8s=
F{>4�><�?�Z?R�?C�>Ɠ?��ǽ��)>H�>�Q"?f�)?���>ӄ�=z�=ӏ->�&2>��p�!;���<�<�Fj=���=�$>W??=#�������`���b��8�d�(��g�=��%=�C�;K��=N=r��>Q-��A:¾K[�])�֋,>h��=>�=�v�=���=�����|�쾠��u���~&�>ŝ�>J�>�#`=p�>���=�]�=���=A�=�Dʽd��=Mk5�s;2�,=��+>�R���<>}����,L_��U*��T>'��=�v=jc?�Ձ?�j?���>�b�80�6��.�K�\��=�/0��s>"��>;<�mD>ǝ۾�����K�̾�\;�22!>$�m<��ܽ��=���=8Ο��?���>#��;M��=���>/G>/�->��>��&�=�����j�!�@u��`e�v������c_=��#>��I�H�&�����&j������=�>j�;K=Ww��=(�������ol�}�[�eq��Zp���ξ���̄�z�g�1SI=��9CUc�9�F.�7����8���Ys������v��]?��-�M��s=؛>�?���>VΧ>�P�=Ǭ_��z�>yV>L�~>Z� ?��l����<7��>�b�>����:
��Q�=�=>�;�<N��=�^�=U��<�{?=Ӊ��g#�Q�ɽ�-%�F��=���=G�=;�S>#&���=��c>����!��C'�S|�w����,>�G�>����>Z���d�}C5�����ZpV>���>�qJ>"਼��a>n��<�ے=�:e>�ν1�>��z=1�8���<3�=B(>��ͼh�8>רl��t���*��S���k�=�� >�0>q�&?ǟ ?w�?�bμCB�Rod���Ƕ7��j����>�=�>��=>��f�o�Լ羌.�$�о���'���n >��=PZ��w>�����:�+=7�?I{���H�=7]w>�������>Z"�=|	>-
>	�d�M� �����q����]޾ӥ!�ˡ2������\��"�`�b�u�Ì���R�`,���o>�5�=�0=<����J�ߘ��X�����=���������ᾌ�`�f����3��K����9����^�ƾpИ���U�ʗ���Sh���� ���3��CX>8s=
F{>4�><�?�Z?R�?C�>Ɠ?��ǽ��)>H�>�Q"?f�)?���>ӄ�=z�=ӏ->�&2>��p�!;���<�<�Fj=���=�$>W??=#�������`���b��8�d�(��g�=��%=�C�;K��=N=r��>Q-��A:¾K[�])�֋,>h��=>�=�v�=���=�����|�쾠��u���~&�>ŝ�>J�>�#`=p�>���=�]�=���=A�=�Dʽd��=Mk5�s;2�,=��+>�R���<>}����,L_��U*��T>'��=�v=jc?�Ձ?�j?���>�b�80�6��.�K�\��=�/0��s>"��>;<�mD>ǝ۾�����K�̾�\;�22!>$�m<��ܽ��=���=8Ο��?���>#��;M��=���>/G>/�->��>��&�=�����j�!�@u��`e�v������c_=��#>��I�H�&�����&j������=�>j�;K=Ww��=(�������ol�}�[�eq��Zp���ξ���̄�z�g�1SI=��9CUc�9�F.�7����8���Ys������v��]?��-�M��s=؛>�?���>VΧ>�P�=Ǭ_��z�>yV>L�~>Z� ?��l����<7��>�b�>����:
��Q�=�=>�;�<N��=�^�=U��<�{?=Ӊ��g#�Q�ɽ�-%�F��=���=G�=;�S>#&���=#1�> ��(U���ž�DY���7=k>�k�>WCϽ�-�=Dɽ�"�=��`�zP���l���=�>e%�>�`2=H@>��:<�����=$��=�>��<�
�TN'�$���~=n�[�="o\�wC�=�|<0�=�1�=E6�<ew��H�:?|q?�f?F����f�x�ƾ�̷��`���W��On�ŀ�=�@R��É�N����4�$���j��T�1�>R�}>�Y>�@�<����gC�y�"=iH=�G�#>���<1IU>���=��=9��=ڼ�Ž6� �4�\1޿q�i�4k��?%����vc���lB=�֨��̘�?�>.=�~�i���n(2=y圼a�K=�����j�4��<�8��Vi��A����0�=���߾h���b��>��P�w>Ɩž�v�>&;�֔	=G�(����,��;����<ƽ��>���=������=���>ә>����p|�r��>̹�=���>��~��=���=�V�>��=>r[�=�=x!��Ľ'��=�>.�� W�u�B����=CD<ƾ=����� �$�=��S��Ż!�ƽ~�:<�ɧ=��>P��=��>p�Ҿ˥ݾd��{���g?>:Kd>ꢐ>"N=e��>�{�<��<�fy���d����0R]>W=>��Q>�@�� ?�����⋾-�R�;�=]�>
��=��@��I>g����=������>d�p=(�.>���<��p=8`=6S"�~�X�7=B?x�{?�Dj?�U�i����i��`u�>��aﾾ�нF"~>���>���h,D�~����I����ws���q����>b2>��->k�=�R��V��eҽ3�����">���=�:N�Z��<\>7>"���֬�)� ��̿�"p������J��ڪ���y��|"�B�>GC���|�=��s���5ߝ���>�D�<d�s=9?ǽ0�]���	�����5|=���<1����62��3�*���u�>HW��U�->��ž�)�=
���k�*�񘦾����JQ��4˼7@=�{�>�Q>�F�vP�=h�9?��e>\�=Xd�=��3=�u�$�F>�m=��>J8�<A>>�3>ز>w�T>Y�>1ԽQ�1�<�1>:P=����+�l�-�H>;>T�=ef>M�b�xɑ��F�qJ���o���&�}>�<�>U��<��>p�Ҿ˥ݾd��{���g?>:Kd>ꢐ>"N=e��>�{�<��<�fy���d����0R]>W=>��Q>�@�� ?�����⋾-�R�;�=]�>
��=��@��I>g����=������>d�p=(�.>���<��p=8`=6S"�~�X�7=B?x�{?�Dj?�U�i����i��`u�>��aﾾ�нF"~>���>���h,D�~����I����ws���q����>b2>��->k�=�R��V��eҽ3�����">���=�:N�Z��<\>7>"���֬�)� ��̿�"p������J��ڪ���y��|"�B�>GC���|�=��s���5ߝ���>�D�<d�s=9?ǽ0�]���	�����5|=���<1����62��3�*���u�>HW��U�->��ž�)�=
���k�*�񘦾����JQ��4˼7@=�{�>�Q>�F�vP�=h�9?��e>\�=Xd�=��3=�u�$�F>�m=��>J8�<A>>�3>ز>w�T>Y�>1ԽQ�1�<�1>:P=����+�l�-�H>;>T�=ef>M�b�xɑ��F�qJ���o���&�}>�<�>U��<��Z=���d��.���,žݶ��&�>i�>䵧�D	�>����\ o=M󟾷Y0�� ��:>f�H>�i�>�>����>�ye�*᝾�6>q��=�_>;�=�.|�k{*����>��k���
>��=�D>:�f=I�9<p�ݽ������<�J3?l�k?��o?#^G�G�ؽ0�z�R��`���rv����I>f�>�1<я�r�����8��E<՚>����>�j�>�O�=3�L=j=ѽE�<�`�������R>,�'����=�b󽇕J��J=�q�>�ݻ�gD���$���ҿ��s�2?���~"�25�2?}��n��ץ�=%]���>'9����<�]<���=l^M�s]˼�½����+�=l���.˽&YD�F���������6־'}>������>KZݾ{�=ʑ��&����(�5�D�S�$寮�j>�@�>B�\=�c��#��=���>qʱ>�n�=�&"=6�>�./�Ǧ�>k>6�3�z>�w�=B�h>y�>��&>��E�i]F=�I�v
�=Ak">�T�Eq���^&=[3+>]�S>�>zj̽�]<�[�=��=� >�ঽ��S�e�M=�M>��B���Z=���d��.���,žݶ��&�>i�>䵧�D	�>����\ o=M󟾷Y0�� ��:>f�H>�i�>�>����>�ye�*᝾�6>q��=�_>;�=�.|�k{*����>��k���
>��=�D>:�f=I�9<p�ݽ������<�J3?l�k?��o?#^G�G�ؽ0�z�R��`���rv����I>f�>�1<я�r�����8��E<՚>����>�j�>�O�=3�L=j=ѽE�<�`�������R>,�'����=�b󽇕J��J=�q�>�ݻ�gD���$���ҿ��s�2?���~"�25�2?}��n��ץ�=%]���>'9����<�]<���=l^M�s]˼�½����+�=l���.˽&YD�F���������6־'}>������>KZݾ{�=ʑ��&����(�5�D�S�$寮�j>�@�>B�\=�c��#��=���>qʱ>�n�=�&"=6�>�./�Ǧ�>k>6�3�z>�w�=B�h>y�>��&>��E�i]F=�I�v
�=Ak">�T�Eq���^&=[3+>]�S>�>zj̽�]<�[�=��=� >�ঽ��S�e�M=�M>��B�w��>Z��������ŷ���,��S>�o?�i>`�>;J�z�=�v�¶���G>̖�=�(
>G+T>c��=Jw�>4y��!۽���<_y�=��>3,�=]�c�͡�*�G=�Ҍ��|?�0��*>d�>2I#=��Ͻ#�]�B$E>d�ľ�R�??q�?/}?[��>���W]�t�;��7׾BH��.X��_��=�=�?���Y��Q��Gz=��VԾi�=���<i�O>5ˮ=>�t��
��d��=�ܑ=1+�=n:�>�kA>i>#�;/3$�դս���</|<̍�:6��3���뿾�j�
9U����n10=q�6��5�ۋ�a�i���8�x=�\%>Ӈ�=y�S=P��:ƿ�<�h�V���:�<A���8������Dľ���o��>���Xq�ٍ���ܯ�����D��k�j�������Y���s����^�>�c���o�d���?g�)?i�?B�?���>��>C
�=n��>	T�>���;�팽y�,;�.�>�.�>N�>�%�3[C�<�X>	�̻�l���k��=$�<=�a�=g伺�t�w7�=2���7���E�=Z�={K�=���=.��t�>+������0��S'�X��> 0p>��?3����P;2��o(ý���<_���ԓ>��>��>5�>��H=�I >5�P>�/?>�;D>���[�=��a�����n���9��=�н�O��ϒ��M�<��=�>�!�<d�l�nHν�.��(�W?�qT?�d]?�s#=�=�3���!�\���%;�=�b<c����5�>��y=>�k��뵾���� ��h��<z�=�V�={��y%��/.=�z��D.<��=�")=��ͽ��G>c�>�/>���=��>
}:;7��c�����n���섿��ľ*1վ�]">p=r��=�G��u��
���5�9�r�( W����=x�<)m黒ă;t��<��=�3��",�ݮ��W����]�L��MSg��]9T�)��b��u�<�������z�z��{�'Hd���>ZN=�s>��D=�7��D��T�6?6�>��T>x=%�w<�>�Q?�=�W>)��>�u�>�/�$�߽�^P>ͼ->�}�>�ށ��?����=^�=��=��=K�>I<@0U>�`�=K,=s+>�KD>�)"=gA����!�u�#�a[<:�`>Tg�>�+;�y
���̾(V��9�\�	��>k��>6�%���M>Y��=�)1=ʰ����t���n>4>⏛>�O�>�
{>+wj> {�<�B���^㽐%b>��;���;�a���u���=�Aý��Q�y>F�����|�!�=�f�;�)�=nVZ<Z�<vn?��q?�GZ?�jq>��������@�p'�<1�=?�W�e,�>�t>t>;Nܿ�{���3�hY�p���Sc�<C+Z>���=�X9��� �s�V^�=]�>=ݼ�>&�=�G�=��<�h�=�ɼY��<��Ǽd����￨�d�����T�A!8��g�>��>M��K�<)��eK"�uս�!KK���[>�ʴ>/L�==_=χ�=sP>59��Z�������Y��J�ғ��l�t�{�gG�:�ڽu�y��X���}Ƚ�Ǌ=�@>at�����\ؐ��2M���?N;j�K�� �2;Z??1=�>���>�ע��)�>U�>{��>v�?]�=�n4�3�རb>_P�>
2�>r�=B�%��i2=���<��$>͹����Q>��O>S�=�E> b]=�"�=z ����E�ّ=螂�D�Ҽ!X�0ƽC�>R3�>����>���"̾�x쾲�A=���>�4�>�'��v
>|�8���5߾��X��
>�U.>�$>0]>E��=YC>>���=�}�=L�;>$oq<��N>w�>�Na�i�G��d>���=y���m��<҉���5�:L��ٲ�S�=l�=5BU�/q?A�n?�Vt?.a�=b��2����*�ֽ4���UFn�T�#���]>
c>.:缫P����q6������́�ez�=�,�=	+j�K%>�3�_���\��>��`>@#<�h؟�ci=]$�=Iѹ=�^���k>p+>��;�EνT���ԁ�����t���1����mك>XL>���=�0n���l��E����=]Cd>Kd=���֨�<�Մ���~�x�������F��־�ξ���yp0�F��=��7����z[*���<C�M�亨�=m��s���[R�roH��/�>%2��8����3�JT$?�o�>~?p:-�_���{>[��<u��=@%D>%WX>x�0���-��s�=N�v>���>Gn�>�V��p�=<�=)L9>�c�<x��=�>^���z��=�ͦ�Ы����h=V#3��"�E�4=n3q�1�=u-<#�g=���>�t����v�Ӿi*�Y�8>��?�	?`�6>�L�=o�?�^��<������9��+>�G�'�=����=&�(>ZQ>��>}�P=*���d>&R>�>�J��d3�x�>o��&�R�.�X��Y̹=実=�=��μ�R$�?^�<�N�?�w�?Y-�?l?<����D�A����ܾ� �_�5�}*"����>��>����_���p?/��~=����0��#�=���=��>�����>G��8��:�*>c�X>�B~<"&E>�R4>���=A��;����:=��<Нܺ9���2���݊��%޾~p��ۮ��C��`��F��8P��H}=w�&�4꽮^1>�w�>�<�>q�>�=l�@;��>K�#���>��������r,��������׽N"=l��#���p�/m�$���%z���qR���5b���ͬ����?~sq�l����戾�D8?��?�d>��A>S�h>��>��>�]>9��Z��_�=�n�>�40?�'? @>u�@�0�G�P�=Z6M>[��=��=J-<�7b;"q= 'n��j�<.K�<�a>��=�n����U�A�W���6�=�H|> 4Q�?c��tݾ�T�_�b�Vi>Q��>rY�<�N@�a䪾Qݬ<�p�P�a����=t����3=����I�B>��>�R�;�����.�+�$>ؾ>��=�or�sf>���T�����"t����|X�å�<�gf�;Z>�'=��P�ev?F��?���?�;?������_��3��GV��p���<=M�>]P�>t�<�T���:-ȾWM?��)�>�ۖ=۲��->@�=���=C��=�_��>B���/>kB�:��&�c=��=��=X�>�%�>�7>E�<�%!�t�� ������V���^����_	E��>P�>����f$>[�����dս}g>�z>�=���>n ������
*��?�����:�� 5�6������j�Y>��ھ:;W>k���h��q���\!���;?鵾�+=��޾�_P�+{�>@��Q箾_釾�\>*=�>~��>8z>�Β>����^�>�Px���A���>$g->_�?TO�>�J�(�d���=E�����=خ�=��=�G;>B%�=:-3�XǻeE�<��=��Y>�|+>����E�ν.r��� >Z��=�
p>���>x�H�/�S��痾�3����y��1>=xZ>��������x1��:�A��s��y8��O(�Gžю�(>a>b��>H�=|��=q>ؼ�ߘ��>\A���!>�Af�����{;J >�%��V"�M���,i��+�=�G�\*>�v�=-���9�?
�?�Bw?U�->����1_�j��/3���"��=1N8=cI�>���\�ܾ/�ݾ�#?��W��Lν"�=+��=#�=:wF=��G�fK�����m1�>�k�<�׽�`�=��">�>�]f>��>�@�=+�;�
5��]I�Z���h�t��<ľGK��^��~'νF>�7I����=3��=K���Z�νɁB�7\8>Zpw>~hD>h�C>ə���L���t��
ؾJiľ^&Ǿ��ھ���F�=�?�s=�셾G(��aO��F0�J���y=q���{�W����ľ�뒾��>�G� ���q?���>��X=�)�>�wE>�8M=Q�\=��>[<U<�=Po? +�>�T?���>�^�k����ê=?k�<��>��j>��Ľ
>��=�Ǩ��y>�ߞ=|\�xd>�"|=�Q9�!S!��rҼ:�|=[��=u6>\�>�@����@ھwa�����F%>6�>�FI�i�>�˘�9h�<����L���t�G�%�b1?�@>��J>��F>�|>��=r̽i5>�d�=	��<� �{E܉��=C�� �F��#������^�p>;i꽖�לP�Zg˽\��?҅�?��c?7��>A{9�4����v-�C�?��>��=��1����>r�C���q�1{�t��>FG�==g�=e�M=��>�e�<Wg�;�r���%ž�>��=���<��>c5�=�ϥ>��:>+j�>�R��;V���\���X��濋���]���y���?�BG���5=@[����|�S0������s�C>`Ǯ�]�6>��^>\�$>Pi4>{I�=�t_���ʾ)i��i��^3��X$�l���"'��9�>]���QI��[Q��ě��(���C����=����eE��*�J�cn	��]�>o`���\��������={�o>0�	?�U�>���<p��Pc>�ʽ��:>��
?:&�>�*�>'�'�����I"�i4���j�c��=��,>6��=�>��>��=�,>O\$=��K��;�=~��<U늽9|*�4��:�g�=�V>�*�>��>�Z$��镾��n�)c�7`r�<��>Y�>��<���>�:����>W����?�9�T8=�@?%�>]h�>jK�=&�g<�X?�ѹϽ�QE>a�G>3l>Qrb�5K�=p��5fr����(۽�9�-�&�
��ZP>9�����=�t����^��͆?���?��W?��5>� �1hr���
���C���>`*����">�M>d� �K����1G��g���B���J���&�:_>���yx=�h
���C���?>���=7��p��=�Y:>�̛>��>O��>U�9�K)ƽi������xͿPI��>�޾]6��p�6,��s�<�~<OL���-�I��1��|W�ם>5Lc>ϧ���6�x��$�3=�f�>)�>�����8�>�����{���{�>�H��{�s>��n��<�=I矾}�<����<3�n��4� R����<s�>fٮ�7PȾ$�Ծ|��=���>�h�>���>Og>�$�?�?�qp�h�>�d?�>��>� ���签��!��o������=�/�=<�׼�6>���=���;J(���>�,�<S >�!ü�V�<����gj�z~>�l�=�w�>*^X>1�<�ꔾ���?}���j��qq>{J�=��R�)D=�	��w�=�����V����9��c�?3��>DK*>�>��+>�<v�?�u�w>$�=��R>�NQ��5G��潟�=5oz�<.���H0�TLp��_=*��*�����ｄ����]?�lq?�L?���>��c�G�����l>��>���8P�=�V=8��-@�1���;¾So�V�=*h�l�[��L>K�>5[ �n�E=�u�!�>��0>�X�<��=�+�=J�>���=e��>��=:ؽ��G�ކ<������+��~#ھ!������A��?h?��D��r�6���A�ξR�z��ݏ�4a>j;�<���>t�4>D�=
B>��=�>l�꾷㪾�{�ek��;Ł<{q>����������YؼT�Խ��(�|�ͽ4�о�q��e慾�N��?�0�XP����~��m)>��>��>�A�>R��=G��Ž?~G:�6��>��	?<�?��4>~C�����I<��Bb2��R�TE=�X>`*$=}*>�=~2�4و<���=��KR>j�-�憴="Gy��i~=�e>z&�>��>�hh=m2��4��	_+�<������e=��=������*�H�����ƾڃ����V=�h�;��\��l�����=�ã>R9�>�4>?U����G<�6�%�4�w=�K���j�=��=:���9(�pڙ���޾���(���T�=+�$>���>Ē"?�vC?��D?T�=-uվ����	Q�=Q�=��>�?&>��<����C5�R�4�5�G�Q���q澶^F>`�[�����,��=�ē��N>\_
=y���Ζ=���=Z��>W�C�	�>���>aÙ>��u>�*j>u"V>�Z�<����39�J�Ϳ��;�oϾCt�M�7�E���e.�=Qo������Ϳ��>.������L%?���>�΃>��g>��n>h��=J����U���Q8Ǿz��`,�U�2����d�/ͤ�����<?a����=C��\�<�%��`%�K�׽�0����>�Tc>!�Ͻ���H�>���>;��>���>Wݏ=�>{�>�5�>Ӕ�>ILI=E�>]�?n��>���>�=��X��;�轫�߼��T>�}C=9�K=��_>�頽}�`=3�?=��K=��~���;��>���=�14�o�T�\Ō=�XP�-ܣ��n��dоz߾�6���&�>���>X�����:+*־�������댽�{>9>	�C�}�^��𯾐�>9A>a .��l�=s0=��3���ݽ���<�P�=6(->����Ћ���=�5)=��g<JtW=C�=�%+�>SC�p�>��?�>:?j�?B[�|�!�k>Ҿܮ���>䘓����=s�9=6@>$+��4���0(}���V��)������}���#>�^>eg���6��ۥ��􃾩�h>h��>(N=�Q>��>�п>*��>ݮ�>��->�O;�"�@�տx�� ���������U���2��~��2'V��i�/��e�����*�z<��ѧ=q��=�6>�>s+D�g���6�����=�5⵾ғ���=󒐾�f�v�ξ
��=mKi���B�S�T�@��(�о��½�>y����>�܁>ޞ=-.>���>�e�>
Z9�1�=��i>^�'=29�>>��=ء<�@=Rc�=&GA>�5�>bLf>M��>�+�;N,=o��=��B��?>��>��=�C�=yE��΁����=Ks׽�$�p8W�(bc���B��3.>�]G>�o���S=ۊ�������(���5�T��>�C�>��=;��xo�vf��LnE�7���5>�r<�������Rܶ�1
{>ba>Jy�=���<�B��Yt��uϼ�����7�=v��>�����f~>a�<>�o��-�z?�=�>��S��#L�d&z>�	?j�;?-�0?z���$������R�q&E�ig�=.�=d6��� �>�͇������O�����6����趼б=f�E�٭�=��=��ܽ4���U�0U}=˥'>1��<=w�>��?��>,�>�,v=|�����ξj��o�Կ�վ,o.���=��:>5礽�6�Hr��`܏�#���׾�[����?�=̏���&>�>(�>y1���q�)�뾚f`�"�r�ɾP̅�i		�|���:潾�Ͼ.^�M���\���7=&�j��GƾHd]�q|��>�)>�t����Ƚ��?@�>���=b�>\����6>6!�>�(0>kU�=2�<�C>*h�>���>��>�/=�3�=��Z���s=��=��f>8�=�(>Ya>��м�v��=#��3����2�_��=e:_��߽cT�>��>RY��|��,���n۾M��e1�Ң�>��w=-z��om��vc;^I8�e඾�g��ђ�>�%l<� g�`�I����2�>V��>8߀=��;3m��̝��f�̽�$��j��<�'=���=�p�<�v��:l���Q=/ .=�wK��}|�ݒ#�Y%�>[0?�[>?6:?2}���y��I����2�����|�&>ք?>�
=���{?�!��d۾����=���؆��֖=-ic=/�>�<w�K�1�I=+"�P�I>��V>��%>�'�>�%6>���=yE�>- �>����@h�o��5����A���<���JT�hiQ:$�5��ˣ��:��ɳ��/;<���A��>LU>��� �Q=�'�=�J����c��Һ���-)�o�_^�������f��b�<۪��!��=�i��T�Z���ݼ�|��/y���L�͍��u��>p��=A5>��=��?	�>�3>5b�>�^>6;	>��>��Լ�>Iz�>��iH�>�c�>A�>W`'>�d!�C��?{�<��"=�-�<~�M>8�y>Iu�=p�=~9�k�󽃋0����u��=b~ýkz��3�	�L|;>�ɰ>RY��|��,���n۾M��e1�Ң�>��w=-z��om��vc;^I8�e඾�g��ђ�>�%l<� g�`�I����2�>V��>8߀=��;3m��̝��f�̽�$��j��<�'=���=�p�<�v��:l���Q=/ .=�wK��}|�ݒ#�Y%�>[0?�[>?6:?2}���y��I����2�����|�&>ք?>�
=���{?�!��d۾����=���؆��֖=-ic=/�>�<w�K�1�I=+"�P�I>��V>��%>�'�>�%6>���=yE�>- �>����@h�o��5����A���<���JT�hiQ:$�5��ˣ��:��ɳ��/;<���A��>LU>��� �Q=�'�=�J����c��Һ���-)�o�_^�������f��b�<۪��!��=�i��T�Z���ݼ�|��/y���L�͍��u��>p��=A5>��=��?	�>�3>5b�>�^>6;	>��>��Լ�>Iz�>��iH�>�c�>A�>W`'>�d!�C��?{�<��"=�-�<~�M>8�y>Iu�=p�=~9�k�󽃋0����u��=b~ýkz��3�	�L|;>�ɰ>�Uc>�]����Ӿh'����V(G>}�|>�������>sʬ������m���T���_=hS>�%�>��[>�ɠ>Pb9>�φ����H�">U5��<���;>�(D>��}=����]�>�i@�-�99]�G���NR9<�i8>��;؜����?�-�?7�Q?�Q0�Gx��S�.�Ҿz#?�Y�b>z�B>RD9�/��){>�a���#C����wt�%��sH=.0��;�=��x=U��Fk�=`R$>l����7>S
�<Ҩ�>9�>�y�=�,=��˽)����q��|���g1������e���������F�<򣁾Dܙ���r���yľ��=�1�>{�<>x�,>q�w=mݒ=�>����/��MǾ��/��|T�����-�ӽaj��� ���>NM������ƽ���:&_�qŨ�/~���m�;"zi��b?A刾8�����<��mE?+�?��>��>��R�X�.>��> �x>�>/_?�FT[>D�>�?k�=r6��@+<��a>E��<΃罍;�=��"���(�=33�=}-�<`���j�]{4�ϊ>�@d>��=��ν�_D=��>[y��"��t��B"�ŰĻN��>uf�
������>g�-���g>��Q�`}��������ʾ���_�=�b1>&��>�>�>�GR>8�=��<x���W׽�E�к�>fA=�Wػ��<�m��*��O�5:����P��x�>��>Zb}�	V�?j��?�q?<���b�V1��:߾��?��e�?F��=�1
�jY���5>��ƾUF���r�[C���D�wa��Ss�=me�;��>>-v@�Y4�>�����F���l[=�-�=L��>j��>�ٓ>��=�3＝mv�ƪh��H�xN��7&ɾ���v$/�����a�;+ҕ�T�Ⱦ�4�=�?�/���Ə"<�l>Q>.Ö>�G�<�	����6ε�/5վZ�߾�S��\	N�?�E�a++�.�b�����*^�e������r�#���F���4���&�V�8��U�� 9�M�?S4�s��&�>�>N?*{?:	>?t�����!�9��=�����>���>�i�;>�@>ߝ>:l?��>Ⴝ�WM=���e��=�9g�'�2��F>=?T=^,=N"�<�3�=�<����b:��N���>=>U�U>�AH����{��>x徽e�쾵��괡���k>�?� �:��+��>s�9��R�<Q쟾x�޾1�i�1"�>�K�>���>֚�=��>�
>�ԏ=���=��
=0"�����ڿ[��$>��ƽ09[�'��=�	��p��ۡ,����=mp>�T�=]��
^�7H�?���?y��>���SZ��倿� �z	?*���_o�>t�@�d�U�03��1Z>Mc���U$�|��L龤�u��
Y��>Ց=�Yл5[�=�P,� �p>�?<�P ����=�'�=ީ�>d�>0�'>P<�;K깽�L��Ȱ��$�@��KD[�FA�B�+2A�&�-�t_�=��&<[�1�n �jgȾ&jл�+�>D��>2��=P�M���=5S,>0%E��=��R��-%��B��Rp�G�����ק�U��=R�7�d��h":<�j����(�ӽ���>��v�7���!?�F���۾yȰ>u�:?J?7�>cߡ>�ZI����>���=V�>�^�>� �>�v���#t�k/s>F?IsF>��{�aVQ=s�Y<�	�<m��<Z=D:�<-c_�n�i=��<�X�<%�Ƚ��n�2��<���=���&߼��A<���=�n�>�򷽄�Ӿ���:A����漩��>�v��l���i?�]C��
�_5��ܺ
�8�r�)�q>AC�><�a>���K�>x�>&�<,�=�ļG.�̪6�r^;�bv>��%�{�νr@ʽ�4*�	��S/����4>��K�>}&?<��Z�:z?1�?j2?K�����W�}I)�I�	���>.:���c�> ٠>�e��!��ط;>ŋ`�R��*�y��V¾ްV�!�y=3��=����@�=Z�#<��E���>�����]�S�>��I>6�>Hm�>�O">��2��.���:������_���4+��w�%-���܍�v��=����9��2^6>����$Ծ���>�Ԗ>X�>*^>��X<�����"��9��������"���f�t��_�H�Dt�=sH=���1�>ꥤ�Y!��?�ͽ�Z�s�=�Ĭ��l6�Q�����;�&?�A޽	Ͼ�ɹ� .)?l�,?�$�=z?�d<�>Ҿ�D�>\�=�+�>)��>P�M2%��>�?�u�>c�}�pL�<��>���=~���p��= �0=3�W=���=$0�=���<q6�=X�!��}�����=ɷ�=��5>�b}��گ��Uc>�]����Ӿh'����V(G>}�|>�������>sʬ������m���T���_=hS>�%�>��[>�ɠ>Pb9>�φ����H�">U5��<���;>�(D>��}=����]�>�i@�-�99]�G���NR9<�i8>��;؜����?�-�?7�Q?�Q0�Gx��S�.�Ҿz#?�Y�b>z�B>RD9�/��){>�a���#C����wt�%��sH=.0��;�=��x=U��Fk�=`R$>l����7>S
�<Ҩ�>9�>�y�=�,=��˽)����q��|���g1������e���������F�<򣁾Dܙ���r���yľ��=�1�>{�<>x�,>q�w=mݒ=�>����/��MǾ��/��|T�����-�ӽaj��� ���>NM������ƽ���:&_�qŨ�/~���m�;"zi��b?A刾8�����<��mE?+�?��>��>��R�X�.>��> �x>�>/_?�FT[>D�>�?k�=r6��@+<��a>E��<΃罍;�=��"���(�=33�=}-�<`���j�]{4�ϊ>�@d>��=��ν�_D=��>�k<nž��)�M�Ѿ��H�,��=�UW=�8s��1>m컽�T�ͩ�Ȕ���Y��=�Ϊ>Č>jA<>��>RC�=pz��C�� %b>� �<!��Pҽx�Y��A�	1>�2�du��kҗ��*ֻ8�=�$=���;�K��
/�=�:^?X�W?��??uA�>B�8��B�K�ܾ�إ���r>��?�bQ��?�)d�B���Ҏ��dھ_;P��,j���	;�>�໽��=�s��`"=��3>*0O>�9a��|�=�vz>�s]>�܈>�� >�=�=�F������� Y޿�&��a��,��#>���<|��=�����X�=D׾D��=�ݻ����>~Y)<���=�ἥF�6D�=�f����b;%�_�tʁ��#Ӿo����@=���=�Q�N,ʼ��Ѿ��l=���� i�n]�����(	7�d'U��C�sI�>n��=9�ʽ�ӆ�¦=#;�>㉉>�L�>H��>@�ƾ�t��^2>5��>Q�>�p>i�<⑟�"!=���$���Խ�s0>:*�>bf��L�<���<M���$?�=y�=�s=�z"���=�����^���hڽhF>U`K>�(>>Y�>�Խ�./� �r�,sn�V�`�#d��_3>�^�,��\��m�L���;i`��<1�L>���>|��>�Yw��Z�>xg�;�n��Xӽ�ix>��>�G����E<�j���uG=��`�����wfA����<&�m=C,=S��m뉽�"����>�N/?��?�HV?��*���1�y��)<-�mڛ<��>r�<�ܼ� ��>,��C;�E��i��͆=H�z�>EZD=��": >�=��j����q>�=�����>m�>xޏ>��>��X=M$��gp=S�=��۽e���������󋪾)3�� �Q�Y>.d�+fڽ��9>E$��L=�؆>�͈>�+>�B�=^�=�n�=�x;>�E��L<)�|]ݾg�E� �����ź��JT�=u����W=�y��iü�uT�te½�g������6���������U��> �h>D���\n���>�)?���>*�>��>��M�>�h1>y�>YO?�>�}>,g�*�.,#�ʻ�S����Wj>��>�S����=���=�ʂ�0��=>l�#��=e{����=.�ݽ�o��Aq�<�(�=�:>Ss!>)�>�	����G����Ue��U&���<��*<��*���<Q�����4��=��ypk:�%Y>��C>���>|p�>�O>��>?|,>+�'�>z�<u�=�*>��=e�ͽK7��)���d-:�s�D��T�<� �<!��=$�l=�9H��<=�g�<g�Q>�E?�v:?�hC?���=A����ʾ�����H�NU�>���>Q��=|愼x����\����龴;�x����E���_�+�ܻ��=1��!m#>����s�
��=p.>���=��T>��>��=|O�=%w=˼�=�x=̴��� �Ùܿ�@���i����2��[��>>��?i{�A�����<�A>)�=B�>>}�=��=��8>��)��T�<�<�/��óʽ�{Լ4�ͽd�վ����q��9⻛����]�r�kW��%���Ͻd ��-Ž��b�ɨ1�����>� �>45��	[;�V�>��>g��>�_�>i˳>e�����޴�=5%�>=�{>�V=����&��tl��5ɻ^�½?��L�=�s>�#=��c=䄤=�@=�<��c<�=J'=H��L�L���5�H��#v>��7>��>��>FڽTM�}.Ծ^���{>���<��>R8�5�D>�RǾ���3�¾�׃���>-�>�o�>�K=���h�>���<U�����e���>'�g=�] =@\�<w��G�R=蛝�M��j��=v`���d� ~��oؼЄ���ͥ=�'>]pN?Y1?�?�e><Ծ�/���� ���k�w�M���>{!5��z�=,���5d��IS�� �ؾPV��(V��fF����>lF�>�=����=�ga��2���`��C�=� ��G�Z>�ܽ��K(=�kV>ls�=�=���9����N	�mꭿ'跾ػ���b����y��T%�0G־'�@=g���P��"�!�<���=�'�=��V>��3>?P7=9��.~1�*6,����t	ݽ���$�1�FH�=ݼ'���=	#�����<�~ý�v�>���_�I����6Z��P-=j��>��>��<��>
(?���>|(�>8�5�GS>��ݽ��?A��>C��>ll>��P���l�*�\��
I>��>6����/��(Z>v�>,��V�M=���=��\=i�>�5��z
=TD�=��<;�<�����=P��=v��<�j>�*�>5iu�'ʾ�����f���4j>��>�>2�#>���=�� <)����'��؄<�� >9�f>%B >��Q>��>�������ʜ�t�=�Z$>���>M-�<��齵%��lw�=_F=h��>��">�C=X6M���\��y��Ä��>@�??c�J?"�)?��>B ��J �����(��u��.����u�G�>w>�Ҷ�uwҾ��žC�
��"�0�G�Ȋ�>���>Z�<M��=Ѧ��P^��J���'� �<��	=7O!�R����^�a��g0>N�]>�6�=0=��᛿�Ͻ��	�z���l�c{k<D�X<4����C�>e�+�����[��>� �=.l
> TL�(�������ZC���K9���O%� %ɾ�V��&���$u�.���=��=阾]����ս�z���.ĥ�nz�,�����֟>a�?>�!ͽ�"���� ?��>�� >��L�0j=+����۪>��<>kb=>����-�&o&=ö>�8�>��>޽�%�����<�[5:Wr=��=��$��u=%�#>��뼗 d<�*u��X����p�A=��+>��!>�Ȥ=]=EO>�P��,[���WJ��#��	B�RA>kd>�;�>ϡ,>�PV�n��Pž�'���ν�"���<��>^[\>�_'>r�+=���	�B2G�GG�;���Da_���?>��V>8�=w\�����~���Y�k�d=��Z;�-ռ���<�?d�Q?�>a?_8m?�e�>ҋ)�{�=�x�q��$뽁�B<�?=�@>�?p�>��kȳ����A�"���-�v�����r>t&�>@j={�_>%&�=is_�uv�<Î\=|`h�Mx2>f�=e��>H�>A}M>8�!>,V�l�Z<#��O����Q���'�f�.�5�m����8�c�/�_>YcS��+�>_q��B�/��]����H����a��<���>ژݼ��{��-�b�齋Sn���I��Z��/
�z��=�C¾��=�峾K�=�`׽;w���j�M���ｽyH�M_���<J�R��t�<�*���>�?���>���>A�L�����b��q��r�|>���>���>��>fс>ݗ?��O�>�l=9RϽJW�=RX7>0AN;���=J�H>�����B�;����="�=:�R=�ʧ<�»6#r;6ь=}�=-�=�q�>�8=���������%ؾ�m>n�>�PI>�?˽�g��=Q߾����r���>�ۙ>�m�>0I���SA�s�>��>����w�s`Q�;֓������">?� =�}=+=#��鿼��>d�Y����n=�B�=�:�Ծ�>b8+>���>��p?1�d?M�?�p�5�-��<k���;1SK>�J�> �/>#:(?.�">)�D�#'0���4���5��d������y.>܅�=�p�=Y)f>T�s=�3_��ʕ���T>뮯=$�D>�>Q>�R>" >?�>�1>�]�=���=�������5���)�.�bž��6>M)=P�>�mY���x�LH���[H<�a�<>��f�>"��=��D>	�M�߷��������K���쾫x����I��c*>r�����O�2;����������;��{B޽�ͻ�Tzܾ.ͽ	����2�=	=��3�!���@m>��1?���>�ɇ>1�r>t�~=��>���>��Y=�?��r�I�>�.>�Л=��>��>j��=��l�
�>L�&>ǌ�=��<��">̞��I�\��ɼ���<O������<�Q��^E=^Z�<�9�<Я=��w���=T���Wg��!�þ3���v��c">���>*����B��DѾ��u��Fξ Q��CҽS(�>�3������ˮ��f�>�1�=���t9�<5E��a<,���=���Jb�@ؽ�g�P�\�ٱ���=���=��Ƚ[�3<n�c���i�>ݧe?*�?,�h?���>�/2��m_�q2k�X%��cP`> �I>�V?غ-?� =Ev�*�ݾ#Ø�=�̓ɽw��s*>td�=�ȼݸ	>����o�����<Z�&>c�b>M�>����>ӻ>��"~�>��!>�+�
E���Aҿ���E����\��& ��>��~�=wQ�:�E�r���V⾗w���믾�F����=|OC�eE<�5>%+�<(1��ҫ�X��;���ƚ�ѯ�MI��	��= 4��(���+Oľ�������d�C�ٽ�9<�'i���o�
�M����>�j+>˦!���D����>�H2?S��>��>vN�>�/=6P�>nI-��>�=�fT>�!m=A�=>�>E��>��>g얼οK��Y >	s>�^>�?>��r>r_��23���`̼�8�=�S�=!�I�h�����d=�Vż�=��=��>�Z�>d�>B���U翾 �X�cG̾���=���>�v�>��	��^���f��Jξ���I-�>��2��5�%5��0ڿ��U>D��=ߛ����=�f�����}�H)�k�ݽ���ïw��Mż���=�����G���̼'�6� zԺ
�ν�2�>�
)?�~z?�Xl?\>��W�K+��e�����Y��>�d�>���=���>>�/���8�S���"��:.�nW���漟=�]�;��8�LX>�K�=����3�=Ь_>x;=I�>A_�=@@�=�TD>���>˕=��F>zM�=yOͽYR���J4�v����5�Dr��<o��<�/ʽg3k���о��U���q�� j<>��>8F>T��=Q2>gSk�❓�P���ݔ��������)�N>0�Z��=3z�#��<������M�|����ϖ���Cܽ�sj�N����ɽ�>�UF=p��<�/7==�?v=?4�>��b=m/=�I���>_��>�vy>#N�>&��e��>��>�ը>d��>6(�7�۽5�= �}=1�=��<S2>����D»z�~=V<�=⤽;��A;�<�W$=\+�<F�k��$ڹ��>��>�ѷ=Ր۾����� �P����>��	?Ǌ���Wu����<*c�'\�ZO����>* =�n^�#g��)þ*R�>߃�=��J���X���<ּ��ͽ��d>����M��$p=ID�\R"����<���zx=d����ܻ��,���-^>�-?oo?�+Q?Ǽ>�	��9�L���C�Vn�>�g�W)9>���>ŢC�g���>e<�X����_��:f`�;Cw�h��=ELA>s��<��>X:���1���n��W�>��>~!>&t> �>�=��1>��Q>=Gp>pB>��I���񿳟п)[�����.����M��F��K�ݽAD�7��>0>!<��ԽA�=6���U�=O��>�s�>9',>K5�>\x��d���w_����������I�����=3���\�������2B==7�L�����MП�d&
������P�>5�$>�=½$؟�B��>Q�)?���>�R.>�ʀ>��]��I�>��=+��=��e>�l=�_�>��~>]/\>M�>P�������y�=���=	ݍ=�>~ot>U���B�a��<2�=�E�c��t�7]<m{=���>���%�(�nb�>vg>#���S�>�t�c�����>`�=X�>��9�6���ٲJ�LӅ���q�ƍ<��,��ұ��"��J�F>r�=�d��0q��N�=�\W=���0@꼱���q��:�=$�{���=tٕ���(� ��̺$���2<�s���>L�m>�,�>�F?��1?�@�>�ә��e��5_�l������'?
?���>$��>9��
����i�5��$�=М��ҙ>�v�~� �8��>MQ=�;�ә���>��=��&>�0>��R>�_�=Ԑ�=_ϟ>��=C��<��6����u����HI��E�����B��=�n�=�A=^�=�`��	�;�3���W����=A��<�[�>�|>������?G|�>t�h���X�eF��x�� ,���	>����pK�=��A�����>$>;뷽lٖ=�N��]?k�^C�����!��>#��>����|�g��==�Z>�y?Ck�>�&= �_>�5t�Q�|�4����Ž�G�>X%�>	�>Y��g��<�=�?���Y>m�N>HW>?�=�_>��=;��=䃾>�:]u��k�����b� ߉�P�:	�>>�A>�m>��=�b�b߾r����k-=*V�>��?�K�>U��$¾�,o���[˾�o�=t4{�L쫾)[�w�0>T��>2t;^Z���<�>
>�廽<��=����B��N�>`����>A`W>�&ӽ��]��ꏾW��=a�L>&�>aѩ>�	�>wd-?�#%?9��>�q��MfH��>G�|'>������>��?AB><}�>VQ#�w�!��{�������=�5��'R=��<x�=H�6>'�)�.�������P>>9^��6�>Ѿ=<�W���>[�d>���>�N<�Fm�8/��a@�X��w��׈�������\���=^�o=�Ơ��t�=t���?��3DI��t�1H>!�f>��=��o��Ϻ�������S=��������A6�H4���y�qIb>S�����<�$;۲߾	�h��ڙ�����w���U��m����a���>D�.>���=b?�=ܯn>��>�>Q>��=�+�> `v>�>��<��ػǡ>I�>8��>C�?uR>����Kn�Z`u�[�=�5k��B�=̎H>M%�=j�>��>Ÿ��C�����e�@��Zý�"=��=�&;=�>��r>{�I�re��<ξ�B��,{>����>��[;�p>]����,>�>Di;����l��[�sȌ>�:�=7~/>e/�>,�>4��>7�<ց���P�k==2��=�
>�T��޹�=9��l��$=��-�;+)��7����;��o!l��pq>��>�LH?D�,?��>��оg�1�P�_%�>%�׾����k�>��6>��>���61 �Y!�M����<VX7�a��;��=�&k>"�=l�9���\+���'���K�2(<+;S>"JJ>�	l>�O{>y��=�K���~Π��Tؿ,����<�3W��am���e����.�U�$>l�置=����:=86��K��>=�a��>���=U�W>�Q>h_-��F��R۳��tξj��D>+��_��f�=o�K����<������E4�;"��i���>�Ҽ�1���2�=��>��>�(�q
��.�н.��=E?1H�>��F=/�?�M�!~�(G�>����>��
>r6�>IF۽ќ��^��;g���Š[=T�6>? >>8H�=��`>��d�2F�='��gC'=pT � ]�'��~�-��Ь��">55>`T{>}t�>�����d��B���rB(����=ĥ<>���>z�þ��t>�h��Oc���=l[��)����*�\>ځ���<�|4P>j�⼿ �;��=z;żd)��<���\��� >��=�,>��w�2G�W��������=-W�=��>��>�]?�+L?;3?5��>���rK���@��ٞ>�頾��?Ga?���=yi�=��վ�@ξƍž5�{<�eW=WT�r{�= x�<���=�X�>"$h>\"�i;⽭(~>|el���(>~�<�V�=���>�x�>?�v>7��V�P�����޿��^���i���*�?>n�7;b��<�֪���<��<�z��L\J�O۾�"��ud�>!j�>FtR>�;�>�ݒ>���F>����}��?�y&���tؽ���>�,���7��PD�i8��ѽ��b�{)�������F�\.���e���V�>�ɜ>hne�62��u�1>G��>�M�>b�>b�Y=���:�~�<��%�ӻ�=��>�><z�>2 y<�a��]�4�齰�2���8>�b@<TlN=��=CH>�j�=�Ȣ;lzy=CnƽD����<�P��;pL<[>)4>�J5>�����Y�>O�_�W�߾����-��̮=x�@><��>��޾��>�7���ƾ�4>٫ɾ� >��D�D��.����>����>71>�o��b=Ǚݽ��b��A�>&������<��=�L+�b�[��`��̈/������ � �Ľd��>ϟ?>��o>7�
?�0?��?�s>DѾ�d=�s�p��=l� �f�><T�>NF<��=���'�@K�BA��꼒|�V��=�:?>]��k�^>f>S$?�C�r�H��=bi��bR>��9>�$>�z�>ۚ�>|�=����p�7�(�=�A���ÿ:=о�Ѿ�=l�U>Qt=��޽�?<])5�!��>�V�����|j>Dv�>b�?sOz>��>���>�̣��t���/O��E�����md��I�a] > |оsZ��a[þ;��?��=Ȍ��B���k"�#��l���;���v�>�Ȫ>�7�<ftB;��F>���=ė�>�>�k�>M��>}��=]>�;ӻ��=X�{>�C�>��?l�'>��w�w$��i
�Grl>$qP>l�E>�AD>4}���x���=' üT��<h_6=�=���#v�0=�=�[<>�i>ΤI>m�v>���='�>!���P�OY��E��q��>y�׾t=!=zo=��/9��a.��]g�ϡȽQ\�P�������Kb��)�>~�>��=���dl=��>�G���='?���I�XMT=�&𽵟������<�k-p��U����<`�@�>��?ߩ�>�.>�����WA���ܽ�A��I�f�a=5o>��==%B���8�tdξw�ҾC�ؾ�aI<���=��ڭ=A�=֦:=S/>C����>1E��:L��x>v6�=�y"> �W>R2>�g	>���u��;���׿�}�N�?�yF�=r0<?U��8�z�X�>��
?G(��?ž�s���>+�=�Q�?��<�4�>��>�j��q����D/=��ֽ�?v�i0���N���V��{큾��8�\�̽42;�^ȫ�Ы����D�>�Y�����|	�7����>�`>|�N�V��>�\?S �>�w*?ɀ�r
?��o����=��2>�	>@e�>�>u�>?��>���>�>ݵ���5ڽ?�!��=�qW<߅����=9=���<��t=-=����*�yJ;�{2=�'K<j�;��>�>�E�=����4b�k�D�W""� J��RK���>-ɞ�����.}��	�B�$!W��پq��nq���꾪3i�XS��xo�>�n>�<����"� ���_��=Ĳg�+j>��FE���:3�=�[�<}�� =N�v=�`�*i��zo����>(��>�
�>�[?=�<�Kᾬﰾ�̾���ę�><k���i =E�=��:ľ����{y�6Xz��ᓾ�Ԏ;g��N�> �0>e�>D�̽u7ѽ�S]�K/�=�0�>!�m�8�.����>^-�>^Fs��ӭ���6> ���Q">��"߿P��2��g���;�=���>���%�=�贽����"N$�.%N�œ�=�+>��>�?(C�>{m�>T̳�W�ɽ:b=%����"n�O�o�LP��]���0q��O�,<���=�˽�ND�)���re���ܽ�S��ۃ��%��?1�>�D�>qm�;Pl<Ak�>t��>D�>��<܄�>򌥽wd�=��!>�ж=FP�>s�>�Bu>��6>���=��E>�O���`�-�C�)�%=��F=+�E=��5>���_W=|oI���>�[j�T�Խg䂼z�$=|'=��=�U�=>i=v�m�EY����O=ɂ�=# Ⱦ�㻽�LǾ�h�>QȾP���뼭��흤��:����!�����7M��(5�=�>ȃ.>v��X�p�I`�=BE>�I��q��=��⼟����k;ɛ�gҝ>X&�=�CZ��hH<��=�랩<A"���8=�g�>v�i>ш>,��F�)�O3���x�Y<�;�=�u;���>���>>PF$������el���ѳ���=�=2�<Q~+=w�*����;�=��=>����T�=�h@=Xbe=��)>d	�pG=ԃռ_��=~�
�W�ǿ�L���來�4;� �uW=���<A{�D=�)<9���ԋp����<(�������<�=�(]>�B�>��>��� >g>֢��FᎾx���Τ�c|����A���+��G�|���OX(�Z�����Qy��3�C�>D7�>)��<��3�>P��>6?�0h��Ab>�p�p��>7�>��<zzz>:E\>���>���>�|�>��=�`E��eU�k��@G�ʊλ��ǽcJ>:1�2M=>��=�D�<[�K=����1�@P�mr�=�U�=Y�$=<� >�s�=1L�X��#�����0�4;��@��!!�>p����#��$辞+E��p�/� �z�޾@@����E������~�>�F�>��;�:�!u����ٽ������M=2���sӼ@_ؽX�����ý;_(�ؽ�s0��Q��L#���	�>��)?��>U��>���*���(�F!�:�D��W�ݑ�dM��0>�&�;�>���q�4�w(�R���Y?���=��=�2">�=���X�=����P<~*<��=�fl>��=��$>]��<@�=��!=,3�̭�����wɿ�	V���[���ü�6�=*�=�����=W>���i�L�ɒ��X�>:}�>J�>n�>��>ڴ�>��̾�w�	��q�}��l��"B��վ��Z�v�ǽ\
�q����#���~<��*���f2�;5@ѽ�C߽L8Q�RL�>|�*>��=	��>N?��?g�
?�⑾:��>�E=��>�D�>��>!u�>�y�<�Q�>��>3b�>���>�IT�R�(�B�ʼޢ<a��=��>�=���=�@�=Z�v='>�pF������=;i�=Ol=�I8<���>��==5
�h1Ǿ\�=bL+��yʾ�Vӽ_������>�����č>�e����}�I�?�������0�樽^	T�����6C>:g�>U>�l��F�-��j�D=�d��_�>�6۽p7� _>�-1���˽�/=<��1>��)<����I�=���41�=KE�>��>�\8?�y�=|�Ҿ��̾�)C�;���98.��!�<(�t>iWW�K ��؋�ⓤ�i��u~�GY�aND�V��=Wn=@B=�4>6��c�=K̽H��=�<�<��-�䨰=)4�=��Y>uG�=��>�/˼F�Y��� =��ڿ(��������پЋE��=+��}���������,�@1�[D��������޻	\�=�7=���=G�>8c>������'Y;�S �i�����ކ��K�
��B6��$��GF�����И�~�x�C�3�<ie�Z�꽅���h ��p�>�%�>���S]8�1�U>d��>�+�>�����>�ԽJ>��r=��>䅼>Z��=!�H>Ʋ>�i>Ԣ���u�Zt����+=�G�;,yh=n�=��>�@6�;hN=.�<���<}F�4-�=�8u��q��ь��f[>��=��=��>NK|=Nǃ�P������@��~�>Sֿ<=M�	��>.z���=2��	�T��Ҿ�6����K��->I�>i>�	���Z �� U=�>��
�	>ɸO��2�|S�<��>F�^>�<s<��<r��cq�;�`=Ou�=�=A�=+�?�O�>fF�>����s��a���B%�S�= 1�����=���>1���U>+a4=.|��7Ⱦ7�t��@��%��>T�>^O��j�>k�Z�k_$�� ?^s���:E����3�m>��4<��>�j�>̇">�m�<�ɾ�E��r��ÿ�ﾉ��+-�.m��� Ž����ﾹR���#���;"I�=<��;���<n�T>��y=�O>��=�گ��N��dOC=�������S1����z�n����#��=�Wh�0^F�k�.��7,����.��wd�4�=�[���^�>Hý=��U���e>��?2~�>�g�T�>p��=Nf=�K	?#A彮B�>/k=,��>lo�>�L?�7�>�8ֻ5ڽ �`��M�=��r>A��uNW>��<=�A򽖼C>��9=MG�b�b�'�=�8������o����$�;��R>�(>[��>3��=]"��jB��u̾i�#=uι>�>�����>�h��F�"������B���#��������~�>�b�>��=��������qa=��=*x�<���vȔ=��J>�N߻׭'���+�B����*�q�>�ԜL��Tɽq�C>{�=M??�9?��?	�1=�E&�'F"��<ɾs��=��8���=���\>DZ1�^轳���n�ҽX�,��]���\��a�=q�\>�8>3Fm=�I���꽘��=7�>,�2�~�[=��+���j>�=>=4l>M��<�l&>�+.��q]����>%ݿ��y��C�羸b���ۍ�?~���Ҿ����+��,s�	R-�G���(e?=vH>�'�<im�=�ʒ<�<�� i�γ>�ȉ���ù�l�1�S�����(�ͯ��i�=�l����=����t���l����ɾƢ��=~>t�<=;/H>y��>C}?3R!?
!�>O�6>3�>��1<Nz?�X> g�>���>�?] 0?��?�R�>/n��~��֊���>j�>���<J�=-P�=�k5����_���
�=�L>��=ۻ��̾���[ѻ�?>N~�>�� >��>NK|=Nǃ�P������@��~�>Sֿ<=M�	��>.z���=2��	�T��Ҿ�6����K��->I�>i>�	���Z �� U=�>��
�	>ɸO��2�|S�<��>F�^>�<s<��<r��cq�;�`=Ou�=�=A�=+�?�O�>fF�>����s��a���B%�S�= 1�����=���>1���U>+a4=.|��7Ⱦ7�t��@��%��>T�>^O��j�>k�Z�k_$�� ?^s���:E����3�m>��4<��>�j�>̇">�m�<�ɾ�E��r��ÿ�ﾉ��+-�.m��� Ž����ﾹR���#���;"I�=<��;���<n�T>��y=�O>��=�گ��N��dOC=�������S1����z�n����#��=�Wh�0^F�k�.��7,����.��wd�4�=�[���^�>Hý=��U���e>��?2~�>�g�T�>p��=Nf=�K	?#A彮B�>/k=,��>lo�>�L?�7�>�8ֻ5ڽ �`��M�=��r>A��uNW>��<=�A򽖼C>��9=MG�b�b�'�=�8������o����$�;��R>�(>t��>���=j�羋B"�8���������+>(:�Oz$?�����N�)����ܾ:�>hN�S/�O��p�4'�>�\L=U��"hc�r=n>���=��!=������;f`�=�r=�$>7�v�#=�9��=[��<��0=�I=��v�P>v	?~�G?s��>����t	�����{��m�=���I�=I�p>�Z���|u=AG����;���x�������Z��8X�>t>���<�ѽ���|Nw�,�c>I�?>�gZ=�eu�Uc9>�v>��q>�	�>�)�=X�*��>ּ8˾����ƿ����Q�7�V�$�4C�h콾n�ƾ`�ľO�̾Q
��(�<�lL>Oj+�=�<��.>��>�>�[���4S�RU+=�����F������y�ݽ2g���!�0�9"k� � ��F�_z�={�V�����;�w������=ݼ�>��=�c�=��>-�>��?�C�>�%�=���>g���;��>8Ơ=���>��K>O��>�í>X'
?i�>0zZ;q}"�{)��=�=�z�=����W=���=9�4�.�V�_(���x�<'AN����<����}!�V�#�<i=�@�=f �=Z0b>|o���yҾ��ž4����SK�h��=+}�>�r��n�;eZþ}�)�D�s��'�����O�ǖ�^WQ>���>�>�	>��_���ܽTM����lԏ���
>�8�Q,Ҽ-��xŽ�����Ѫ)��Hܽ#⽛�|=ٟ�="��s�?��Y?l�Q? ��r"㾪4
��=��>jJ>Ky,>i<�>�.�=��?�����������<V�Z���ܾ�o���UW>�FH>[w1>�> <C��̚��Z�=��#�"�j>�U�=bv�-Z=�=}.>O����휽�[P��տ�*�����U ���X�4��(ٻ=�����־^$1��&�����~�]�nŔ��6˽�v�=Ik<�u���1>�oy�!U�<m}�=a[�;.0�[�¾[�X��fN�!㜾��>�Fྦ���wr�&��N��S���1����uv�,���o>�T;Gl�<��A=�&?���>�8>�>�nW>��K�葿>�'���p>H��>�,?0�> T�>:k?�s`������{���1`=�*��آ6���
>�s{>/�
z�=J��=��[��H�=�f�=XU>��:>I-&>��>H=p�R�iV�>m{�=|��������h���� ���D�>�j�<�5j�;�H����2�����J���N>�pl�d�ھ?��>%c>�0�=�^�?��<0��=d�X=ٰ��y$$���=�:J=W5h���3�H�|=r�=��Y��="7S��(�=N�I>w�=��>܃;?'"%?�l�y� ����@���d�I��= �>�pɽӒ=�]>��e�Y�߾ 2k�K��=���Z]=�F�;^3>�a0>1�2��T=���<���=�=�t>�[�>�I�>�w�>���>��>Ղ=>�1F��ѧ��- �sȫ�������0�}���������zn ��	e=ݻU�����F���>?>�����4���
�z=J��=��>�lt>�"3>�Պ�=�6�w�ƾ�G׾��=�j�����4ҽӒ-��i����7ل����ܾ��۾�K��:�>i�=�D��u�>&?c%?C��>���=�>�=`�>~�> U�>�)�>���>?��&>p�>�?/�B>�QE��rR�J𼙮��.=�V�= �:>g��=*&K=��ټc���e �$O6��u����=%�<M��=]ӈ=+=�*�>0&�>��:� �=���?�&��}����rI?č�my�����8�"��G���	p>Hɾ��{���\�>�Bj>����i�dܐ=��
���;>���=z�r��v�q06��9>�y�;̔�r�:��!c��E ���>�Qu>YnT>yy?w;?�??�)��`�r��&���FV�\Mm>��>χ�<֪�>�V>��ؾo����,!��^�g�����X>G�n<N��=���>���\���\O7���?�G>q:>֧�=_��=[ ?��>C�>�ڤ=�bY�|ξe���7�Ϳ#B��CY �!ċ���
�߆V�?��4Z��f�
���5�(�þP羥Y=�6>�K >�C>�tZ>Ǚ�>�թ��Ҁ���o�FO��%�9} �/�Ǽ-K���^����=9�B��p������_����,4�ys<�' Ƚ���>�SM=���>���>�@?�38?.�?|z9��`�>l��>�o>b��>�7?>O��>P�=uC ?��?�Ҁ>�1��'D�0ߊ=��m=Y ���)>�Wp>�X�<�(V�M��:��1~Ͻ�i���[���Լ'Sݼ֏>tg�=���=M��>�z>��X^��L�<E_�^Gw��#?���,�`=TܾU�@�Enj�3�־����t[>�}�,J��_���n+f>VWN=P����=7�a���
��p�>C�'=�����!�)=�3=u
���)����o���Ԕ;h�>t��>�f>E�>wO?��=?�d)��*����9>��=�<F����>�=e��Y�J:����%��� �����~��;W���m>?1t�E�����>v��j��>6;=H��>�y�=�D�=�W�<��>�B�>���>?�b>��W>᭾__˾�4�n�K���05��R��uȽ��H=]ƽ|ž[�^���0�]~����r�H|>��)>�Ev>Lݎ=�~=^����Ϙ��1=��=u�������_�?��;2�����b>^L6�?@ܽ}ʽ'Y&�T�
�\����p�p�0�Ď!�D�>j�s>�%j>G�>o�>?k.�>ﶸ> �����?��O>(��>��>HH	?奕>�>DV�=�`�>!�2?�-�>1��}����=��<>��H>�Ӄ>o(z>&e���;�:R�=������ʽ}�ӽ��]=f{�=]�?�O�<c�=���>�Q�=����t����=1/���"	?m̻��e-�4��(۾����~ž�X>d������$=�1�>q]=F�r=��s=�Cz�H�M�,�>�Y���v���4>��>��=�T>FOh�5���|C�=H�2�x�)>Cq=�>cV ?b??B<��%eG�f�����RX�ن�>��>�<�>�4{>������h��5徶>��V��j�G>$M���W�=Ȋ�>i�{=n�={�{>Q|�>ɮ���)S>o[=��<L�>�d?��m=^��>I���t�# ���Ŀ/��8y�����8>�~>�'w=�����������&��bM >H��>*��<܎�=v�=t6�=$������=&��-ž��������%��=�:���a>(�ͽB���T��Aֺ���D��	��8�!�N��[�ܽc�@>6;�=��Q>�a�>�-?]>��>�.��~>U�"=�C�>:��>���>���>3e�>�Ǟ�C?r*?��q>��ٽ*�g����<�M�=쟺=�ul>�t=��Ǽ%�=�,��H0��0���n��l�*;�m=f;;<B���.-<,�&>���>�Q�=����t����=1/���"	?m̻��e-�4��(۾����~ž�X>d������$=�1�>q]=F�r=��s=�Cz�H�M�,�>�Y���v���4>��>��=�T>FOh�5���|C�=H�2�x�)>Cq=�>cV ?b??B<��%eG�f�����RX�ن�>��>�<�>�4{>������h��5徶>��V��j�G>$M���W�=Ȋ�>i�{=n�={�{>Q|�>ɮ���)S>o[=��<L�>�d?��m=^��>I���t�# ���Ŀ/��8y�����8>�~>�'w=�����������&��bM >H��>*��<܎�=v�=t6�=$������=&��-ž��������%��=�:���a>(�ͽB���T��Aֺ���D��	��8�!�N��[�ܽc�@>6;�=��Q>�a�>�-?]>��>�.��~>U�"=�C�>:��>���>���>3e�>�Ǟ�C?r*?��q>��ٽ*�g����<�M�=쟺=�ul>�t=��Ǽ%�=�,��H0��0���n��l�*;�m=f;;<B���.-<,�&>�h�>͉��Խ0�C��ԙ�= /r>�=>��> �<��k˽���<�Oi�6[�H}��5k�y����꽗��>5]�>ڿ�=<�U�=�}t=�a=ў�í��獮=�5y���=)"9z O=�q>�?�=.C��K]�pA>��.>��<�>��?��(?��>7B�}� � �3��r�`�&��>�X>��[>�R1�W�R��%˾ai�cC���>�`)��. =o�1>7����Ć=*->
��������4=��_���9���S=�n�<�����.>��>�;�M`��J�F�
���cG�������,��(� �����]�.�-->�?��OǼ^�ۼ�z������O��b�>m:O��l�>h���۾�h\=B�fI�$ɯ�}�Q�a3��\'0����G���F[�\�=��\l�&	�#sg��b�����e�B�{x���O;�>O�
>�%����ӽm0m>�!�>���> ��>��>V�C��Pҽ0>��V1A>���>�>?(�>�C�>δ�2ν�O�����%=V��@=:7�>+=>JRJ�"1�=9X=�>w��<��>������"P>�s:��$>�,e>=��>��_=�ܼ����"=��<���@v�>���<e½��̽����Ӿ���`A�=�A�$o���Y�>,A>�{>;�=~�T=y�<����E��2(���=_�>S��G-��Q�<ᨛ��y�<��?>� L���k��=�ûԒP>h�?6q�>^��>::������#��v�􈬾Wr#<��7>"t�>�蚽(=�=0?�M���ؽx+վ��Ծ�eܼ�O�=Bt�=<��=m*T>'�d>��<Cd꽎}l��ȏ� �c=E��^� ��=m{���S>%>�Ģ��č�S��S|ۿ���L��)��j�=�>r��>��h>�9x�����b쮾\��|�4=�tm>��>ʍ�>n*�>��F� �8~�=&��Tn��Z¾�Xξ�5��UX=��ŗp=����t��z?�ڦB��/S��u�<��/�/v��D�� �>��p>ѽ�̉>�y�>o6�>�,?Nq���V�=^�B>���='�	=g��>�'>�CN>�?���=38D��Zh>��k�UhA��Q��ؚ<��h=��?=w�<Ū<c�=i�W>[�h>�p�= >!�+=�'[=���<W4*=�qZ>�}y>���>�b�=cs�=�RQ��/R�c�������� �>��s���N<��>�h%>��ؾ�.�+I=���!ё��`>�`�>�	u>�30>��}��-ܽ�S$�'�ӽZ�����=媻]�"��S׼�)�=��j�\U������Ҽ���w�< R�:�H>X?S:"?�
�>͏u�}x羫3#��#��R�P>�=��>Q��=^�;�����W��ñ�����54޾M���J�;�э=��=�aX>m��>��>���=L�{=�沽+$�Z^��j-��4T=0�=d�E�7m;=��>�ɽ�􂽎��Bݿe�l��}N�~�����=�[>Q��={wP���ѽ����Tk¾���>ǵ?��=�+>f}|=�/I>��>eѥ���˽ڶ�fJL�b�ᾘ%��?l���QW��&(>C�O�gPｦ�&��a�61f�����l_n��M�}���f�>L�"=�3���>�z�>���>��? �u>�&?�r���
�/᤽0|�=/�t>WO�>�]�>iF�>[K>cy��ω���'�AM��\�A�6r<5>2=<�=F���H6>i��=��=�>Ez=,%�=���=X�<�=�=�>u,
>=��=�κ��%"�Pc������nE�ޒ�q3C>�y	�ŋ�9���+��Q߾=�l��C��x<���������c=�	�>�=�F�����A����<�o7=T��]�+<1n�=��=��>��ɼN>�ˆ>QF�Q��=S�M=�-4�#�>0�?Z�*?p��>�X��ϧ�8n������[���E�=2��=ƠV��S�>�ɶ��:ξ֨$������¾���<���=�h>y|+>��<q˒=�,�=|d=�����;��~�>nxf=8���:=d�/� ��<���<�W� �ѿ��.���3��v����
���=F��}���'��y���(=������5�<e�>��>��z>Gy�>jA�>Qq�����=\�v�~ؾ�举�����(���:��=�o5�g�1���>��G��匾[}���m��{���U�xX�>��ݺ-ت�
 X=��j>
��>��?6�>��?% =S�>f0>���=hr�>4@?>��>��>2��>ms>�h���>�K��<��K=���=(x�=_-�MKR;/R=!d<��;n򻰻����潹�Z=��; �?=Є�<n�>Q�>=����=�<�B5�WX�=�>��G><͗=�D׽�Ȃ� �k�S�qѾ	����t��l���/>�ǘ>��>L�T==�]�bZ�闩�6#��C:��C=��=�oi=��	b>�u=��=e���k�`=�=xji>�lL���^>�?L:?鉍>,y��l_�+�'��
�6*����>⎟=�T�=[�>���<0�vh��-g��־9���{7<��=l?K�[�>�g>���=��>�2v=� ���67����<3f��Ǵ5>;����<n~�=�M> ~�~�&�7k��=ƿ	��X�2��Q��R�a�jM���ŵ��
�=��	�^9[�����1�I���6A�M�;��g����=�р>u�ξ��ɽ�<�;H�����m�E�-�f�b�C�o�]B�=�A�᛽�O]�
����4νY��پ7π�l"Ľ�©>�Gt=u"����4���>.,�>3��>oX�>�ߟ>�����@>�>�]�>(��>�X?��	?���>�%0>�L��0��m�ؽ��E=�(>c=����:� 淼�fؼ��>J�6���~=���<����xC@=?΃=����/@	�9�
=D%I>ȡ�>�[D�Cf>n^?=��9��4>6y�hR�>����R��ϼgq�׮�=��˾d`��?\P��^�>�P=�&y>�>�x�����=}T��/�e9R�[;b>�̑=𢷽���<f.>��=>��=1s���Ϩ>��4;����E�|�\�B>B?5[�>�?,?��� �+�x�	��hw�M���*�>�C_=1��G�>�=��V����i��"޾�Y�< @�=��E>�ʘ=�-�=	�Q�:��9�ؽ.�2=Z=�=0z��n<�|S;}0>�� =���HQ>��'��4�x��m�ٿ>zb��r��Y	����=5��>&l��E�˾�(�]��l#�L�T��i�>�?>�uľ�=�����*>W����� �N�����<�um�"a���"��P3;�E������ �������K���+����
��/�(���]��>���>�E�=�k�=l�	?��>�Q�>5{d>��>�<_=b*"�=s�>.b$>.<���p>�����>0)�>�E>�!��vԽm�x��|��v�w=��>#�!>^�x��*;kt=|ו=�"�Ib��˭��=Ǌ�9�Ľ�Q�=��:>f��=����/��,�@=+"�`1Q�������>q][�q�i=_�H>w���Gݾ��>�Ǝ�1~��i>��>7� =�f9>U��=u����3�
�>�@>�6<���=����`�g,=��:AI>�q�>��:�ث=�쌽|�=�D=>"�#>���>?�6?�&�=�*b����Θ+�R3%>P��=M�_=j"���8��1w�;
m��>X�uf�ť�� �8�Q='�t>/��=n僽,e=*F�%ʽ=iH��߈=��=�ŧ����<��=�>�<��<	.@>^	>�	1=�S��M����ƿ��4��tU�8��bY��ׄ�?M����6� �>�kY�  �>|w>grl�-H�>�p:�mߗ�<*��(И�������	�n	�<�-�Ϛ��Oƾ]�6�1���5<7=�=�v��9����<����,�<�&������ ��U���T�>���>�"<_��?�#?�,�>�~�>�F>5ǋ�]<��g_�ȍ�>]�>���->��H>�d�=L>�=,�N>35M�*���!=��(>�� �=�]=�\=������(=Tl"=�l�=�<����'�>�,ܼ4�*���Z��ut�=4�#=���\�<?�V>+��L�k�CG���+�=��>S�z>�q��I�H���a1Ҿ��>ƀ>2��QH!=8��>?��>�k��� ,�t�=s���ܶ����>�_s�|=����>-ע=���73�����=6�>=A��o=>��$=	��>;��>��)?�'?�Խ����O�[����c�*��~>�.>�<�h�=�p�=��ž����O�w���˾�9�!�~��h(�i+�>�>#�d����;�*����*�>������7>�v�>6D%=|�м]C�<��>�j�Ʈ��>����¿�B�v�=� ��2˽�f�щ2��t-=��=�X&����>�q�>�"i>������<`��v�����X��V�w�G��*��\���������=�����0��=�v��,���L�	=/�*�`�f��Yʽ�h)��Q}�~�>�s�>p�'�5I����>/e
>J��>���>�G���x���"�>l(>d���U�=VD�>D�=}��� �>c��=0���S�̽��F<�R���=���<��=A4���P >��=vb�=�V=������ʼ|㻸_�!�=
�(���=�
�>-r�&+񼙢k>s9:�*cԽ%�R��=�+=ر>Ǘ<����hJ���9⾥�&=��>���=AN�=X2)�<�B>1�[>�=�}��� ]=GS]>����gk�>��<u��=�k�=��=�>Y>����8e���c}�u�w<sS�<2�A>��>��>���>�v?�S�=�2�l�M��Y���y"����=���>�	�>�%�����zd���u��G#�w����#�a��;�Y�<o���1
��2��w�=�yP��&= �x:�>G��Y��RT>�B�=I�I>�[�=;S���ѽ:����ϿS�fbJ������M�l�W�|��l�$�������+�=�Js� �=V�8=/�>=��>��> s'=옍�� ��;�;�=����d��	n<���M��ʽ�V[��5� �&��"�k����Յ��y��V��'ƽ�N���J�>�� ?2>��9Zҽ�'?u�^>
,>wq>L�m>��ܽ��ͽ�D�=�)�>.�>
b4>�d;R>h<Xو�a&>�骼>�˽��}<<8i>u��=��e�4�T>_�<�C�)�L�9����UT<��W���?�`�p:3�;/�ְ�=�N����A>��*���O�Pn�>|�#��kξ�kW�*3�>�!=�Z>>]������X����U>�')����=�>0R�>�T�����>#�=luH=�z8����WJ�<x�?=�P�>�|�<G�1�����a>k87>ӫ�=jD̼�mc>��<�,)>g+$>^>�}&?�C?��>�"�>#�<3OT����:)˾���>�6�>�P���>������4�(���~����KI>گ���>�(>2��=~�ںsԽ�Ur=߾X��Jt9�Ss>�E�G��-RZ��>��.>FM=��>&�(�
-��
�ԒտU����{��虾H�ü?5>�C�W�M�?a��y�=��2<ƭ	���J����W2(�u��=!���w�����=��8<7���.�=i�پﶜ�m�˽;c_�4�g�������ڽĠ����q��:�'����:�B���߽��>�_�>h�>��K���!�f�>�v>��#>\�!>bMb>�]�	�B=�7>S=��0��'�>��[>´-���k���=H�U=B�����h�<ʨ>�	�=7�q� ��b=�&��Pl>����P/=M�@�Y�����
��a�@o�<1R>~[7=JA�KGƾT\���U�J^���>u���3|�����vZ��ϴ�K�����=�L��G��zi�����;��>�a�=�&�Df<�O>1��&軰�(=�X��^����v��=�R>�>cr*��T"�s��Dp\=����A�>�[�>���>+S?}�K�Bu���$��S���Y.�H3>E뭽$" ;��ڻ|��b��+ξ2��m��t�%���_���	>Ʒ�=駂�ԑT>�'����;�4�ߎ�>%�߼�������;2=�/p>���>���>�>G��>����@ҿ�����F�Y�Ž��l��3��[��ٻ?��t2��`�B(g>��>�=@�۾/ɠ=�tZ=D�=Ϭk=dg�`�>��������:�޾���T�>�<j>�J�-���G�(���G6���#��}��.���ҽ�Ge��!z�0�x�Le�>�\�>G��=���>���=Nk�>I�>�b>ز�>�=m�>hg�=/>�2 >��=���>�<�>��>��>�$�OLI�q��=�ʼ9�֢�6B=%�=f�w=F"�:�m�=۴=d�ȼ�I������N'�P=���=	!"=���=���=j�ؼm7���W�� ����<�6��[3�>��\���"=a��uA�����3z=&D?�H*U��i�Ī%����oR�>�/�Ϟ�-r��la>#E>w�:>%T��=�j�eȽ���>�Կ'�9T����_�K�=I��E�>�x��Z�=���>�-/?|�?_�=!��`�	�#��X�������=���>9��JѽC>�ɲ�TL��oQ��Q`(�-���»�>1�Q>2��=��;��N���.�v>K��Z=Z�x�
�B��U>)��>��>��r>��1�L>L�o�x��%�￾[�� g�r���3��/c�<L��=
�1�vcD�)�f=�ӽq���-1�������!��黒&��4ͽ��>��>�|6����=����Xؾ�I��$�<�ʗ���;0ڡ��?�k�Ⱥ��= �� ��𛖾�z��ۆ����>Th�=_i3=��=�=���=�D�>$ˏ��1�>����,�>�߽`&�>��<'��=��>p�<>Ef�>��e>��w��C(�DU>�Z�='�U��M�e��<�a=� e=j&�=sp��$8<��1ӽ�, >�8|=)��=3k�<�6�=D)g>c˽N�������J��H	��,Gƽɾ�>��Ѿ�4>�v����6�����˙��W�Z.���O��o'���þyG�>5��=�*�;�����^>k暻���<��]��#���:)=��_���=P�����h��d*">O�=L��=%V�A^~>���>�{?��>J%ཿ�'�d���Ǿ�Ԭ�4>�Ĥ=���=F��>��H�`K>&����ܾ��5����;޻6�c>� *�S�<��h=6[>��(�Y�P<�!�=n�����=�s��;~>�/K>x=���5=>�'<���0
�=����ʿ�� ���=��0�w�PȾ��ٽ8�ؽ��������k+�P�3�	�&>nǽ{�X���ڻ��q>>������
_9��Q����r����#9 > �5��;�����o��B-�y���'k�:�����˾���C�b��.�>T�2>K�=�w
>I[�>���>[�?2d:�\�>^m���M�>m��=�G���A>��;<��	?�t?�Ͻ>�Ñ>���&]���=��j=���-�A=�p>�}�=]�>e��<��<9��<�K�(�?:�� >CV>��i=ϡ�=*�=>]a=	����r�zW��'���<��:�_�Z;�9��S%�= 6�=;�o����QV>8n�<~cؾ�G�<Y�=�%�=��>��)=��꽀�s�܆�=���犋��`�=��۾HmF<���<�6=N颽�'>���noF>�����Vi=��b���4>��>E� ?��?���=�-(����8M�����T|>]�@>>1s>]�>O$,���>�'Ҿ₂�u���e=8'���K>]�>�ݼ!6��"�=�����pU>w�>>�j<��E���>K>U�=s�0�>]���m/��K3;��������,¿���ͷA�����ٗ�m:���ȼvu�����K�Sھ�ҟ�\H>})?>8,�>"��=
�����<��/>�Q�2�;5>`վ-����侙�'��#���:��*��ۆ�L뜼� 0��A�����v�ؾ�҉�)ow���>*�l>m�W��.����=�8'>��?k�>��>}�g�cմ���=Vl>�Ξ���Z�2��>�>�f�>/��e�A����M�<N�%����=�v<��>���L>�>Y�=h���l���U��#��XG�#V�>��b=�U>�D�>1�x�_���RP����
���1'�P,�>j����H�ƿ���σ��vi��oE��*�Ժ�~ھ�ߠ��D׾��=!O�����=� <�6k>!���f�=Srٽ{t>�<e��v��&9:>j�����=��'�<�u�(`�=��<��>tUA?&?V�>�Yؽ�p�Y�#�n�)��>Z=Rع=͝�>�;�u�����y۽c߾�V >�����r�>�D$��8�;OP)>h,>������2>�L��d[�==� >�$	>]$9>?K>�輼2�G>1�$��l=<���Fɿ�{ �T��G��Q���H_�b? ��g{�"���.z��m���A�ؼ̐[>ݟ�=S�\>��_>�ԧ>�G>C��>똊>��|���T�9�9�YĔ�i1��N�>���I�V���<x$��5CN���ν��A��Ř�����r��Ń7�3͝>�.�>Z������<E��>��>���>�ؠ�>?	?��I�S�>��q>y�ɽv�<>���=r2�>���>��>?�>�N���O��ύ=-���"�}��佹�S>ӱb=�>��y=p���i��Ǫ;ZU���C�<�Z�=d!>���=�IY=��>}��K�װ�jc���G�t\��r��>�~���
��J[�>U���\���=7���9�T| ���k>�(��(`�>��s>�f|�)�7�j�E�^�>����;��w�ϰ���6��
>��%<��=�	��pվ;�_C>182>� L>·�>~��>��>�
�>�P%�dl������ؖT�7S>xX>�,���/>�`O=������N敾nZ�����<�~���ýɉ5>w(~>e7&>��@�����D�ڀ�>��~>^^>�<����א!���>�a�>?�I=9*a�qʾ�G�*ݿ�lH��^��ֽ �>ec����Ӵ!>gLվ��p��r�:��=d�M=�i=v!ƾ}d��^�W>��b>X�=cb�=�=��5�.Q��(�Q�wa���T��D�=��>�2J��FA����F���^M������Y�<����>��>'C�=��S>J��>n�>h@>JH	���5>����`=�o>��>x����>_�>�a�>��=�!>��P�Rh���O=E��[n��U���xy>�>g�B��������=ћ=�t�=�@��R�����%���=��P=�;%���������� �-����F���t?Oо���ε>��o���>���M�$��.[���>4o>U��z�>D�>���<�Gֽ�(��$� ����<7�8>	D<ؗ�=��n>����w���$���N[|�)��<&�a���)�G�>�7�>K9�>�L?B!:?d>��8�S����賾�A��O��$>1š���>�>���)��ؾ������瘈����='�8>; ��$>�ґ=��龠���Õ�=ؘ>x=�=9&�����>+��<�^�=��>/�;\O>��J���
���ȿn�|�SUP�i�-��=�͝�7��X����>�¾�w����<>D�j������:���l�_>"̾K�X��q��t�s��W��/�ۆ��h!�u|1�jsl��k�����=u�>���=K����T�V�@>��߼[r���>�8�>7�@>�1�>XS�>��U>��>�R���>��X��T8��p�=�1���	�=���>1�=�>=W8 >�V{>\F����/��l�;�D�=*>�C�=��n>@��=<��:W�u�w���{��=�v<�{4;���<4��0�.�癬��;F��H�=tg��w¾zm����`��3jU��?"����M=��8�a���Ӿ�}�������)���ܽH��=g[d��(�>F�0>�Ք=c��;�J@�N�]�,Kټ�,=�W���_�3+�=�">B˜�^,�<T2�;X����M�z�=�$����>���>��?�?�^c�T�ƾ� �P.Ⱦ�'潅��RY >�y���/&>!��>5|Q�b�������2��;ʾPֱ����=Տ�<���<�1`>��=8Ǘ��H����;>=.ý�?�;KH�.��>]n�=$t��Q>=�>[-M�1��������οV4~�� ߾��>k���X�������T>�"��`o=��x)=��=�������qI?�[?�2-=�KP>E�ʾ�Tj��/���>�z\��֟���~�;LF�[~�����h4��/�'̾�*�Y2!���׽g�ٽ�ZȽQu�>�xX>�i�=�;={��>���>�S?7
�=�ӊ>q�q>`n1>Y<,>�AG=?��S!�>!��>o�^>�Y�>Ѕ�>��[�Joʽם�;=w�<�Ɠ�1��<ǰ>,�=��=��=<�-���7�qTE��E�Gy�=DbƼm�m��>�Z>������7����;���P���ea[�0V�>	V{�x�s�p���x��EF����=½�D຾���<쐳��=���>@�>_�k>��>m@���Z��{���cb7�x���3��=���=��輅Y�����������I?<�O�=uh-=�\�=Vс>ά�>pf?F$?	d=�ž;�mľX+_�W-C����>_,ɽ��=�%��M �l-���꾾y��𱾥(�=,F>3Խ���6c�=ՠ�=�G��Ѳ"�
��jK��4�<G�5>Xv�>�C.>�m>�(>p~���9u��RT�	�������@P����:�=���=?O>:��=��>~�z��5�@>��_>3��>9K��1ɾA��>tE#>�n�>�`.��Z��\Hƾ,0�������7N�(���u�����="U-�ã��Z�6���=m�������v����-Ƚ�j����>TR�>�b>bd��1i�>���>�U�>����=���>ܜ8>�9>>;z[��j>4��> �7>�j�>�"�=���E��n<z6�=�=`s�;J\�=�>��=gT={��W=�DЏ�Z����:6=��p�o�̷>-��=��>>9�؂��t���ݾ��>k>��ٽv�ξd"��OE�򶴼�~���l>YH<7	������u�������>�>ꏼ<�'=^�<3�<�΂����<�c3�������z;B��rҽ\;�>ѧ�j��q��~�ʾ�M���?a>�X�>��E?j�X?s�@>�M'��I�=/���F�Z���?2
�>ha�t�q>��<��E�Ծ_a�iq�[)`�h�{>�=�k3����=�/�=�d۽&LŽ���=�2�=��<44~=c��> ��=�o�ĉc>r��>�/�=U�#�~��B�%�4��6꾴���6�'F=��5���>e!?�B��W��#�׾`hֽ����Tlf���>�+x>��>��þ1�E���l�5���B�������As���k����<3 �>�ɂ��E<�U������2��8���C�s����H�e>7��>t�<;�z��Xr>����&�9�t�>f�>���=�\���2j>�Ug���>M	?C��>���>2��>!	��=
�hA=?��<=#=K<��>���=�==��=3cλ@�t<��ü� 2�+(,>c�=G�g�e�>`��=B��>2�%>��>�Z�=>�྆א=�"f�@)s>z�y>	`d����=:� �L���%��w7�<���>{%>������.>~>j������>�>v򾽚�T���=n&M�S��=�Q�=�ս�?=)�-�?2>���<���>+X�>.��>�r?!?��c?m��>�ܾ`�X=h�(�����y�>e��=�=߇��ژ�����z�	{���6�EľZ��+[��� �>0�>�J�<�:D<����H-=�ܨ=.|���6OԽ|�=E=Տk>a��T �-辰1��A?���]ҿ�!�qF�:
��8��DТ=�f��/�����>���g*�z;���>�L>������6Ծc%f��x>a?��>F/�!�缁�˾v�������:>�xƽ=(�{��6i2������G��x9��N7=�>9�;�R���>��>�á�F�Ѿ�_W>���>hr�=M��>��9����ɒ����>Te�>�ɤ>�U�>['ʽjs�=2?��>��"��Uʂ�S��;G�y=��H8�>ڑ���X�9�">R���X�=6�<�Nh��j�;�mc˽�ֽ:�=hʸ>�2=I6=n*��־�vP�R����>�\��-[�>����9ێ�#�%�hb��pU=l�>O�伡?|� )]��L/>A��<�	Q�#b��#�>�?�=�_�=�v�;�+�}��<��=��>8<�;>��~5ּ��=@�e>F�]>�wm>��	?���>��!?g��� s���	�������==�	�g�>�A��zH��Z��F����gg�4����<���|�OA?�D��h�9>�U>N@W��߽#����c9>�#�=C�u��4=Α1��F�����#>K>��=��S�E�u�Գ�sqɿB Ǿ���mO���v�w�k>�c>N�>A/=rrt�f��G9>�٣=@R2>���=�>�>�#�="�O�;�<1�)���U�o^񾆳m�4�������A ��!��e����_��V�LQ&��qn�c &���*��/�����	w>��4>\��+P����>�M>}B�>j؍=G��=�ᔾ��>v^�>�H;>��>��/<�3��:Z<~��>wny>{���0<��>��|=D�,=,&=�>X��K>S
=Ra?��Oy�fJ=�>ڽ�q�<�$�㹦�ۥ9���=�S�>�{�=��<�Eo���[9�������*�>�s��XE8>=���籾cv-����ܫ�=O *>�[��+�0 ��P>��>�Z��w8�9-�=
��=D�=y�6>:�</�9=�*���=.���9�Z�?t�=�#�<�Z<��>��>��^>:O�>D�>E4G?4m;hZɾʹ��Y��5tֽ�w���M�>��_��e�`��=�ھ͆�|Z��d4ӾP*6�h1���u��Ϩe>y::>\��=���j���BV�8��<�L���>�[
�
Q��'���D��<�)�=c$\>����b.�kl���ٿAf־�_(�S$1�p���C>��Q<Yyм�F�=$쑾��*����<��=�Ǽ���=��&>��=���>vI ��P�=��f�H�5���۾H��������=�q2��#(��l ���H��U�nu��c���B��m�W��@��}�;����>re�>4O�����?5�>�T�>,N�=!�>�z����<�'�>8�A=z`>�d<>��F�n+Z=���>X��>Z:��;\6�/炼���=�j<QQ{=��>�h���<R~9pƨ=ؑ=�ƭ=֞ >�'.��"d���������K>��S>���=M�0>��}��ׄ����B���>�]�=t�4>8�Ծ�!$���)�s'p�T����M�>k˼�e�W�w�q>�� >z��#�]�>KV>�F�==G=���'<����&>`�q>��Z=w�S��]���;�IYt����>"|�>Q�p>��>�y�>Q�]?�a0=����L�c�Ԫ�ڏ�<
HI��߂>����;"�R��=��ƾVO����@��9��g{�tp*�
G׼��>)bf>Y
%�o^ֹ�*��aV=������������i%��Q>l.}>F�>!
��cL�=)�����r	�A�ؿė��;h���ջ�Rb=��>��)�Xz���ǡ��?���;��H�=<y>�7�= g�;ߤ-�b�{��=>�r�̼��lƼ$��C�@	�Δʾ�=ҽ���
	D>$�b����;�ľ����bT=*N��ATl������o���?�>5�3>WQy� ]U��h+>�^�>�Z�>�R�=�-�����$o�>ReW>��%>l�~=��:>�Z7�{I�=�7�>�2)>q%�<������=3=�=K�N����<|P�=�C��{�=h�G>e��hV��9J<z颽mؽ})�=t=�[��5z	<r�+>�m׼?6%=�Qо1�=j�ɽM�+>��!����>DD�D5����I�4�=��X�=&L>`=��#��?jQ�	S>(>��V��B��?j>>�aν�t��j~>9? �Y����B>?�= p��U�=^:=��<�=>i�>�=�>���>��?67?`�y�갾�H���M-�.�=����>>�&M>�|�	s���Vk��y��\���]�o w�#&ѽ/|?���x>Q7�>l�X=�B=��˽������=c���ӡ���~'���<Z|�>`Gk>���=o)>B�!�y���m����Կ8XݾZ�ؾͩ�I����=�ʠ�0xǽƅ����m�t	m��H��3���:���Vھ��s��>d�>'���q[���m�����3N���e����"�V<�>�\���(��}-��ʡ���.��yɽ�vr�g�B��ν:
�>#j�>B�-���k�>8lU>�h6>���>f��kl�0s+>%��>w�>���>��>��<�r�>��>$�^> 2�)4�����=��W=g�M��0>��z>1׽kP�)N�=O���T�6V->i�ݽ��̽;tH�&MF�����>z�>�q9>���#�,7�B����3e>�?��;��@d�[C�`߿�������ٽ����q�J���S7�=
B�:j��=���:~�=a^��)�W>��>�����43���=�=sb�$�C=G�ν��*1�`�"�f,>��>�2i>��?vT?��/?W�>��k���P��	����=�� �=B�>/� ?t>j���	?���D���0���Ǿ��=�K�<�w�>�E���$����:�������>�l�>�r�4����B>W�>�z�>��?��>1@��Y�|�
�Ο�YNƿ����ξ%=����;�c����l���2��W>sG�=�OȾ�nо��t=V�j=�f>8|�>��U>�x�<��[�)����O���G����¾zs�� {�&[(>&Z[��=��� �*�����n���QҴ<���.�����
����.$�>��>��>���>��>�B�>؍>��{�^+?��b`����<�;�>��j>q��>u��>���>8���ij��|/��0KK��Hn=�S>ơ�=i�>Y)�>����ͽ�_�>�>�(;�D�\0��8=z��θ&>��k>��_>ٺ?s�<Å� ���xH������=�Hw>p�.�轓`N��6�>9�m�nW�k�	�N[��#��z�>�Y�>�=>�4=nNp<՝=KZ����务=���=Gu���~�>�!=��U�=/�0��6׽rS�A6�=75=���=bɂ>Rw9?i�f?'�b?0�>\�߽�0Y��m>��F��=F�>s{?�Y�>�e�>L�|�}翾oG��>��а��Ȁ*�plu��.?�d��A�<��S>�[��Ob�����C�>s�e���>�A�=^[�>夽>.�>H�>�\>􎆾Q5�|���d�9�2��h��x��
����F>0<�=��v<�Dp�zp޾�	��O�~��9�>��>n�U>�O)�.���졾�f���
�#|����msJ��,���7��=�S4�P����<v��4�3t���*���_u��[��ƾ��'�t=�<,��=`T��� �=.2*>���>�;�>D�9>^�+=s�?,��=8�2>��k�y�c>��>�6�>��?�i?,����x#���<�k���>���=�o�=o3�>��=�i����6�0 ��ިX�!�y=G��.��� �=�{=��=��M>X��=���>�����%��h��L���	<��=��>���LSB�S��>nQ��K���tf���󔾐,��> ��>!��>��>+�۽M:{=r�?��$�:F��=.��=�=�ef�=���=��>k�[�� ���.@�Xdͽ`���#N
>QLq>�s�>Z?�a? �@?6M�>Ez�x�S��G[�vߋ��l>��>!�O>��><�����پ�р��F�Z��'��5Fa>�8�=(�<�5��>���=<���eu轌t>�aP����<�O���Ma>�q?>��>��>�(��D��!	����ֿ�Ъ�[���z��А��v�y6���t��=�k:�#������ʾ�uM�J��>}�>F,#���1��ֽ��Uꔾg�X��P��	�оo�ƾ����'n>�|��:��q�˾��1����:`�FS"���Ľ����Bh��y��ߋ>U��>�<��:$���=I;8>R9?v=�>��>Vt����?�
�<�=��3?��>��>2��>x;R����'^s��W��Y0>=e>�$�=@��=N�W����*e>.M>:�=��5�����g3�f�����7>�%M>�>yaE>���=����k
�i�"��y����> #?6-%�� Q���~��%�=q�=5��5�3��ű��b����ԽW��<�͚>�.>\�|��y=�3���zt*�h��=��=�������LӨ;2,$>I��=�t��%G��.J��]K��⽽��=�9�>Y�!?	�>?�}I?�>��:��b_�R33���0=`_�>��
?S��>��ֽв
����ɧ �y��.�#��u$>�ͮ�ٴ��a�=���=�6�>-�t;�F��O��07>��ֽ���<�����QN=�kg>/��>x��>��>�7���<�;��6!���оN/߾NiP��z�y2���%�E	D���=C��Ծ6h�5���ɘ>e�,>��=ݍ��^0���]���=t;=Ջ�;�ɾ�r���l��J>�(߽NŽ-�ּ��=t��������2����N���LZ����E|�>��\>�\>lp{>�}?u?�{>3�ڐ"?�Ԍ�I���!����>�n�>s\@>�B�>�v?�7,>�3��&����;���#>z&�=͏D=ԎH>B�=����6�); @(>���[:"�˯���o��y7�<ؘ>9��=)ǻ>��D>>���5>����
"��*�3�����?ֺ���dC��T�>�4�/��-��{���E��k�=��>�=w�p=�ٽ���qR0=[�$I>Sm=1���B=��7=�g�=�q�?��{�C�%�T��;���>#��=�DZ=���>��?!�>ܶz=�����DF��z��#+>Ϫ�>,�>��ͽi�ڽ�.ɾ�4�/������������'�ֆ�=;�>JN,=>�@>I%>��������g�>����=�jI>�x(��V=���=��4>7<>�C�|�rK���(������Og��ؼn���� �L\ɽS8�=1{�)ʒ�ppF��Hֽ�)R���=��=�b���ǽ&�	��4���o����I���&����Xa۾����f>�V =��:�3FO� �t��>�)�=hA�=/ *;�Ӿ�%ͽ�Q?r=���>�>&�>+�?8o�>������>��>���<g��G��>�?:�>}�?��!?��=B�Q���=M�P� -�;�>���=c�=���= �<荿���*=�x �<��X\=��!=`>"=��h=��=Vpq=�=5]�=�F��g�ɾ����g��cƽ��;>U����߾ؗ��o�D<�#���I���H��q�I趻�=ۜ>�ְ>��>>1�8;x29�?���Q��_�o5��߲���a=i��=�{�=U�����e�,t�bk�p'�=�u=�#�='��=��J>ݚF?�^X?/c?r�>u����{�E"�A�=�5��>�C?�2<�������V�޾l(�y��Ya��/0{�F\�=?)�<w�����><�<e�<�>�=T�j�؟b��+<^c8>ن�>;��>oph>R��S�b=�� ��Qj����$̿�O�I�x�E��P��o�� %}�}u����ٽ�����9��Ia�;o{�>��=ǻ�=W"= ӽ�.�ϛ�>��p>)�~���r>��{����(E�h-X>=��􋤽&�����H&��w������XT_��р���Ǽ"��>���>��=��I=��> D�>1�>��>��>a[>r���4�7���>}�>]7|>�-S>��&>?U>��%�Ek���C��=HXx���=2'2>�8=a����=9��<g%��U�=�q#>�V>��=Q�L=)=7�>ʺ�#�;���>>��6]���Z������K��%g>G��=�O"��C�>u���wԦ�x�����<�_>˙5>���=���="�l=�Z	>*��=���<|�L�e��<X�l=9A�� 7����>���ERO�#�4=�c�<�@۽��#�������b��c���D>u��겁?t?�<u?򅹽�aӾ�eo��l�3y�>��L���ֽC�>�cw�_:����|����r	�m�_���ʾ�{<!)�>
E�<�CH>f�>�9����j�O�>ƞ�<�>H����>7Na>�T�>���=z�%�.���ﴔ=�|>��o�m��N�~��:ɾC���}I���,�L=��A>�#�;�x���"_>���=`��=�3u��>6<Fv9>e>���;�����|)վ'ξ�W��q��ԛ�<�B�<0�
N)<��)�W$:���P��,��L��)O<���=-D�='�>���->ݒ|�[酾�kW�$��>��>yw�>rL=��7��3��Ŭ�=f �<\u�>�05>͎S�6�<�`?>e��>p�o>��>:g�48K>���=�����*7>t�>����� �:��J>�:�=����#����=�(w>�,>u�=��g�s�|�a_�>��{����پT�ʾ�*~����>�%�<�����C>��ɾtu�N:(>�Z:>nE�=�8>��3� �>��>JK�=&�X>�c�=)�L��9��nUq�6i��J���v=ޝ)�>�v��OL�{S罰�k�aw�={)k>'�F�K��M>/O�;�}?��o?�e?�ڼŝY�� S�܄�=³�>���UZ��
�>�l������S���@�@'�F+�TS��q/��YbJ=�9%>~Nx=�kG>QC;�Z׽�fY=ͬ'>g�I>�Y�>ZE:>"��=M�u=��=�Z�<���<r�����q�������z�*����;䯴���4�������{1�*��z��I�=��=sw=؞>r �H����}X=˟?WYn�7�?O߽�����)	={'B>T�Ӿ�=>l��)ȣ�\C+��E��2��������Y�=�<>�u>�Z�r)���gs��>C�;>�"�>r��<��
=|�7>���>eQa>�᡼�M2����;��>��?�)�>�c8�b@��U��O��>>A�	>��y>��<�"�=�*�`�l����<�=i�=��n=�o�^�^��Ͱ=J,>NU^�5]�=�F��g�ɾ����g��cƽ��;>U����߾ؗ��o�D<�#���I���H��q�I趻�=ۜ>�ְ>��>>1�8;x29�?���Q��_�o5��߲���a=i��=�{�=U�����e�,t�bk�p'�=�u=�#�='��=��J>ݚF?�^X?/c?r�>u����{�E"�A�=�5��>�C?�2<�������V�޾l(�y��Ya��/0{�F\�=?)�<w�����><�<e�<�>�=T�j�؟b��+<^c8>ن�>;��>oph>R��S�b=�� ��Qj����$̿�O�I�x�E��P��o�� %}�}u����ٽ�����9��Ia�;o{�>��=ǻ�=W"= ӽ�.�ϛ�>��p>)�~���r>��{����(E�h-X>=��􋤽&�����H&��w������XT_��р���Ǽ"��>���>��=��I=��> D�>1�>��>��>a[>r���4�7���>}�>]7|>�-S>��&>?U>��%�Ek���C��=HXx���=2'2>�8=a����=9��<g%��U�=�q#>�V>��=Q�L=)=7�>ʺ�#�;���>>��6]���Z������K��%g>G��=�O"��C�>u���wԦ�x�����<�_>˙5>���=���="�l=�Z	>*��=���<|�L�e��<X�l=9A�� 7����>���ERO�#�4=�c�<�@۽��#�������b��c���D>u��겁?t?�<u?򅹽�aӾ�eo��l�3y�>��L���ֽC�>�cw�_:����|����r	�m�_���ʾ�{<!)�>
E�<�CH>f�>�9����j�O�>ƞ�<�>H����>7Na>�T�>���=z�%�.���ﴔ=�|>��o�m��N�~��:ɾC���}I���,�L=��A>�#�;�x���"_>���=`��=�3u��>6<Fv9>e>���;�����|)վ'ξ�W��q��ԛ�<�B�<0�
N)<��)�W$:���P��,��L��)O<���=-D�='�>���->ݒ|�[酾�kW�$��>��>yw�>rL=��7��3��Ŭ�=f �<\u�>�05>͎S�6�<�`?>e��>p�o>��>:g�48K>���=�����*7>t�>����� �:��J>�:�=����#����=�(w>�,>u�=��g�s�|�J��=ŭ��KOƾg/���̾	6?�_ԽjlU>��Q�k�ؽU��@x����Tg�u�z��1�=[8<���=��2�M��>mtQ�x���Q�<ȴh>h:+>u<�&q����<��>5ށ=�T>��O���=/����1�<��>��	=�S<��<�[?ŞK?�?h�K��%��������.=��>p��=�S��N�_i�=��=F*���u��"�;������T�=�(�=;C�����h��L-��쑣=�R=i��a�!�)���<!Y>�vg>i��h�c���=kd��U���4��,����GU�`��bߝ<�4�<{.�������I�e�~�0+<��[����<�j�=�xw�i��J);0�	=�?��>HA���|ؽ]���VӾ����	4�=*�����]��}�=�I�t���>X������ӛ�YG�\ڽ�����8��>�of��c�|�>�G$?�@?q!�>8sp>!ә>,�=�%�=Ms�=o�2>å�>��ؽ����=@=�̧=��8>܎������i�>�2<�2+=���=-��<������R�>=�	�=-�B=,�+=�v0�Z���c�=\D��
�<��=r1�>�⟾lV�e�վ��C�b��=��h=�/�>)����Ľ��6��H���fD<�*��
�=\{{>v��U��=��p> �>�h�<z#��K��=�[>�%��^c=�F��0�M���$�=�m>#ʙ<�����mfb>��Q=&:Ž81=�����z(?�l@?�f�>�����'�m���R��Ⱦ><~�>��>�٨=`���%�����78����v�����1<"<����=*�->����/��=�L=4|�=�=��r�7���l���!|>)=X>V�<=�?�����=�2=�H��U������Y���M��#+ѽ�S��$�������u�f�1=׾���\p����֒=�7>㧘=��<7"=��=��>�U鍾ng�"�Q��0
��w��(#e�gv�=Q@ؽ�%>���5{�sK�Ϧ/�#\��ю��kk��'����<Ϟ>��=e��=���>p*�>���>���>�~=Ɲ� �#��CR����="n�>uu�>�����?%�Zs�>�>�ם���Ƚ2���s>���=�w�<=�;��g��B����>5z>&Z<0Į��k��<���=���?�?�%=n>ʈ>Kj|�`�վ�8�ʾcЏ�2J��h�?��y�m����&���t�g�S�w�m>K�<�*�r̦=��>�ih�g��=rcD=���1���μx�<γ˽I��<��H�>��>l�U>=-��Y���[>�M�>�������@>Ed̽.�$?O�Y?�%?��ƾ�?��þ;�	>�8�>`ܺ=�K}=�W"�De5�X>�wB�*8���c�OrF>�y:�c�;=�F>l3���a>
4�;���+$>�{�?lu��)<*�>�_=k`�=ϭ=��=�?=�8�� 9���7��,��;������5�^�.<�W��S=j��9S6�&۠�/:�!���7�=��=�>B=�i�=/�>HИ=P��>'��=�a���虾�����NQȾ��>�C���	���Ŭ�=���;�Ԯ�c�p�8c�{1~=^6T��ߠ>��'������;	>t�?1��>��[>H�'��>�����4>-,`>=">µ��*#�d;A>�b�=�t�+�Խ�~.��潣��=�;3>�,ż��><N�V>1��=�>}�=����=����mN=�xQ>�x�;
H�X>aYp>�ؽ/=�Ã��T<�\۽�懾/��M&>ѳ�>˾>�P�=k���������<պ�>��<2s����=���>��#���k=��>����3����섽u�Y�Yh�S�&���ɼ�{��d7���N|=���<����TмEƻ=Oʁ� �=�d@<~�=�?��O?ԷG?1j���X��_߾���ҽ���m��=�8>ec,>����h� i+��U��%;�U*½]�ŽM�>b��E�6>P5>k�>n��<㌀>t�=�s;X$p>�����<ү>�J>"��=i�y��B�����U|����q�m��i��NG==]<���9��ș�`�R��M���j��6�=�&Q�8+��e��=ID>��5� 载�r?> �\���þ�p����^�۽� A�X#t���<�7
���G���=a��=��=��.�����W�C��}���t�PI�z̏>�����ͼ���a�?N��>;��=\\὜*������8z�>=��>�*X�Y���=s��>:i=�A���Q>>��z=�8����=D�w<.��<Q�C=nu�=9ˀ=�n=�l>mf�W��� =��->�
D���I�%�f>���=��=J��=ŭ��KOƾg/���̾	6?�_ԽjlU>��Q�k�ؽU��@x����Tg�u�z��1�=[8<���=��2�M��>mtQ�x���Q�<ȴh>h:+>u<�&q����<��>5ށ=�T>��O���=/����1�<��>��	=�S<��<�[?ŞK?�?h�K��%��������.=��>p��=�S��N�_i�=��=F*���u��"�;������T�=�(�=;C�����h��L-��쑣=�R=i��a�!�)���<!Y>�vg>i��h�c���=kd��U���4��,����GU�`��bߝ<�4�<{.�������I�e�~�0+<��[����<�j�=�xw�i��J);0�	=�?��>HA���|ؽ]���VӾ����	4�=*�����]��}�=�I�t���>X������ӛ�YG�\ڽ�����8��>�of��c�|�>�G$?�@?q!�>8sp>!ә>,�=�%�=Ms�=o�2>å�>��ؽ����=@=�̧=��8>܎������i�>�2<�2+=���=-��<������R�>=�	�=-�B=,�+=�v0�Z���c�=\D��
�<��=,*�>>6=������	��.������>I��>x��T2�>�6�"�����~W	����Hh>��>$)�>Pj�U�>m"�<G���5L>�<>G.L<c2�Jx�y��.�= �f>�����"�����ʽ�<�2I>�1A>�J˽�;нU9^?��?9^??��<�b���t�,�:�\sK>����>P'$>̝޼�ڇ>>.x>�c���*EL�"���^�����=�G���c�=x�=����8��v>tV>>��c=$=���=4֗>���>�[�>�<�L�y�Ȼ�0l�zr�ކ��eU9�q����=�j����]=�[=�G����b��S��o�ͽ*νI93>wZt>�6>ru�<��8�):�=ٿ�u���J[�� �[$ݾL��n ���� �=�AF.�C���/o>�;��sR�AI�s�)��3��韾���a?k �"���<e�=��$?U�?gٌ>w1�=e]�=ɘ2�9�{���{=_x?U�f>��齤�C�&w��.�>�@?&=6�1�Wʔ>��=��n�>GZ�>�5�?��=��=K���-Q��#>��	>>r��ռ�z׽�S��o@>	|�>��C�p. �x̾�iV��8�����>~ ?;߿����>��>j/k�g���ɾ���L�=X3u>��>�)=0t'>�z<�շ�I2~>Ck�>��	>��<v����Ͻ� `>|l�=�Ģ=\�<���M��������>�E>�P+<��V��?
@�?��3?���>� �d�����O�0��>_�$�y��>�$>�V&>&�>��=/3������?�j^̾M1꼟��=����f�1�=�X��ɽK�=y�&>�D���H�=B@'>=��>9ב>{�z=|�_�&=+T =������U㘿��о�:�����i��=O>#1����ټ��½p�k��b��`�R=��O=��>�#�=�������6Ϊ;���wF�<�轓c�iԾ�̑��=�����S�R���S��N���y|��욾T`b�Y��@a����(}��?R���M���G#>�� ?��-?��>�;�e��;FJ>@ �g!r>�5�>�ɡ=�Ҽ�_V>@K�>I̯>p~�>�ڼ�����~;>���m��(��<��>�-�;��^=ե��K��nF�P��w'=y%>��>L�����Խ��>b��>L�����Ǿ�-s��-����<Mv>?���� ���<ج¾n���ɾ[Lɾ�ͽޚ\>�Dd>��Q>����oGV>K30����=�hw>�����&O>�/H��[��� >����3>橧=�kH�)�߽0��L����Dּ"c>0�=q䇽��Y?�@?�"?�(�:Yr��>_���B���>*sR����>7μ�K>��2<�A���K̾�I�ݵ���	�;�Wν��?>2t]�1�X��C�>�Ƚ`d�-\�=���=T�׻=q�;炊=�U->�m>CxS>��a�����+���Z���0޿A���-��
����;��U�]�%�6>å�=��q��<�H����݋�z�=�N�=!��>�w;= ��;�2��=�d��u��d>cq��vhþ�Y�b���};�t?��2f��
˽e�m�{���:�o��Æ�q�t�ۊ��!��U�ؾ�-����>o�����ݽ�����6?�b�>cz�>kx�>�Dн��3>�$�=���=w] >S�>�>� �=�x�>�x�>�G<��]�ԦȽ�8�>Vu�<�f;>~>ܲ�>#��>�����>��y�&����H<�|�<�vM>��6>]�>UE<��=,*�>>6=������	��.������>I��>x��T2�>�6�"�����~W	����Hh>��>$)�>Pj�U�>m"�<G���5L>�<>G.L<c2�Jx�y��.�= �f>�����"�����ʽ�<�2I>�1A>�J˽�;нU9^?��?9^??��<�b���t�,�:�\sK>����>P'$>̝޼�ڇ>>.x>�c���*EL�"���^�����=�G���c�=x�=����8��v>tV>>��c=$=���=4֗>���>�[�>�<�L�y�Ȼ�0l�zr�ކ��eU9�q����=�j����]=�[=�G����b��S��o�ͽ*νI93>wZt>�6>ru�<��8�):�=ٿ�u���J[�� �[$ݾL��n ���� �=�AF.�C���/o>�;��sR�AI�s�)��3��韾���a?k �"���<e�=��$?U�?gٌ>w1�=e]�=ɘ2�9�{���{=_x?U�f>��齤�C�&w��.�>�@?&=6�1�Wʔ>��=��n�>GZ�>�5�?��=��=K���-Q��#>��	>>r��ռ�z׽�S��o@>	|�>��C�p. �x̾�iV��8�����>~ ?;߿����>��>j/k�g���ɾ���L�=X3u>��>�)=0t'>�z<�շ�I2~>Ck�>��	>��<v����Ͻ� `>|l�=�Ģ=\�<���M��������>�E>�P+<��V��?
@�?��3?���>� �d�����O�0��>_�$�y��>�$>�V&>&�>��=/3������?�j^̾M1꼟��=����f�1�=�X��ɽK�=y�&>�D���H�=B@'>=��>9ב>{�z=|�_�&=+T =������U㘿��о�:�����i��=O>#1����ټ��½p�k��b��`�R=��O=��>�#�=�������6Ϊ;���wF�<�轓c�iԾ�̑��=�����S�R���S��N���y|��욾T`b�Y��@a����(}��?R���M���G#>�� ?��-?��>�;�e��;FJ>@ �g!r>�5�>�ɡ=�Ҽ�_V>@K�>I̯>p~�>�ڼ�����~;>���m��(��<��>�-�;��^=ե��K��nF�P��w'=y%>��>L�����Խ��>j7?��I�+��(�����o�={�>� ?�f�����=���>��2<B��6W���Y����A��J�>-��>�>�7>��;�"�=B��<KQ>�T�=�m�=�������#�|b�Ӭ�r��-�ν(�7�=��>�v��=,n=F>>�G?	@I?�5H?�c����:�<���&����>1��
�����=zҽ��B�\�W�����5��#F�  =OQ>;�P��儽��#=��&=l<>� Ew=OZ>�aq��	>74:>���>qT�> �=�'�����ɥ�����<ӱ�7��ˁ��+���j�=Cu���҃<nC���-����پ�`ݾ�W��g���V=K��<�ٽc��`��>�x$���(�AMᾫY��,��7j�rH.���;>=M������읜����397��g=J�FY�#��k��-��>g��>���>d�6=d?���>i��>�*�<��>﹤>y�B�eN�;#��>-?�F?�û>3����O��:X��:@����/`>�fv>ӊ{���;�>�ӽ�����='a!<0x���3���l��¼���=v�7>���k:ϼ���>,�n��(�J���S�����)�N��i(?Έ侾t&��&���ھ���~��/�;�Zg>���>���>�Ϗ=<W>n>�=p��=�d=�^L>c�=J*O�9kE�s,���T����"��v�ۼ�����$�W�!>G���,�=��=z�n>��V?/*?��>|Ͼ6k�r�'���痲>4�[�ӰI>m�->_��=���E�Ѿ2�$&'�@�Ծ[�<"g��xi>7>������:��ؽ%y+���<>rWh>�!=�#<p�=4��>S��=���=�&���q�8���>�.���Q¿��۾��5�؋����e=��,>Ǫ[�$�� ��+U����ý+>-8m>	mg>�x>$>m>%l7>b-|>��J�h��=|
��k������2���p���T&>�S���L�h��C��z=���
����;��$�W}�.ą��u���+>� �=���>jL�> #?�y�>Q&?��� R>�,
?Q�A>��>m �>2z�>r�3>4=�E>��?o���׽�����4�k�7>R�ý���=�ۓ>Û�:f7C;�� >�t.>|�a=-ĥ�;��=�QU�����&x>���=��F>���>,�n��(�J���S�����)�N��i(?Έ侾t&��&���ھ���~��/�;�Zg>���>���>�Ϗ=<W>n>�=p��=�d=�^L>c�=J*O�9kE�s,���T����"��v�ۼ�����$�W�!>G���,�=��=z�n>��V?/*?��>|Ͼ6k�r�'���痲>4�[�ӰI>m�->_��=���E�Ѿ2�$&'�@�Ծ[�<"g��xi>7>������:��ؽ%y+���<>rWh>�!=�#<p�=4��>S��=���=�&���q�8���>�.���Q¿��۾��5�؋����e=��,>Ǫ[�$�� ��+U����ý+>-8m>	mg>�x>$>m>%l7>b-|>��J�h��=|
��k������2���p���T&>�S���L�h��C��z=���
����;��$�W}�.ą��u���+>� �=���>jL�> #?�y�>Q&?��� R>�,
?Q�A>��>m �>2z�>r�3>4=�E>��?o���׽�����4�k�7>R�ý���=�ۓ>Û�:f7C;�� >�t.>|�a=-ĥ�;��=�QU�����&x>���=��F>8��>n=�p����������B��R�>�V�>6�����&=�������3�־E=�+�=�ON>r4>%���y�>��>D���L=�>b=��Q=��=1 ��B="x��&b=�]��J��[�˽�Nؽ�!>�D�>�M>x�=��!��0>T@?�$D?5?�"���PȾm:�x?�ys�=��=�Li�����>�}�>�eY��n轠��qf4��\��|�c�J���_=b��=h=`=n6=]0L�20v�n�=���=:�Q��<h=�e�=���=bpZ=X��=�R�=��=�G�<
l>������ʿ��žz?
��~�=5#ٽ�w=	ב��^<������o�!>1>�k�>چ]>�}��{b���æ=5x>�闾,��2�ڙ���o����ʾ�YZ�!8�>�2��Z��o�,��'��~�8�ݽ��I�x�����iн2 �����>��=�X>�5���.?�,?ۻ����>B��=0%S>u �>'�P�JY-���k�.�Ͻ�|�>N��>�G?�<��+�V��V�<���=U=�H=J@�=�B>�co���<M�C>���=���>W�5>@r�=���gF��a	�)D�"�=>8��>n=�p����������B��R�>�V�>6�����&=�������3�־E=�+�=�ON>r4>%���y�>��>D���L=�>b=��Q=��=1 ��B="x��&b=�]��J��[�˽�Nؽ�!>�D�>�M>x�=��!��0>T@?�$D?5?�"���PȾm:�x?�ys�=��=�Li�����>�}�>�eY��n轠��qf4��\��|�c�J���_=b��=h=`=n6=]0L�20v�n�=���=:�Q��<h=�e�=���=bpZ=X��=�R�=��=�G�<
l>������ʿ��žz?
��~�=5#ٽ�w=	ב��^<������o�!>1>�k�>چ]>�}��{b���æ=5x>�闾,��2�ڙ���o����ʾ�YZ�!8�>�2��Z��o�,��'��~�8�ݽ��I�x�����iн2 �����>��=�X>�5���.?�,?ۻ����>B��=0%S>u �>'�P�JY-���k�.�Ͻ�|�>N��>�G?�<��+�V��V�<���=U=�H=J@�=�B>�co���<M�C>���=���>W�5>@r�=���gF��a	�)D�"�=>Ɓ>ԳR�%����Y�A������]=��=K�:=�B��Jj=\e���߾G��Z�羄�=�T5>n��>M�O>/h�>�g%>�oP��ҍ�=/�=��=љ���H�=7�c>�2�<��%>���<�5��$��(:�=�5�>N�=@M ����=�~o?.R�?
�Z?�;�>A�2���j����oA>��>�ܾ5+>qܨ�d���٣�䰂���	�]�S�D)�&|=��-=O������=�@6=�]ƽ��=U��$"�=!�1=6�V�3�Z>c�>_��=w[$�����v��Nc�<5��^Ŀ�ʾ�N&��>���>$���a�g.�����v�-\��P�۽�>��-?$w�>����'��M��6���X�?��ak����}��	�X�D�E0�=c�o��޾zֽ�ᙾ/갾/�p�#Qd�Ώ��桾�e�R�	�f�>�<烸�*P����<B��>21?9�>J���]��萶>��>���>�W�>{�_<�Ћ�=J>?Ϋ>�(�>���4�k�[S>pf>3Bd�ļ����	=�����d�</J�ųɼSx*<���oF>rT�=`:�	����g=�u�<��~>�����T��u��������ٽ�N�>�ư>Uw�N*�f4�������� �o�6>S�k>��b>kt�> �=��=�d�=��w=�>�sg>Ya�=���<�wu���ϼ��=������<=�g���<�d�1�=Mw>g��;�;���hʽ	܁?���?h\?���>X�c{�1 o��z�����>F���k��`N��	^�Ԑ��Cp%�P`Y���!�=����>>fO�<F�}��i�<��h�>&j
>�k<䳋>N��=P�=�=Ǖ�=�1�>�����==�B=���}w�e边��8�m���:�`�<��=w��E֠�C:a�, ݽe��=c�>}*�=� �=MH��=�<E���Qv��R�@����B��b5$�±ž�ѽ�C�>.ˍ�`s��"x��=NG�|$�:����d#�!iw�r��x�c���<B��>%��ª�b���a�\>H�	?�gp>�Oo>�D~>�v�J�L>���>���>cd>�	>��<$~�>,y�=��>Y���0�<�؇=9��F�o=�_��ނ=�?����<���<��
ݼ�j�@/��/>¼>�� >��,"��Ɓ>ԳR�%����Y�A������]=��=K�:=�B��Jj=\e���߾G��Z�羄�=�T5>n��>M�O>/h�>�g%>�oP��ҍ�=/�=��=љ���H�=7�c>�2�<��%>���<�5��$��(:�=�5�>N�=@M ����=�~o?.R�?
�Z?�;�>A�2���j����oA>��>�ܾ5+>qܨ�d���٣�䰂���	�]�S�D)�&|=��-=O������=�@6=�]ƽ��=U��$"�=!�1=6�V�3�Z>c�>_��=w[$�����v��Nc�<5��^Ŀ�ʾ�N&��>���>$���a�g.�����v�-\��P�۽�>��-?$w�>����'��M��6���X�?��ak����}��	�X�D�E0�=c�o��޾zֽ�ᙾ/갾/�p�#Qd�Ώ��桾�e�R�	�f�>�<烸�*P����<B��>21?9�>J���]��萶>��>���>�W�>{�_<�Ћ�=J>?Ϋ>�(�>���4�k�[S>pf>3Bd�ļ����	=�����d�</J�ųɼSx*<���oF>rT�=`:�	����g=�u�<��~>�����T��u��������ٽ�N�>�ư>Uw�N*�f4�������� �o�6>S�k>��b>kt�> �=��=�d�=��w=�>�sg>Ya�=���<�wu���ϼ��=������<=�g���<�d�1�=Mw>g��;�;���hʽ	܁?���?h\?���>X�c{�1 o��z�����>F���k��`N��	^�Ԑ��Cp%�P`Y���!�=����>>fO�<F�}��i�<��h�>&j
>�k<䳋>N��=P�=�=Ǖ�=�1�>�����==�B=���}w�e边��8�m���:�`�<��=w��E֠�C:a�, ݽe��=c�>}*�=� �=MH��=�<E���Qv��R�@����B��b5$�±ž�ѽ�C�>.ˍ�`s��"x��=NG�|$�:����d#�!iw�r��x�c���<B��>%��ª�b���a�\>H�	?�gp>�Oo>�D~>�v�J�L>���>���>cd>�	>��<$~�>,y�=��>Y���0�<�؇=9��F�o=�_��ނ=�?����<���<��
ݼ�j�@/��/>¼>�� >��,"��OI��	���龼������Q�	;��>�Ѿ	;����>�T��������%c��BA��b!,>��*?�v?>�ܧ>r'���i��̕�h��=�j>VB>�K	>d�=p<��:����=髦=�W >7�P=rF >�C>��>Pί;�з=?@b?�{?\g?��>y�Ǿ��M��D�US�>��=˾=aq>��^���ω�08��FLu=�bϾ�]T��Qɾf�|�>L��>rd�=.�==F������{�:>yX��#�<ࢂ<Pz`�B韽Y�W��"(=s�J����;��<���T��Ϳ�_ �LF�yz�0�>9h^���</m�L���~���S�T0*�ϟ�=��?ꀄ>�>(��A*K�G>��Ͼ���Qr=�q��zǛ��pG�G��ai�:w��f���I�# ��|Q��15�dtľ�M̾�������V'>���>}��=W��=��>}�0>s5?4��>c3�=�{}>.dɺ*��f�
>��>�?9�?TKR>�I�=�4�Ӯ��o�� =v[,=��<|�z�Og6���D=�/��N
>�Iܼq��={��<��e<ۥ�=�7�=j;�Q%�4½��=